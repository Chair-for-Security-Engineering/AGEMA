/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_Pipeline_d1 (SI_s0, clk, SI_s1, Fresh, SO_s0, SO_s1);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [867:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(1)) U1938 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_943, n2796}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1939 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_945, n2810}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1940 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_947, n2462}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1941 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_949, n2760}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1942 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_951, n2791}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1944 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_953, n2813}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1945 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_955, n2630}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1946 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_957, n2765}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_927 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( new_AGEMA_signal_2745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( new_AGEMA_signal_2747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( new_AGEMA_signal_2749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( new_AGEMA_signal_2751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( new_AGEMA_signal_2753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( new_AGEMA_signal_2755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( new_AGEMA_signal_2757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( new_AGEMA_signal_2759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_2761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_2763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C ( clk ), .D ( n2630 ), .Q ( new_AGEMA_signal_2765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C ( clk ), .D ( new_AGEMA_signal_955 ), .Q ( new_AGEMA_signal_2767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( new_AGEMA_signal_2769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( new_AGEMA_signal_2771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C ( clk ), .D ( n2462 ), .Q ( new_AGEMA_signal_2773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C ( clk ), .D ( new_AGEMA_signal_947 ), .Q ( new_AGEMA_signal_2775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C ( clk ), .D ( n2760 ), .Q ( new_AGEMA_signal_2777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C ( clk ), .D ( new_AGEMA_signal_949 ), .Q ( new_AGEMA_signal_2779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C ( clk ), .D ( n2796 ), .Q ( new_AGEMA_signal_2781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C ( clk ), .D ( new_AGEMA_signal_943 ), .Q ( new_AGEMA_signal_2783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C ( clk ), .D ( n2765 ), .Q ( new_AGEMA_signal_2785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C ( clk ), .D ( new_AGEMA_signal_957 ), .Q ( new_AGEMA_signal_2787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C ( clk ), .D ( n2791 ), .Q ( new_AGEMA_signal_2789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C ( clk ), .D ( new_AGEMA_signal_951 ), .Q ( new_AGEMA_signal_2791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_2793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_2795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C ( clk ), .D ( n2813 ), .Q ( new_AGEMA_signal_2797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C ( clk ), .D ( new_AGEMA_signal_953 ), .Q ( new_AGEMA_signal_2799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C ( clk ), .D ( n2810 ), .Q ( new_AGEMA_signal_2801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C ( clk ), .D ( new_AGEMA_signal_945 ), .Q ( new_AGEMA_signal_2803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_3317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_3323 ) ) ;

    /* cells in depth 2 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1937 ( .a ({new_AGEMA_signal_943, n2796}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[0] ), .c ({new_AGEMA_signal_970, n2719}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1943 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1023, n2672}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1947 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[1] ), .c ({new_AGEMA_signal_958, n2635}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1948 ( .a ({new_AGEMA_signal_947, n2462}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[2] ), .c ({new_AGEMA_signal_971, n2641}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1949 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[3] ), .c ({new_AGEMA_signal_959, n2790}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1950 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[4] ), .c ({new_AGEMA_signal_960, n2519}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1951 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_972, n2750}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1952 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[5] ), .c ({new_AGEMA_signal_973, n2615}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1953 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1024, n2640}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1955 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[6] ), .c ({new_AGEMA_signal_974, n2699}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1956 ( .a ({new_AGEMA_signal_974, n2699}), .b ({new_AGEMA_signal_1025, n2737}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1957 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[7] ), .c ({new_AGEMA_signal_975, n2816}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1958 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1026, n2767}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1961 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[8] ), .c ({new_AGEMA_signal_976, n2780}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1962 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1027, n2789}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1963 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .r ( Fresh[9] ), .c ({new_AGEMA_signal_977, n2317}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1965 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[10] ), .c ({new_AGEMA_signal_978, n2694}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1966 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1028, n2769}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1969 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[11] ), .c ({new_AGEMA_signal_979, n2073}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1970 ( .a ({new_AGEMA_signal_979, n2073}), .b ({new_AGEMA_signal_1029, n2707}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1971 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[12] ), .c ({new_AGEMA_signal_961, n2315}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1972 ( .a ({SI_s1[0], SI_s0[0]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[13] ), .c ({new_AGEMA_signal_962, n2682}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1973 ( .a ({new_AGEMA_signal_962, n2682}), .b ({new_AGEMA_signal_980, n2713}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1975 ( .a ({new_AGEMA_signal_953, n2813}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[14] ), .c ({new_AGEMA_signal_981, n2723}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1976 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1031, n2688}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1978 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[15] ), .c ({new_AGEMA_signal_982, n2725}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1979 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1032, n2541}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1984 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[16] ), .c ({new_AGEMA_signal_983, n2815}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1985 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1033, n2086}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1987 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[17] ), .c ({new_AGEMA_signal_984, n2600}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1990 ( .a ({new_AGEMA_signal_947, n2462}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[18] ), .c ({new_AGEMA_signal_985, n2538}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1991 ( .a ({new_AGEMA_signal_985, n2538}), .b ({new_AGEMA_signal_1035, n2786}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1995 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[19] ), .c ({new_AGEMA_signal_963, n2595}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1996 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_986, n2742}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1999 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[20] ), .c ({new_AGEMA_signal_987, n2753}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2000 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1037, n2577}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2004 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[21] ), .c ({new_AGEMA_signal_988, n2400}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2008 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[22] ), .c ({new_AGEMA_signal_989, n2785}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2009 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1039, n2792}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2013 ( .a ({new_AGEMA_signal_953, n2813}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[23] ), .c ({new_AGEMA_signal_990, n2609}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2014 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_1040, n2724}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2017 ( .a ({new_AGEMA_signal_949, n2760}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[24] ), .c ({new_AGEMA_signal_991, n2661}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2018 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1041, n2174}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2020 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[25] ), .c ({new_AGEMA_signal_964, n2708}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2021 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_992, n2493}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2025 ( .a ({new_AGEMA_signal_943, n2796}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[26] ), .c ({new_AGEMA_signal_993, n2587}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2028 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1044, n2570}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2029 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[27] ), .c ({new_AGEMA_signal_965, n2559}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2035 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[28] ), .c ({new_AGEMA_signal_994, n2643}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2036 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1045, n2442}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2038 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_995, n2739}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2044 ( .a ({new_AGEMA_signal_947, n2462}), .b ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .r ( Fresh[29] ), .c ({new_AGEMA_signal_996, n2437}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2045 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[30] ), .c ({new_AGEMA_signal_966, n2261}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2046 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_997, n2778}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2052 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[31] ), .c ({new_AGEMA_signal_998, n2452}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2055 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1050, n2766}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2068 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[32] ), .c ({new_AGEMA_signal_1000, n2772}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2070 ( .a ({new_AGEMA_signal_951, n2791}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[33] ), .c ({new_AGEMA_signal_1001, n2824}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2071 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1053, n2612}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2074 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_1054, n2313}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2089 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[34] ), .c ({new_AGEMA_signal_1002, n2395}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2090 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1058, n2818}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2094 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[35] ), .c ({new_AGEMA_signal_967, n2779}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2096 ( .a ({new_AGEMA_signal_955, n2630}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[36] ), .c ({new_AGEMA_signal_1003, n2624}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2097 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[37] ), .c ({new_AGEMA_signal_968, n2242}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2100 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[38] ), .c ({new_AGEMA_signal_1004, n2356}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2119 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_1063, n2823}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2122 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[39] ), .c ({new_AGEMA_signal_1005, n2611}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2131 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1065, n2828}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2133 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[40] ), .c ({new_AGEMA_signal_1006, n2616}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2134 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1066, n2679}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2138 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[41] ), .c ({new_AGEMA_signal_1007, n2563}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2139 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1067, n2809}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2150 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_1068, n2709}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2163 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .r ( Fresh[42] ), .c ({new_AGEMA_signal_1008, n2401}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2211 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[43] ), .c ({new_AGEMA_signal_1010, n2061}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2232 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[44] ), .c ({new_AGEMA_signal_1011, n2721}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2276 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .r ( Fresh[45] ), .c ({new_AGEMA_signal_1012, n2298}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2278 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_1080, n2118}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2307 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[46] ), .c ({new_AGEMA_signal_1013, n2346}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2341 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[47] ), .c ({new_AGEMA_signal_1015, n2430}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2383 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[48] ), .c ({new_AGEMA_signal_969, n2712}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2402 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[49] ), .c ({new_AGEMA_signal_1017, n2777}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2615 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_947, n2462}), .clk ( clk ), .r ( Fresh[50] ), .c ({new_AGEMA_signal_1019, n2463}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2627 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[51] ), .c ({new_AGEMA_signal_1020, n2474}) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C ( clk ), .D ( new_AGEMA_signal_2745 ), .Q ( new_AGEMA_signal_2746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C ( clk ), .D ( new_AGEMA_signal_2747 ), .Q ( new_AGEMA_signal_2748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C ( clk ), .D ( new_AGEMA_signal_2749 ), .Q ( new_AGEMA_signal_2750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C ( clk ), .D ( new_AGEMA_signal_2751 ), .Q ( new_AGEMA_signal_2752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C ( clk ), .D ( new_AGEMA_signal_2753 ), .Q ( new_AGEMA_signal_2754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C ( clk ), .D ( new_AGEMA_signal_2755 ), .Q ( new_AGEMA_signal_2756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C ( clk ), .D ( new_AGEMA_signal_2757 ), .Q ( new_AGEMA_signal_2758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C ( clk ), .D ( new_AGEMA_signal_2759 ), .Q ( new_AGEMA_signal_2760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C ( clk ), .D ( new_AGEMA_signal_2761 ), .Q ( new_AGEMA_signal_2762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C ( clk ), .D ( new_AGEMA_signal_2763 ), .Q ( new_AGEMA_signal_2764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C ( clk ), .D ( new_AGEMA_signal_2765 ), .Q ( new_AGEMA_signal_2766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C ( clk ), .D ( new_AGEMA_signal_2767 ), .Q ( new_AGEMA_signal_2768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C ( clk ), .D ( new_AGEMA_signal_2769 ), .Q ( new_AGEMA_signal_2770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C ( clk ), .D ( new_AGEMA_signal_2771 ), .Q ( new_AGEMA_signal_2772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C ( clk ), .D ( new_AGEMA_signal_2773 ), .Q ( new_AGEMA_signal_2774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C ( clk ), .D ( new_AGEMA_signal_2775 ), .Q ( new_AGEMA_signal_2776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C ( clk ), .D ( new_AGEMA_signal_2777 ), .Q ( new_AGEMA_signal_2778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C ( clk ), .D ( new_AGEMA_signal_2779 ), .Q ( new_AGEMA_signal_2780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C ( clk ), .D ( new_AGEMA_signal_2781 ), .Q ( new_AGEMA_signal_2782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C ( clk ), .D ( new_AGEMA_signal_2783 ), .Q ( new_AGEMA_signal_2784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C ( clk ), .D ( new_AGEMA_signal_2785 ), .Q ( new_AGEMA_signal_2786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C ( clk ), .D ( new_AGEMA_signal_2787 ), .Q ( new_AGEMA_signal_2788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C ( clk ), .D ( new_AGEMA_signal_2789 ), .Q ( new_AGEMA_signal_2790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C ( clk ), .D ( new_AGEMA_signal_2791 ), .Q ( new_AGEMA_signal_2792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C ( clk ), .D ( new_AGEMA_signal_2793 ), .Q ( new_AGEMA_signal_2794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C ( clk ), .D ( new_AGEMA_signal_2795 ), .Q ( new_AGEMA_signal_2796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C ( clk ), .D ( new_AGEMA_signal_2797 ), .Q ( new_AGEMA_signal_2798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C ( clk ), .D ( new_AGEMA_signal_2799 ), .Q ( new_AGEMA_signal_2800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C ( clk ), .D ( new_AGEMA_signal_2801 ), .Q ( new_AGEMA_signal_2802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C ( clk ), .D ( new_AGEMA_signal_2803 ), .Q ( new_AGEMA_signal_2804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C ( clk ), .D ( new_AGEMA_signal_3317 ), .Q ( new_AGEMA_signal_3318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C ( clk ), .D ( new_AGEMA_signal_3323 ), .Q ( new_AGEMA_signal_3324 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_987 ( .C ( clk ), .D ( n2769 ), .Q ( new_AGEMA_signal_2805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_2807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C ( clk ), .D ( new_AGEMA_signal_2794 ), .Q ( new_AGEMA_signal_2809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C ( clk ), .D ( new_AGEMA_signal_2796 ), .Q ( new_AGEMA_signal_2811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C ( clk ), .D ( new_AGEMA_signal_2750 ), .Q ( new_AGEMA_signal_2813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C ( clk ), .D ( new_AGEMA_signal_2752 ), .Q ( new_AGEMA_signal_2815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C ( clk ), .D ( n2174 ), .Q ( new_AGEMA_signal_2817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C ( clk ), .D ( new_AGEMA_signal_1041 ), .Q ( new_AGEMA_signal_2819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C ( clk ), .D ( new_AGEMA_signal_2746 ), .Q ( new_AGEMA_signal_2821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C ( clk ), .D ( new_AGEMA_signal_2748 ), .Q ( new_AGEMA_signal_2823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C ( clk ), .D ( new_AGEMA_signal_2758 ), .Q ( new_AGEMA_signal_2825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C ( clk ), .D ( new_AGEMA_signal_2760 ), .Q ( new_AGEMA_signal_2827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C ( clk ), .D ( n2570 ), .Q ( new_AGEMA_signal_2829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_2831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C ( clk ), .D ( n2792 ), .Q ( new_AGEMA_signal_2833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C ( clk ), .D ( new_AGEMA_signal_1039 ), .Q ( new_AGEMA_signal_2835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C ( clk ), .D ( n2635 ), .Q ( new_AGEMA_signal_2837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C ( clk ), .D ( new_AGEMA_signal_958 ), .Q ( new_AGEMA_signal_2839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C ( clk ), .D ( n2587 ), .Q ( new_AGEMA_signal_2841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C ( clk ), .D ( new_AGEMA_signal_993 ), .Q ( new_AGEMA_signal_2843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C ( clk ), .D ( n2725 ), .Q ( new_AGEMA_signal_2845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C ( clk ), .D ( new_AGEMA_signal_982 ), .Q ( new_AGEMA_signal_2847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C ( clk ), .D ( n2708 ), .Q ( new_AGEMA_signal_2849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_2851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C ( clk ), .D ( n2818 ), .Q ( new_AGEMA_signal_2853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_2855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C ( clk ), .D ( n2790 ), .Q ( new_AGEMA_signal_2857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C ( clk ), .D ( new_AGEMA_signal_959 ), .Q ( new_AGEMA_signal_2859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C ( clk ), .D ( n2786 ), .Q ( new_AGEMA_signal_2861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C ( clk ), .D ( new_AGEMA_signal_1035 ), .Q ( new_AGEMA_signal_2863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C ( clk ), .D ( n2400 ), .Q ( new_AGEMA_signal_2865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C ( clk ), .D ( new_AGEMA_signal_988 ), .Q ( new_AGEMA_signal_2867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C ( clk ), .D ( new_AGEMA_signal_2762 ), .Q ( new_AGEMA_signal_2869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C ( clk ), .D ( new_AGEMA_signal_2764 ), .Q ( new_AGEMA_signal_2871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C ( clk ), .D ( n2815 ), .Q ( new_AGEMA_signal_2873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C ( clk ), .D ( new_AGEMA_signal_983 ), .Q ( new_AGEMA_signal_2875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C ( clk ), .D ( n2723 ), .Q ( new_AGEMA_signal_2877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C ( clk ), .D ( new_AGEMA_signal_981 ), .Q ( new_AGEMA_signal_2879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C ( clk ), .D ( n2709 ), .Q ( new_AGEMA_signal_2881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_2883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C ( clk ), .D ( n2753 ), .Q ( new_AGEMA_signal_2885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C ( clk ), .D ( new_AGEMA_signal_987 ), .Q ( new_AGEMA_signal_2887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C ( clk ), .D ( n2401 ), .Q ( new_AGEMA_signal_2889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_2891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C ( clk ), .D ( new_AGEMA_signal_2786 ), .Q ( new_AGEMA_signal_2893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C ( clk ), .D ( new_AGEMA_signal_2788 ), .Q ( new_AGEMA_signal_2895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C ( clk ), .D ( new_AGEMA_signal_2766 ), .Q ( new_AGEMA_signal_2897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C ( clk ), .D ( new_AGEMA_signal_2768 ), .Q ( new_AGEMA_signal_2899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C ( clk ), .D ( n2615 ), .Q ( new_AGEMA_signal_2901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C ( clk ), .D ( new_AGEMA_signal_973 ), .Q ( new_AGEMA_signal_2903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C ( clk ), .D ( n2643 ), .Q ( new_AGEMA_signal_2905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C ( clk ), .D ( new_AGEMA_signal_994 ), .Q ( new_AGEMA_signal_2907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C ( clk ), .D ( n2563 ), .Q ( new_AGEMA_signal_2909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_2911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C ( clk ), .D ( n2612 ), .Q ( new_AGEMA_signal_2913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C ( clk ), .D ( new_AGEMA_signal_1053 ), .Q ( new_AGEMA_signal_2915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C ( clk ), .D ( n2824 ), .Q ( new_AGEMA_signal_2917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C ( clk ), .D ( new_AGEMA_signal_1001 ), .Q ( new_AGEMA_signal_2919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C ( clk ), .D ( n2816 ), .Q ( new_AGEMA_signal_2921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C ( clk ), .D ( new_AGEMA_signal_975 ), .Q ( new_AGEMA_signal_2923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C ( clk ), .D ( n2073 ), .Q ( new_AGEMA_signal_2925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C ( clk ), .D ( new_AGEMA_signal_979 ), .Q ( new_AGEMA_signal_2927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C ( clk ), .D ( n2519 ), .Q ( new_AGEMA_signal_2929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C ( clk ), .D ( new_AGEMA_signal_960 ), .Q ( new_AGEMA_signal_2931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C ( clk ), .D ( n2616 ), .Q ( new_AGEMA_signal_2933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_2935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C ( clk ), .D ( new_AGEMA_signal_2790 ), .Q ( new_AGEMA_signal_2937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C ( clk ), .D ( new_AGEMA_signal_2792 ), .Q ( new_AGEMA_signal_2939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C ( clk ), .D ( n2780 ), .Q ( new_AGEMA_signal_2941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C ( clk ), .D ( new_AGEMA_signal_976 ), .Q ( new_AGEMA_signal_2943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C ( clk ), .D ( new_AGEMA_signal_2798 ), .Q ( new_AGEMA_signal_2945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C ( clk ), .D ( new_AGEMA_signal_2800 ), .Q ( new_AGEMA_signal_2947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C ( clk ), .D ( n2742 ), .Q ( new_AGEMA_signal_2949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C ( clk ), .D ( new_AGEMA_signal_986 ), .Q ( new_AGEMA_signal_2951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C ( clk ), .D ( n2724 ), .Q ( new_AGEMA_signal_2953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C ( clk ), .D ( new_AGEMA_signal_1040 ), .Q ( new_AGEMA_signal_2955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C ( clk ), .D ( n2317 ), .Q ( new_AGEMA_signal_2957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C ( clk ), .D ( new_AGEMA_signal_977 ), .Q ( new_AGEMA_signal_2959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C ( clk ), .D ( n2688 ), .Q ( new_AGEMA_signal_2961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_2963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C ( clk ), .D ( n2609 ), .Q ( new_AGEMA_signal_2965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C ( clk ), .D ( new_AGEMA_signal_990 ), .Q ( new_AGEMA_signal_2967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C ( clk ), .D ( n2672 ), .Q ( new_AGEMA_signal_2969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C ( clk ), .D ( new_AGEMA_signal_1023 ), .Q ( new_AGEMA_signal_2971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C ( clk ), .D ( n2640 ), .Q ( new_AGEMA_signal_2973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C ( clk ), .D ( new_AGEMA_signal_1024 ), .Q ( new_AGEMA_signal_2975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C ( clk ), .D ( n2713 ), .Q ( new_AGEMA_signal_2977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C ( clk ), .D ( new_AGEMA_signal_980 ), .Q ( new_AGEMA_signal_2979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C ( clk ), .D ( n2777 ), .Q ( new_AGEMA_signal_2981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C ( clk ), .D ( new_AGEMA_signal_1017 ), .Q ( new_AGEMA_signal_2983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C ( clk ), .D ( n2789 ), .Q ( new_AGEMA_signal_2985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_2987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C ( clk ), .D ( n2661 ), .Q ( new_AGEMA_signal_2989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C ( clk ), .D ( new_AGEMA_signal_991 ), .Q ( new_AGEMA_signal_2991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C ( clk ), .D ( new_AGEMA_signal_2774 ), .Q ( new_AGEMA_signal_2993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C ( clk ), .D ( new_AGEMA_signal_2776 ), .Q ( new_AGEMA_signal_2995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C ( clk ), .D ( n2694 ), .Q ( new_AGEMA_signal_2997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C ( clk ), .D ( new_AGEMA_signal_978 ), .Q ( new_AGEMA_signal_2999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C ( clk ), .D ( new_AGEMA_signal_2778 ), .Q ( new_AGEMA_signal_3001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C ( clk ), .D ( new_AGEMA_signal_2780 ), .Q ( new_AGEMA_signal_3003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C ( clk ), .D ( n2682 ), .Q ( new_AGEMA_signal_3005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C ( clk ), .D ( new_AGEMA_signal_962 ), .Q ( new_AGEMA_signal_3007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C ( clk ), .D ( new_AGEMA_signal_2802 ), .Q ( new_AGEMA_signal_3009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C ( clk ), .D ( new_AGEMA_signal_2804 ), .Q ( new_AGEMA_signal_3011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C ( clk ), .D ( n2624 ), .Q ( new_AGEMA_signal_3013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_3015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C ( clk ), .D ( n2356 ), .Q ( new_AGEMA_signal_3017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_3019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C ( clk ), .D ( n2778 ), .Q ( new_AGEMA_signal_3021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C ( clk ), .D ( new_AGEMA_signal_997 ), .Q ( new_AGEMA_signal_3023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C ( clk ), .D ( n2766 ), .Q ( new_AGEMA_signal_3025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C ( clk ), .D ( new_AGEMA_signal_1050 ), .Q ( new_AGEMA_signal_3027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C ( clk ), .D ( n2767 ), .Q ( new_AGEMA_signal_3029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_3031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C ( clk ), .D ( n2641 ), .Q ( new_AGEMA_signal_3033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C ( clk ), .D ( new_AGEMA_signal_971 ), .Q ( new_AGEMA_signal_3035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C ( clk ), .D ( n2719 ), .Q ( new_AGEMA_signal_3037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C ( clk ), .D ( new_AGEMA_signal_970 ), .Q ( new_AGEMA_signal_3039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C ( clk ), .D ( n2707 ), .Q ( new_AGEMA_signal_3041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C ( clk ), .D ( new_AGEMA_signal_1029 ), .Q ( new_AGEMA_signal_3043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C ( clk ), .D ( n2493 ), .Q ( new_AGEMA_signal_3045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C ( clk ), .D ( new_AGEMA_signal_992 ), .Q ( new_AGEMA_signal_3047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C ( clk ), .D ( n2577 ), .Q ( new_AGEMA_signal_3049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C ( clk ), .D ( new_AGEMA_signal_1037 ), .Q ( new_AGEMA_signal_3051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C ( clk ), .D ( n2541 ), .Q ( new_AGEMA_signal_3053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_3055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C ( clk ), .D ( n2679 ), .Q ( new_AGEMA_signal_3057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_3059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C ( clk ), .D ( n2699 ), .Q ( new_AGEMA_signal_3061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C ( clk ), .D ( new_AGEMA_signal_974 ), .Q ( new_AGEMA_signal_3063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C ( clk ), .D ( n2611 ), .Q ( new_AGEMA_signal_3065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C ( clk ), .D ( new_AGEMA_signal_1005 ), .Q ( new_AGEMA_signal_3067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C ( clk ), .D ( n2739 ), .Q ( new_AGEMA_signal_3069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C ( clk ), .D ( new_AGEMA_signal_995 ), .Q ( new_AGEMA_signal_3071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C ( clk ), .D ( n2772 ), .Q ( new_AGEMA_signal_3073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C ( clk ), .D ( new_AGEMA_signal_1000 ), .Q ( new_AGEMA_signal_3075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C ( clk ), .D ( n2442 ), .Q ( new_AGEMA_signal_3085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_3089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C ( clk ), .D ( n2779 ), .Q ( new_AGEMA_signal_3137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C ( clk ), .D ( new_AGEMA_signal_967 ), .Q ( new_AGEMA_signal_3141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C ( clk ), .D ( n2721 ), .Q ( new_AGEMA_signal_3173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C ( clk ), .D ( new_AGEMA_signal_1011 ), .Q ( new_AGEMA_signal_3177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C ( clk ), .D ( n2823 ), .Q ( new_AGEMA_signal_3201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C ( clk ), .D ( new_AGEMA_signal_1063 ), .Q ( new_AGEMA_signal_3205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C ( clk ), .D ( n2346 ), .Q ( new_AGEMA_signal_3221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C ( clk ), .D ( new_AGEMA_signal_1013 ), .Q ( new_AGEMA_signal_3225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C ( clk ), .D ( n2315 ), .Q ( new_AGEMA_signal_3241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C ( clk ), .D ( new_AGEMA_signal_961 ), .Q ( new_AGEMA_signal_3245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C ( clk ), .D ( new_AGEMA_signal_3318 ), .Q ( new_AGEMA_signal_3319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C ( clk ), .D ( new_AGEMA_signal_3324 ), .Q ( new_AGEMA_signal_3325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C ( clk ), .D ( new_AGEMA_signal_2754 ), .Q ( new_AGEMA_signal_3341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C ( clk ), .D ( new_AGEMA_signal_2756 ), .Q ( new_AGEMA_signal_3345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C ( clk ), .D ( n2600 ), .Q ( new_AGEMA_signal_3361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C ( clk ), .D ( new_AGEMA_signal_984 ), .Q ( new_AGEMA_signal_3365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C ( clk ), .D ( n2750 ), .Q ( new_AGEMA_signal_3397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C ( clk ), .D ( new_AGEMA_signal_972 ), .Q ( new_AGEMA_signal_3401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C ( clk ), .D ( new_AGEMA_signal_2782 ), .Q ( new_AGEMA_signal_3413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C ( clk ), .D ( new_AGEMA_signal_2784 ), .Q ( new_AGEMA_signal_3417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C ( clk ), .D ( n2737 ), .Q ( new_AGEMA_signal_3561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C ( clk ), .D ( new_AGEMA_signal_1025 ), .Q ( new_AGEMA_signal_3567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C ( clk ), .D ( n2785 ), .Q ( new_AGEMA_signal_3613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C ( clk ), .D ( new_AGEMA_signal_989 ), .Q ( new_AGEMA_signal_3619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C ( clk ), .D ( n2595 ), .Q ( new_AGEMA_signal_3845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C ( clk ), .D ( new_AGEMA_signal_963 ), .Q ( new_AGEMA_signal_3853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C ( clk ), .D ( n2437 ), .Q ( new_AGEMA_signal_3865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C ( clk ), .D ( new_AGEMA_signal_996 ), .Q ( new_AGEMA_signal_3873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C ( clk ), .D ( n2828 ), .Q ( new_AGEMA_signal_4017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C ( clk ), .D ( new_AGEMA_signal_1065 ), .Q ( new_AGEMA_signal_4025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C ( clk ), .D ( n2538 ), .Q ( new_AGEMA_signal_4189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C ( clk ), .D ( new_AGEMA_signal_985 ), .Q ( new_AGEMA_signal_4197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C ( clk ), .D ( n2809 ), .Q ( new_AGEMA_signal_4249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_4257 ) ) ;

    /* cells in depth 4 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1954 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ( Fresh[52] ), .c ({new_AGEMA_signal_1127, n2575}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1959 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[53] ), .c ({new_AGEMA_signal_1128, n1962}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1964 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ( Fresh[54] ), .c ({new_AGEMA_signal_1129, n1922}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1974 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[55] ), .c ({new_AGEMA_signal_1030, n2755}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1977 ( .a ({new_AGEMA_signal_977, n2317}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ( Fresh[56] ), .c ({new_AGEMA_signal_1130, n1926}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1980 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1032, n2541}), .clk ( clk ), .r ( Fresh[57] ), .c ({new_AGEMA_signal_1131, n1925}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1986 ( .a ({new_AGEMA_signal_1033, n2086}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ( Fresh[58] ), .c ({new_AGEMA_signal_1132, n2151}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1988 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[59] ), .c ({new_AGEMA_signal_1034, n2631}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U1989 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_1133, n2734}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1992 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ( Fresh[60] ), .c ({new_AGEMA_signal_1134, n2763}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1997 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[61] ), .c ({new_AGEMA_signal_1036, n1930}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2005 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ( Fresh[62] ), .c ({new_AGEMA_signal_1038, n2492}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2006 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1135, n2732}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2010 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2746}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[63] ), .c ({new_AGEMA_signal_1136, n1937}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2022 ( .a ({new_AGEMA_signal_2752, new_AGEMA_signal_2750}), .b ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .r ( Fresh[64] ), .c ({new_AGEMA_signal_1042, n1942}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) U2026 ( .a ({new_AGEMA_signal_993, n2587}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ( Fresh[65] ), .c ({new_AGEMA_signal_1043, n2676}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2030 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ( Fresh[66] ), .c ({new_AGEMA_signal_1139, n1944}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2037 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[67] ), .c ({new_AGEMA_signal_1140, n1950}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2039 ( .a ({new_AGEMA_signal_2756, new_AGEMA_signal_2754}), .b ({new_AGEMA_signal_995, n2739}), .clk ( clk ), .r ( Fresh[68] ), .c ({new_AGEMA_signal_1046, n1949}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2042 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[69] ), .c ({new_AGEMA_signal_1047, n2677}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2043 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1141, n2662}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2047 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[70] ), .c ({new_AGEMA_signal_1048, n2627}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2053 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_998, n2452}), .clk ( clk ), .r ( Fresh[71] ), .c ({new_AGEMA_signal_1049, n1957}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2056 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[72] ), .c ({new_AGEMA_signal_1142, n2088}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2062 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[73] ), .c ({new_AGEMA_signal_999, n1964}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2063 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2758}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[74] ), .c ({new_AGEMA_signal_1051, n2736}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2069 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2762}), .clk ( clk ), .r ( Fresh[75] ), .c ({new_AGEMA_signal_1052, n2673}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2072 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[76] ), .c ({new_AGEMA_signal_1144, n2761}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2073 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1323, n2720}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2075 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ( Fresh[77] ), .c ({new_AGEMA_signal_1145, n2412}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2076 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_1324, n2417}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2079 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_966, n2261}), .clk ( clk ), .r ( Fresh[78] ), .c ({new_AGEMA_signal_1055, n2571}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2080 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1146, n2505}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2081 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ( Fresh[79] ), .c ({new_AGEMA_signal_1056, n2651}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2083 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2762}), .clk ( clk ), .r ( Fresh[80] ), .c ({new_AGEMA_signal_1147, n2359}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2086 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[81] ), .c ({new_AGEMA_signal_1057, n2101}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2087 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1148, n2625}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2091 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[82] ), .c ({new_AGEMA_signal_1059, n2190}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2095 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[83] ), .c ({new_AGEMA_signal_1060, n1976}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2098 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ( Fresh[84] ), .c ({new_AGEMA_signal_1150, n2535}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2101 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .r ( Fresh[85] ), .c ({new_AGEMA_signal_1151, n1973}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2105 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[86] ), .c ({new_AGEMA_signal_1061, n2690}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2111 ( .a ({new_AGEMA_signal_992, n2493}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2766}), .clk ( clk ), .r ( Fresh[87] ), .c ({new_AGEMA_signal_1062, n2817}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2113 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[88] ), .c ({new_AGEMA_signal_1153, n2741}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2118 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ( Fresh[89] ), .c ({new_AGEMA_signal_1154, n1992}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2120 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[90] ), .c ({new_AGEMA_signal_1155, n1991}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2123 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ( Fresh[91] ), .c ({new_AGEMA_signal_1064, n1993}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2125 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[92] ), .c ({new_AGEMA_signal_1156, n1995}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2132 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[93] ), .c ({new_AGEMA_signal_1157, n2241}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2135 ( .a ({new_AGEMA_signal_2772, new_AGEMA_signal_2770}), .b ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .r ( Fresh[94] ), .c ({new_AGEMA_signal_1158, n2003}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2140 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ( Fresh[95] ), .c ({new_AGEMA_signal_1159, n2008}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2141 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ( Fresh[96] ), .c ({new_AGEMA_signal_1160, n2572}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2143 ( .a ({new_AGEMA_signal_1067, n2809}), .b ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .r ( Fresh[97] ), .c ({new_AGEMA_signal_1161, n2004}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2147 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[98] ), .c ({new_AGEMA_signal_1162, n2009}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2151 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2766}), .clk ( clk ), .r ( Fresh[99] ), .c ({new_AGEMA_signal_1163, n2533}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2157 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[100] ), .c ({new_AGEMA_signal_1069, n2026}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2158 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .r ( Fresh[101] ), .c ({new_AGEMA_signal_1164, n2022}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2159 ( .a ({new_AGEMA_signal_2776, new_AGEMA_signal_2774}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ( Fresh[102] ), .c ({new_AGEMA_signal_1070, n2227}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2167 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2766}), .clk ( clk ), .r ( Fresh[103] ), .c ({new_AGEMA_signal_1009, n2027}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2171 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ( Fresh[104] ), .c ({new_AGEMA_signal_1167, n2214}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2173 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[105] ), .c ({new_AGEMA_signal_1168, n2290}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2174 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2758}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[106] ), .c ({new_AGEMA_signal_1169, n2376}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2178 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .r ( Fresh[107] ), .c ({new_AGEMA_signal_1072, n2034}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2182 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ( Fresh[108] ), .c ({new_AGEMA_signal_1073, n2171}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2183 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[109] ), .c ({new_AGEMA_signal_1170, n2039}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2188 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[110] ), .c ({new_AGEMA_signal_1172, n2042}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2191 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[111] ), .c ({new_AGEMA_signal_1173, n2754}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2192 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_959, n2790}), .clk ( clk ), .r ( Fresh[112] ), .c ({new_AGEMA_signal_1174, n2044}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2198 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .r ( Fresh[113] ), .c ({new_AGEMA_signal_1175, n2654}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2202 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1037, n2577}), .clk ( clk ), .r ( Fresh[114] ), .c ({new_AGEMA_signal_1176, n2055}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2205 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[115] ), .c ({new_AGEMA_signal_1177, n2057}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2208 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[116] ), .c ({new_AGEMA_signal_1178, n2407}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2212 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1010, n2061}), .clk ( clk ), .r ( Fresh[117] ), .c ({new_AGEMA_signal_1179, n2062}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2216 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ( Fresh[118] ), .c ({new_AGEMA_signal_1180, n2731}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2220 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1181, n2068}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2224 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ( Fresh[119] ), .c ({new_AGEMA_signal_1074, n2642}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2225 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ( Fresh[120] ), .c ({new_AGEMA_signal_1182, n2252}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2228 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ( Fresh[121] ), .c ({new_AGEMA_signal_1075, n2075}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) U2233 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ( Fresh[122] ), .c ({new_AGEMA_signal_1076, n2081}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2234 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[123] ), .c ({new_AGEMA_signal_1183, n2080}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2237 ( .a ({new_AGEMA_signal_984, n2600}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ( Fresh[124] ), .c ({new_AGEMA_signal_1077, n2498}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2238 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_1184, n2773}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2239 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[125] ), .c ({new_AGEMA_signal_1185, n2083}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2244 ( .a ({new_AGEMA_signal_2772, new_AGEMA_signal_2770}), .b ({new_AGEMA_signal_1033, n2086}), .clk ( clk ), .r ( Fresh[126] ), .c ({new_AGEMA_signal_1186, n2562}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2247 ( .a ({new_AGEMA_signal_2760, new_AGEMA_signal_2758}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ( Fresh[127] ), .c ({new_AGEMA_signal_1078, n2087}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2251 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1041, n2174}), .clk ( clk ), .r ( Fresh[128] ), .c ({new_AGEMA_signal_1187, n2156}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2260 ( .a ({new_AGEMA_signal_1028, n2769}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ( Fresh[129] ), .c ({new_AGEMA_signal_1188, n2100}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2277 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_1012, n2298}), .clk ( clk ), .r ( Fresh[130] ), .c ({new_AGEMA_signal_1079, n2544}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2279 ( .a ({new_AGEMA_signal_1004, n2356}), .b ({new_AGEMA_signal_1080, n2118}), .clk ( clk ), .r ( Fresh[131] ), .c ({new_AGEMA_signal_1191, n2121}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2284 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ( Fresh[132] ), .c ({new_AGEMA_signal_1193, n2122}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2286 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[133] ), .c ({new_AGEMA_signal_1194, n2811}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2294 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[134] ), .c ({new_AGEMA_signal_1081, n2647}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2297 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[135] ), .c ({new_AGEMA_signal_1082, n2132}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2304 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[136] ), .c ({new_AGEMA_signal_1199, n2220}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2305 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2746}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[137] ), .c ({new_AGEMA_signal_1200, n2138}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2312 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_2780, new_AGEMA_signal_2778}), .clk ( clk ), .r ( Fresh[138] ), .c ({new_AGEMA_signal_1201, n2555}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2322 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2782}), .clk ( clk ), .r ( Fresh[139] ), .c ({new_AGEMA_signal_1202, n2429}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2328 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2766}), .clk ( clk ), .r ( Fresh[140] ), .c ({new_AGEMA_signal_1083, n2162}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2337 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ( Fresh[141] ), .c ({new_AGEMA_signal_1014, n2545}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2340 ( .a ({new_AGEMA_signal_965, n2559}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[142] ), .c ({new_AGEMA_signal_1085, n2178}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2342 ( .a ({new_AGEMA_signal_1015, n2430}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[143] ), .c ({new_AGEMA_signal_1204, n2176}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2343 ( .a ({new_AGEMA_signal_1041, n2174}), .b ({new_AGEMA_signal_2772, new_AGEMA_signal_2770}), .clk ( clk ), .r ( Fresh[144] ), .c ({new_AGEMA_signal_1205, n2175}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2348 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2782}), .clk ( clk ), .r ( Fresh[145] ), .c ({new_AGEMA_signal_1016, n2182}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2353 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .r ( Fresh[146] ), .c ({new_AGEMA_signal_1206, n2188}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2355 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[147] ), .c ({new_AGEMA_signal_1207, n2189}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2357 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[148] ), .c ({new_AGEMA_signal_1208, n2446}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2362 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ( Fresh[149] ), .c ({new_AGEMA_signal_1087, n2576}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2363 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_2788, new_AGEMA_signal_2786}), .clk ( clk ), .r ( Fresh[150] ), .c ({new_AGEMA_signal_1088, n2748}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) U2368 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_1375, n2674}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2378 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[151] ), .c ({new_AGEMA_signal_1089, n2213}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2380 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_2760, new_AGEMA_signal_2758}), .clk ( clk ), .r ( Fresh[152] ), .c ({new_AGEMA_signal_1090, n2215}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2384 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[153] ), .c ({new_AGEMA_signal_1211, n2218}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2386 ( .a ({new_AGEMA_signal_1012, n2298}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[154] ), .c ({new_AGEMA_signal_1212, n2219}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2405 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[155] ), .c ({new_AGEMA_signal_1217, n2240}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2407 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ( Fresh[156] ), .c ({new_AGEMA_signal_1218, n2561}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2408 ( .a ({new_AGEMA_signal_2772, new_AGEMA_signal_2770}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ( Fresh[157] ), .c ({new_AGEMA_signal_1219, n2243}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2411 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ( Fresh[158] ), .c ({new_AGEMA_signal_1220, n2245}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2422 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .r ( Fresh[159] ), .c ({new_AGEMA_signal_1221, n2540}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2423 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ( Fresh[160] ), .c ({new_AGEMA_signal_1222, n2259}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2426 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ( Fresh[161] ), .c ({new_AGEMA_signal_1091, n2262}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2431 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[162] ), .c ({new_AGEMA_signal_1092, n2266}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2432 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_2784, new_AGEMA_signal_2782}), .clk ( clk ), .r ( Fresh[163] ), .c ({new_AGEMA_signal_1093, n2645}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2436 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2746}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ( Fresh[164] ), .c ({new_AGEMA_signal_1094, n2268}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2443 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ( Fresh[165] ), .c ({new_AGEMA_signal_1225, n2278}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2448 ( .a ({new_AGEMA_signal_2792, new_AGEMA_signal_2790}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[166] ), .c ({new_AGEMA_signal_1095, n2383}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2455 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ( Fresh[167] ), .c ({new_AGEMA_signal_1228, n2774}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2458 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[168] ), .c ({new_AGEMA_signal_1229, n2287}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2470 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[169] ), .c ({new_AGEMA_signal_1231, n2438}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2471 ( .a ({new_AGEMA_signal_1012, n2298}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[170] ), .c ({new_AGEMA_signal_1096, n2299}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2481 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1054, n2313}), .clk ( clk ), .r ( Fresh[171] ), .c ({new_AGEMA_signal_1232, n2371}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2484 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ( Fresh[172] ), .c ({new_AGEMA_signal_1018, n2316}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2486 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ( Fresh[173] ), .c ({new_AGEMA_signal_1098, n2318}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2492 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[174] ), .c ({new_AGEMA_signal_1235, n2325}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2494 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[175] ), .c ({new_AGEMA_signal_1236, n2328}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2495 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ( Fresh[176] ), .c ({new_AGEMA_signal_1099, n2327}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2505 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .r ( Fresh[177] ), .c ({new_AGEMA_signal_1237, n2343}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2510 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[178] ), .c ({new_AGEMA_signal_1239, n2344}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) U2512 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1013, n2346}), .clk ( clk ), .r ( Fresh[179] ), .c ({new_AGEMA_signal_1100, n2348}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2513 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ( Fresh[180] ), .c ({new_AGEMA_signal_1101, n2347}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2520 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ( Fresh[181] ), .c ({new_AGEMA_signal_1102, n2363}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2521 ( .a ({new_AGEMA_signal_1067, n2809}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2762}), .clk ( clk ), .r ( Fresh[182] ), .c ({new_AGEMA_signal_1243, n2353}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2524 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[183] ), .c ({new_AGEMA_signal_1244, n2355}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2530 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[184] ), .c ({new_AGEMA_signal_1245, n2364}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2543 ( .a ({new_AGEMA_signal_2748, new_AGEMA_signal_2746}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ( Fresh[185] ), .c ({new_AGEMA_signal_1103, n2415}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2558 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ( Fresh[186] ), .c ({new_AGEMA_signal_1104, n2700}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2563 ( .a ({new_AGEMA_signal_2796, new_AGEMA_signal_2794}), .b ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .r ( Fresh[187] ), .c ({new_AGEMA_signal_1105, n2594}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2564 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2766}), .clk ( clk ), .r ( Fresh[188] ), .c ({new_AGEMA_signal_1106, n2402}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2585 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ( Fresh[189] ), .c ({new_AGEMA_signal_1255, n2428}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2588 ( .a ({new_AGEMA_signal_1015, n2430}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ( Fresh[190] ), .c ({new_AGEMA_signal_1256, n2431}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2594 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[191] ), .c ({new_AGEMA_signal_1107, n2483}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2599 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[192] ), .c ({new_AGEMA_signal_1258, n2443}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2606 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[193] ), .c ({new_AGEMA_signal_1259, n2693}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2608 ( .a ({new_AGEMA_signal_998, n2452}), .b ({new_AGEMA_signal_2800, new_AGEMA_signal_2798}), .clk ( clk ), .r ( Fresh[194] ), .c ({new_AGEMA_signal_1108, n2453}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2616 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1019, n2463}), .clk ( clk ), .r ( Fresh[195] ), .c ({new_AGEMA_signal_1109, n2464}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2620 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[196] ), .c ({new_AGEMA_signal_1110, n2468}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2624 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2762}), .clk ( clk ), .r ( Fresh[197] ), .c ({new_AGEMA_signal_1111, n2473}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2625 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ( Fresh[198] ), .c ({new_AGEMA_signal_1112, n2472}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2628 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1020, n2474}), .clk ( clk ), .r ( Fresh[199] ), .c ({new_AGEMA_signal_1113, n2475}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2632 ( .a ({new_AGEMA_signal_2804, new_AGEMA_signal_2802}), .b ({new_AGEMA_signal_1065, n2828}), .clk ( clk ), .r ( Fresh[200] ), .c ({new_AGEMA_signal_1263, n2480}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2638 ( .a ({new_AGEMA_signal_1037, n2577}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[201] ), .c ({new_AGEMA_signal_1264, n2487}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2641 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ( Fresh[202] ), .c ({new_AGEMA_signal_1114, n2488}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2665 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ( Fresh[203] ), .c ({new_AGEMA_signal_1270, n2520}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2667 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_993, n2587}), .clk ( clk ), .r ( Fresh[204] ), .c ({new_AGEMA_signal_1115, n2521}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2674 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_963, n2595}), .clk ( clk ), .r ( Fresh[205] ), .c ({new_AGEMA_signal_1271, n2531}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2689 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ( Fresh[206] ), .c ({new_AGEMA_signal_1273, n2553}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2691 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[207] ), .c ({new_AGEMA_signal_1274, n2554}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) U2695 ( .a ({new_AGEMA_signal_965, n2559}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[208] ), .c ({new_AGEMA_signal_1116, n2560}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2698 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .r ( Fresh[209] ), .c ({new_AGEMA_signal_1275, n2564}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2714 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .r ( Fresh[210] ), .c ({new_AGEMA_signal_1278, n2586}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2720 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[211] ), .c ({new_AGEMA_signal_1117, n2597}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2721 ( .a ({new_AGEMA_signal_1024, n2640}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[212] ), .c ({new_AGEMA_signal_1280, n2596}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2723 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ( Fresh[213] ), .c ({new_AGEMA_signal_1281, n2598}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2725 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_2760, new_AGEMA_signal_2758}), .clk ( clk ), .r ( Fresh[214] ), .c ({new_AGEMA_signal_1021, n2599}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2732 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ( Fresh[215] ), .c ({new_AGEMA_signal_1283, n2610}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2734 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ( Fresh[216] ), .c ({new_AGEMA_signal_1284, n2614}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2735 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[217] ), .c ({new_AGEMA_signal_1285, n2613}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2737 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[218] ), .c ({new_AGEMA_signal_1119, n2617}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2742 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ( Fresh[219] ), .c ({new_AGEMA_signal_1120, n2629}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2751 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ( Fresh[220] ), .c ({new_AGEMA_signal_1287, n2784}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2757 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[221] ), .c ({new_AGEMA_signal_1121, n2650}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2775 ( .a ({new_AGEMA_signal_2780, new_AGEMA_signal_2778}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[222] ), .c ({new_AGEMA_signal_1022, n2683}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2789 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[223] ), .c ({new_AGEMA_signal_1294, n2711}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2790 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[224] ), .c ({new_AGEMA_signal_1295, n2710}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2792 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_969, n2712}), .clk ( clk ), .r ( Fresh[225] ), .c ({new_AGEMA_signal_1122, n2714}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2797 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1011, n2721}), .clk ( clk ), .r ( Fresh[226] ), .c ({new_AGEMA_signal_1123, n2722}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2799 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .r ( Fresh[227] ), .c ({new_AGEMA_signal_1297, n2726}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2806 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ( Fresh[228] ), .c ({new_AGEMA_signal_1298, n2738}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2822 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .r ( Fresh[229] ), .c ({new_AGEMA_signal_1301, n2768}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2828 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[230] ), .c ({new_AGEMA_signal_1124, n2782}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2829 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[231] ), .c ({new_AGEMA_signal_1125, n2781}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2832 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_989, n2785}), .clk ( clk ), .r ( Fresh[232] ), .c ({new_AGEMA_signal_1303, n2787}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2834 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[233] ), .c ({new_AGEMA_signal_1304, n2794}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2835 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_2792, new_AGEMA_signal_2790}), .clk ( clk ), .r ( Fresh[234] ), .c ({new_AGEMA_signal_1305, n2793}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2844 ( .a ({new_AGEMA_signal_2804, new_AGEMA_signal_2802}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ( Fresh[235] ), .c ({new_AGEMA_signal_1306, n2812}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2847 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ( Fresh[236] ), .c ({new_AGEMA_signal_1126, n2820}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2851 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ( Fresh[237] ), .c ({new_AGEMA_signal_1308, n2825}) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C ( clk ), .D ( new_AGEMA_signal_2805 ), .Q ( new_AGEMA_signal_2806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C ( clk ), .D ( new_AGEMA_signal_2807 ), .Q ( new_AGEMA_signal_2808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C ( clk ), .D ( new_AGEMA_signal_2809 ), .Q ( new_AGEMA_signal_2810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C ( clk ), .D ( new_AGEMA_signal_2811 ), .Q ( new_AGEMA_signal_2812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C ( clk ), .D ( new_AGEMA_signal_2813 ), .Q ( new_AGEMA_signal_2814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C ( clk ), .D ( new_AGEMA_signal_2815 ), .Q ( new_AGEMA_signal_2816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C ( clk ), .D ( new_AGEMA_signal_2817 ), .Q ( new_AGEMA_signal_2818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C ( clk ), .D ( new_AGEMA_signal_2819 ), .Q ( new_AGEMA_signal_2820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C ( clk ), .D ( new_AGEMA_signal_2821 ), .Q ( new_AGEMA_signal_2822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C ( clk ), .D ( new_AGEMA_signal_2823 ), .Q ( new_AGEMA_signal_2824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C ( clk ), .D ( new_AGEMA_signal_2825 ), .Q ( new_AGEMA_signal_2826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C ( clk ), .D ( new_AGEMA_signal_2827 ), .Q ( new_AGEMA_signal_2828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C ( clk ), .D ( new_AGEMA_signal_2829 ), .Q ( new_AGEMA_signal_2830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C ( clk ), .D ( new_AGEMA_signal_2831 ), .Q ( new_AGEMA_signal_2832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C ( clk ), .D ( new_AGEMA_signal_2833 ), .Q ( new_AGEMA_signal_2834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C ( clk ), .D ( new_AGEMA_signal_2835 ), .Q ( new_AGEMA_signal_2836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C ( clk ), .D ( new_AGEMA_signal_2837 ), .Q ( new_AGEMA_signal_2838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C ( clk ), .D ( new_AGEMA_signal_2839 ), .Q ( new_AGEMA_signal_2840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C ( clk ), .D ( new_AGEMA_signal_2841 ), .Q ( new_AGEMA_signal_2842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C ( clk ), .D ( new_AGEMA_signal_2843 ), .Q ( new_AGEMA_signal_2844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C ( clk ), .D ( new_AGEMA_signal_2845 ), .Q ( new_AGEMA_signal_2846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C ( clk ), .D ( new_AGEMA_signal_2847 ), .Q ( new_AGEMA_signal_2848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C ( clk ), .D ( new_AGEMA_signal_2849 ), .Q ( new_AGEMA_signal_2850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C ( clk ), .D ( new_AGEMA_signal_2851 ), .Q ( new_AGEMA_signal_2852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C ( clk ), .D ( new_AGEMA_signal_2853 ), .Q ( new_AGEMA_signal_2854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C ( clk ), .D ( new_AGEMA_signal_2855 ), .Q ( new_AGEMA_signal_2856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C ( clk ), .D ( new_AGEMA_signal_2857 ), .Q ( new_AGEMA_signal_2858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C ( clk ), .D ( new_AGEMA_signal_2859 ), .Q ( new_AGEMA_signal_2860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C ( clk ), .D ( new_AGEMA_signal_2861 ), .Q ( new_AGEMA_signal_2862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C ( clk ), .D ( new_AGEMA_signal_2863 ), .Q ( new_AGEMA_signal_2864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C ( clk ), .D ( new_AGEMA_signal_2865 ), .Q ( new_AGEMA_signal_2866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C ( clk ), .D ( new_AGEMA_signal_2867 ), .Q ( new_AGEMA_signal_2868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C ( clk ), .D ( new_AGEMA_signal_2869 ), .Q ( new_AGEMA_signal_2870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C ( clk ), .D ( new_AGEMA_signal_2871 ), .Q ( new_AGEMA_signal_2872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C ( clk ), .D ( new_AGEMA_signal_2873 ), .Q ( new_AGEMA_signal_2874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C ( clk ), .D ( new_AGEMA_signal_2875 ), .Q ( new_AGEMA_signal_2876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C ( clk ), .D ( new_AGEMA_signal_2877 ), .Q ( new_AGEMA_signal_2878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C ( clk ), .D ( new_AGEMA_signal_2879 ), .Q ( new_AGEMA_signal_2880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C ( clk ), .D ( new_AGEMA_signal_2881 ), .Q ( new_AGEMA_signal_2882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C ( clk ), .D ( new_AGEMA_signal_2883 ), .Q ( new_AGEMA_signal_2884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C ( clk ), .D ( new_AGEMA_signal_2885 ), .Q ( new_AGEMA_signal_2886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C ( clk ), .D ( new_AGEMA_signal_2887 ), .Q ( new_AGEMA_signal_2888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C ( clk ), .D ( new_AGEMA_signal_2889 ), .Q ( new_AGEMA_signal_2890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C ( clk ), .D ( new_AGEMA_signal_2891 ), .Q ( new_AGEMA_signal_2892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C ( clk ), .D ( new_AGEMA_signal_2893 ), .Q ( new_AGEMA_signal_2894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C ( clk ), .D ( new_AGEMA_signal_2895 ), .Q ( new_AGEMA_signal_2896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C ( clk ), .D ( new_AGEMA_signal_2897 ), .Q ( new_AGEMA_signal_2898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C ( clk ), .D ( new_AGEMA_signal_2899 ), .Q ( new_AGEMA_signal_2900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C ( clk ), .D ( new_AGEMA_signal_2901 ), .Q ( new_AGEMA_signal_2902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C ( clk ), .D ( new_AGEMA_signal_2903 ), .Q ( new_AGEMA_signal_2904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C ( clk ), .D ( new_AGEMA_signal_2905 ), .Q ( new_AGEMA_signal_2906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C ( clk ), .D ( new_AGEMA_signal_2907 ), .Q ( new_AGEMA_signal_2908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C ( clk ), .D ( new_AGEMA_signal_2909 ), .Q ( new_AGEMA_signal_2910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C ( clk ), .D ( new_AGEMA_signal_2911 ), .Q ( new_AGEMA_signal_2912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C ( clk ), .D ( new_AGEMA_signal_2913 ), .Q ( new_AGEMA_signal_2914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C ( clk ), .D ( new_AGEMA_signal_2915 ), .Q ( new_AGEMA_signal_2916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C ( clk ), .D ( new_AGEMA_signal_2917 ), .Q ( new_AGEMA_signal_2918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C ( clk ), .D ( new_AGEMA_signal_2919 ), .Q ( new_AGEMA_signal_2920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C ( clk ), .D ( new_AGEMA_signal_2921 ), .Q ( new_AGEMA_signal_2922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C ( clk ), .D ( new_AGEMA_signal_2923 ), .Q ( new_AGEMA_signal_2924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C ( clk ), .D ( new_AGEMA_signal_2925 ), .Q ( new_AGEMA_signal_2926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C ( clk ), .D ( new_AGEMA_signal_2927 ), .Q ( new_AGEMA_signal_2928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C ( clk ), .D ( new_AGEMA_signal_2929 ), .Q ( new_AGEMA_signal_2930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C ( clk ), .D ( new_AGEMA_signal_2931 ), .Q ( new_AGEMA_signal_2932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C ( clk ), .D ( new_AGEMA_signal_2933 ), .Q ( new_AGEMA_signal_2934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C ( clk ), .D ( new_AGEMA_signal_2935 ), .Q ( new_AGEMA_signal_2936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C ( clk ), .D ( new_AGEMA_signal_2937 ), .Q ( new_AGEMA_signal_2938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C ( clk ), .D ( new_AGEMA_signal_2939 ), .Q ( new_AGEMA_signal_2940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C ( clk ), .D ( new_AGEMA_signal_2941 ), .Q ( new_AGEMA_signal_2942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C ( clk ), .D ( new_AGEMA_signal_2943 ), .Q ( new_AGEMA_signal_2944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C ( clk ), .D ( new_AGEMA_signal_2945 ), .Q ( new_AGEMA_signal_2946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C ( clk ), .D ( new_AGEMA_signal_2947 ), .Q ( new_AGEMA_signal_2948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C ( clk ), .D ( new_AGEMA_signal_2949 ), .Q ( new_AGEMA_signal_2950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C ( clk ), .D ( new_AGEMA_signal_2951 ), .Q ( new_AGEMA_signal_2952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C ( clk ), .D ( new_AGEMA_signal_2953 ), .Q ( new_AGEMA_signal_2954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C ( clk ), .D ( new_AGEMA_signal_2955 ), .Q ( new_AGEMA_signal_2956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C ( clk ), .D ( new_AGEMA_signal_2957 ), .Q ( new_AGEMA_signal_2958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C ( clk ), .D ( new_AGEMA_signal_2959 ), .Q ( new_AGEMA_signal_2960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C ( clk ), .D ( new_AGEMA_signal_2961 ), .Q ( new_AGEMA_signal_2962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C ( clk ), .D ( new_AGEMA_signal_2963 ), .Q ( new_AGEMA_signal_2964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C ( clk ), .D ( new_AGEMA_signal_2965 ), .Q ( new_AGEMA_signal_2966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C ( clk ), .D ( new_AGEMA_signal_2967 ), .Q ( new_AGEMA_signal_2968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C ( clk ), .D ( new_AGEMA_signal_2969 ), .Q ( new_AGEMA_signal_2970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C ( clk ), .D ( new_AGEMA_signal_2971 ), .Q ( new_AGEMA_signal_2972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C ( clk ), .D ( new_AGEMA_signal_2973 ), .Q ( new_AGEMA_signal_2974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C ( clk ), .D ( new_AGEMA_signal_2975 ), .Q ( new_AGEMA_signal_2976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C ( clk ), .D ( new_AGEMA_signal_2977 ), .Q ( new_AGEMA_signal_2978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C ( clk ), .D ( new_AGEMA_signal_2979 ), .Q ( new_AGEMA_signal_2980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C ( clk ), .D ( new_AGEMA_signal_2981 ), .Q ( new_AGEMA_signal_2982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C ( clk ), .D ( new_AGEMA_signal_2983 ), .Q ( new_AGEMA_signal_2984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C ( clk ), .D ( new_AGEMA_signal_2985 ), .Q ( new_AGEMA_signal_2986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C ( clk ), .D ( new_AGEMA_signal_2987 ), .Q ( new_AGEMA_signal_2988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C ( clk ), .D ( new_AGEMA_signal_2989 ), .Q ( new_AGEMA_signal_2990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C ( clk ), .D ( new_AGEMA_signal_2991 ), .Q ( new_AGEMA_signal_2992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C ( clk ), .D ( new_AGEMA_signal_2993 ), .Q ( new_AGEMA_signal_2994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C ( clk ), .D ( new_AGEMA_signal_2995 ), .Q ( new_AGEMA_signal_2996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C ( clk ), .D ( new_AGEMA_signal_2997 ), .Q ( new_AGEMA_signal_2998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C ( clk ), .D ( new_AGEMA_signal_2999 ), .Q ( new_AGEMA_signal_3000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C ( clk ), .D ( new_AGEMA_signal_3001 ), .Q ( new_AGEMA_signal_3002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C ( clk ), .D ( new_AGEMA_signal_3003 ), .Q ( new_AGEMA_signal_3004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C ( clk ), .D ( new_AGEMA_signal_3005 ), .Q ( new_AGEMA_signal_3006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C ( clk ), .D ( new_AGEMA_signal_3007 ), .Q ( new_AGEMA_signal_3008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C ( clk ), .D ( new_AGEMA_signal_3009 ), .Q ( new_AGEMA_signal_3010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C ( clk ), .D ( new_AGEMA_signal_3011 ), .Q ( new_AGEMA_signal_3012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C ( clk ), .D ( new_AGEMA_signal_3013 ), .Q ( new_AGEMA_signal_3014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C ( clk ), .D ( new_AGEMA_signal_3015 ), .Q ( new_AGEMA_signal_3016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C ( clk ), .D ( new_AGEMA_signal_3017 ), .Q ( new_AGEMA_signal_3018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C ( clk ), .D ( new_AGEMA_signal_3019 ), .Q ( new_AGEMA_signal_3020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C ( clk ), .D ( new_AGEMA_signal_3021 ), .Q ( new_AGEMA_signal_3022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C ( clk ), .D ( new_AGEMA_signal_3023 ), .Q ( new_AGEMA_signal_3024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C ( clk ), .D ( new_AGEMA_signal_3025 ), .Q ( new_AGEMA_signal_3026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C ( clk ), .D ( new_AGEMA_signal_3027 ), .Q ( new_AGEMA_signal_3028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C ( clk ), .D ( new_AGEMA_signal_3029 ), .Q ( new_AGEMA_signal_3030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C ( clk ), .D ( new_AGEMA_signal_3031 ), .Q ( new_AGEMA_signal_3032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C ( clk ), .D ( new_AGEMA_signal_3033 ), .Q ( new_AGEMA_signal_3034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C ( clk ), .D ( new_AGEMA_signal_3035 ), .Q ( new_AGEMA_signal_3036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C ( clk ), .D ( new_AGEMA_signal_3037 ), .Q ( new_AGEMA_signal_3038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C ( clk ), .D ( new_AGEMA_signal_3039 ), .Q ( new_AGEMA_signal_3040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C ( clk ), .D ( new_AGEMA_signal_3041 ), .Q ( new_AGEMA_signal_3042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C ( clk ), .D ( new_AGEMA_signal_3043 ), .Q ( new_AGEMA_signal_3044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C ( clk ), .D ( new_AGEMA_signal_3045 ), .Q ( new_AGEMA_signal_3046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C ( clk ), .D ( new_AGEMA_signal_3047 ), .Q ( new_AGEMA_signal_3048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C ( clk ), .D ( new_AGEMA_signal_3049 ), .Q ( new_AGEMA_signal_3050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C ( clk ), .D ( new_AGEMA_signal_3051 ), .Q ( new_AGEMA_signal_3052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C ( clk ), .D ( new_AGEMA_signal_3053 ), .Q ( new_AGEMA_signal_3054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C ( clk ), .D ( new_AGEMA_signal_3055 ), .Q ( new_AGEMA_signal_3056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C ( clk ), .D ( new_AGEMA_signal_3057 ), .Q ( new_AGEMA_signal_3058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C ( clk ), .D ( new_AGEMA_signal_3059 ), .Q ( new_AGEMA_signal_3060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C ( clk ), .D ( new_AGEMA_signal_3061 ), .Q ( new_AGEMA_signal_3062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C ( clk ), .D ( new_AGEMA_signal_3063 ), .Q ( new_AGEMA_signal_3064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C ( clk ), .D ( new_AGEMA_signal_3065 ), .Q ( new_AGEMA_signal_3066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C ( clk ), .D ( new_AGEMA_signal_3067 ), .Q ( new_AGEMA_signal_3068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C ( clk ), .D ( new_AGEMA_signal_3069 ), .Q ( new_AGEMA_signal_3070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C ( clk ), .D ( new_AGEMA_signal_3071 ), .Q ( new_AGEMA_signal_3072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C ( clk ), .D ( new_AGEMA_signal_3073 ), .Q ( new_AGEMA_signal_3074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C ( clk ), .D ( new_AGEMA_signal_3075 ), .Q ( new_AGEMA_signal_3076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C ( clk ), .D ( new_AGEMA_signal_3085 ), .Q ( new_AGEMA_signal_3086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C ( clk ), .D ( new_AGEMA_signal_3089 ), .Q ( new_AGEMA_signal_3090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C ( clk ), .D ( new_AGEMA_signal_3137 ), .Q ( new_AGEMA_signal_3138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C ( clk ), .D ( new_AGEMA_signal_3141 ), .Q ( new_AGEMA_signal_3142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C ( clk ), .D ( new_AGEMA_signal_3173 ), .Q ( new_AGEMA_signal_3174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C ( clk ), .D ( new_AGEMA_signal_3177 ), .Q ( new_AGEMA_signal_3178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C ( clk ), .D ( new_AGEMA_signal_3201 ), .Q ( new_AGEMA_signal_3202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C ( clk ), .D ( new_AGEMA_signal_3205 ), .Q ( new_AGEMA_signal_3206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C ( clk ), .D ( new_AGEMA_signal_3221 ), .Q ( new_AGEMA_signal_3222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C ( clk ), .D ( new_AGEMA_signal_3225 ), .Q ( new_AGEMA_signal_3226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C ( clk ), .D ( new_AGEMA_signal_3241 ), .Q ( new_AGEMA_signal_3242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C ( clk ), .D ( new_AGEMA_signal_3245 ), .Q ( new_AGEMA_signal_3246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C ( clk ), .D ( new_AGEMA_signal_3319 ), .Q ( new_AGEMA_signal_3320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C ( clk ), .D ( new_AGEMA_signal_3325 ), .Q ( new_AGEMA_signal_3326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C ( clk ), .D ( new_AGEMA_signal_3341 ), .Q ( new_AGEMA_signal_3342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C ( clk ), .D ( new_AGEMA_signal_3345 ), .Q ( new_AGEMA_signal_3346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C ( clk ), .D ( new_AGEMA_signal_3361 ), .Q ( new_AGEMA_signal_3362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C ( clk ), .D ( new_AGEMA_signal_3365 ), .Q ( new_AGEMA_signal_3366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C ( clk ), .D ( new_AGEMA_signal_3397 ), .Q ( new_AGEMA_signal_3398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C ( clk ), .D ( new_AGEMA_signal_3401 ), .Q ( new_AGEMA_signal_3402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C ( clk ), .D ( new_AGEMA_signal_3413 ), .Q ( new_AGEMA_signal_3414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C ( clk ), .D ( new_AGEMA_signal_3417 ), .Q ( new_AGEMA_signal_3418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C ( clk ), .D ( new_AGEMA_signal_3561 ), .Q ( new_AGEMA_signal_3562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C ( clk ), .D ( new_AGEMA_signal_3567 ), .Q ( new_AGEMA_signal_3568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C ( clk ), .D ( new_AGEMA_signal_3613 ), .Q ( new_AGEMA_signal_3614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C ( clk ), .D ( new_AGEMA_signal_3619 ), .Q ( new_AGEMA_signal_3620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C ( clk ), .D ( new_AGEMA_signal_3845 ), .Q ( new_AGEMA_signal_3846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C ( clk ), .D ( new_AGEMA_signal_3853 ), .Q ( new_AGEMA_signal_3854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C ( clk ), .D ( new_AGEMA_signal_3865 ), .Q ( new_AGEMA_signal_3866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C ( clk ), .D ( new_AGEMA_signal_3873 ), .Q ( new_AGEMA_signal_3874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C ( clk ), .D ( new_AGEMA_signal_4017 ), .Q ( new_AGEMA_signal_4018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C ( clk ), .D ( new_AGEMA_signal_4025 ), .Q ( new_AGEMA_signal_4026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C ( clk ), .D ( new_AGEMA_signal_4189 ), .Q ( new_AGEMA_signal_4190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C ( clk ), .D ( new_AGEMA_signal_4197 ), .Q ( new_AGEMA_signal_4198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C ( clk ), .D ( new_AGEMA_signal_4249 ), .Q ( new_AGEMA_signal_4250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C ( clk ), .D ( new_AGEMA_signal_4257 ), .Q ( new_AGEMA_signal_4258 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1259 ( .C ( clk ), .D ( n2755 ), .Q ( new_AGEMA_signal_3077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_3079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C ( clk ), .D ( n2151 ), .Q ( new_AGEMA_signal_3081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C ( clk ), .D ( new_AGEMA_signal_1132 ), .Q ( new_AGEMA_signal_3083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C ( clk ), .D ( new_AGEMA_signal_3086 ), .Q ( new_AGEMA_signal_3087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C ( clk ), .D ( new_AGEMA_signal_3090 ), .Q ( new_AGEMA_signal_3091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C ( clk ), .D ( new_AGEMA_signal_2838 ), .Q ( new_AGEMA_signal_3093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C ( clk ), .D ( new_AGEMA_signal_2840 ), .Q ( new_AGEMA_signal_3095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C ( clk ), .D ( new_AGEMA_signal_2826 ), .Q ( new_AGEMA_signal_3097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C ( clk ), .D ( new_AGEMA_signal_2828 ), .Q ( new_AGEMA_signal_3099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C ( clk ), .D ( n1964 ), .Q ( new_AGEMA_signal_3101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C ( clk ), .D ( new_AGEMA_signal_999 ), .Q ( new_AGEMA_signal_3103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C ( clk ), .D ( n2673 ), .Q ( new_AGEMA_signal_3105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C ( clk ), .D ( new_AGEMA_signal_1052 ), .Q ( new_AGEMA_signal_3107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C ( clk ), .D ( n2359 ), .Q ( new_AGEMA_signal_3109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C ( clk ), .D ( new_AGEMA_signal_1147 ), .Q ( new_AGEMA_signal_3111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C ( clk ), .D ( n1973 ), .Q ( new_AGEMA_signal_3113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C ( clk ), .D ( new_AGEMA_signal_1151 ), .Q ( new_AGEMA_signal_3115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C ( clk ), .D ( n2690 ), .Q ( new_AGEMA_signal_3117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_3119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C ( clk ), .D ( n2741 ), .Q ( new_AGEMA_signal_3121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C ( clk ), .D ( new_AGEMA_signal_1153 ), .Q ( new_AGEMA_signal_3123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C ( clk ), .D ( n1993 ), .Q ( new_AGEMA_signal_3125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_3127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C ( clk ), .D ( n2241 ), .Q ( new_AGEMA_signal_3129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C ( clk ), .D ( new_AGEMA_signal_1157 ), .Q ( new_AGEMA_signal_3131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C ( clk ), .D ( new_AGEMA_signal_2946 ), .Q ( new_AGEMA_signal_3133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C ( clk ), .D ( new_AGEMA_signal_2948 ), .Q ( new_AGEMA_signal_3135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C ( clk ), .D ( new_AGEMA_signal_3138 ), .Q ( new_AGEMA_signal_3139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C ( clk ), .D ( new_AGEMA_signal_3142 ), .Q ( new_AGEMA_signal_3143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C ( clk ), .D ( n2290 ), .Q ( new_AGEMA_signal_3145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C ( clk ), .D ( new_AGEMA_signal_1168 ), .Q ( new_AGEMA_signal_3147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C ( clk ), .D ( n2171 ), .Q ( new_AGEMA_signal_3149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_3151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C ( clk ), .D ( n2042 ), .Q ( new_AGEMA_signal_3153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C ( clk ), .D ( new_AGEMA_signal_1172 ), .Q ( new_AGEMA_signal_3155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C ( clk ), .D ( n2754 ), .Q ( new_AGEMA_signal_3157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C ( clk ), .D ( new_AGEMA_signal_1173 ), .Q ( new_AGEMA_signal_3159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C ( clk ), .D ( new_AGEMA_signal_2806 ), .Q ( new_AGEMA_signal_3161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C ( clk ), .D ( new_AGEMA_signal_2808 ), .Q ( new_AGEMA_signal_3163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C ( clk ), .D ( n2535 ), .Q ( new_AGEMA_signal_3165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C ( clk ), .D ( new_AGEMA_signal_1150 ), .Q ( new_AGEMA_signal_3167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C ( clk ), .D ( n2642 ), .Q ( new_AGEMA_signal_3169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_3171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C ( clk ), .D ( new_AGEMA_signal_3174 ), .Q ( new_AGEMA_signal_3175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C ( clk ), .D ( new_AGEMA_signal_3178 ), .Q ( new_AGEMA_signal_3179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C ( clk ), .D ( n2773 ), .Q ( new_AGEMA_signal_3181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C ( clk ), .D ( new_AGEMA_signal_1184 ), .Q ( new_AGEMA_signal_3183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C ( clk ), .D ( n2627 ), .Q ( new_AGEMA_signal_3185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C ( clk ), .D ( new_AGEMA_signal_1048 ), .Q ( new_AGEMA_signal_3187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C ( clk ), .D ( new_AGEMA_signal_2886 ), .Q ( new_AGEMA_signal_3189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C ( clk ), .D ( new_AGEMA_signal_2888 ), .Q ( new_AGEMA_signal_3191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C ( clk ), .D ( n2631 ), .Q ( new_AGEMA_signal_3193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C ( clk ), .D ( new_AGEMA_signal_1034 ), .Q ( new_AGEMA_signal_3195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C ( clk ), .D ( n2376 ), .Q ( new_AGEMA_signal_3197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C ( clk ), .D ( new_AGEMA_signal_1169 ), .Q ( new_AGEMA_signal_3199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C ( clk ), .D ( new_AGEMA_signal_3202 ), .Q ( new_AGEMA_signal_3203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C ( clk ), .D ( new_AGEMA_signal_3206 ), .Q ( new_AGEMA_signal_3207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C ( clk ), .D ( new_AGEMA_signal_2978 ), .Q ( new_AGEMA_signal_3209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C ( clk ), .D ( new_AGEMA_signal_2980 ), .Q ( new_AGEMA_signal_3211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C ( clk ), .D ( new_AGEMA_signal_2906 ), .Q ( new_AGEMA_signal_3213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C ( clk ), .D ( new_AGEMA_signal_2908 ), .Q ( new_AGEMA_signal_3215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C ( clk ), .D ( new_AGEMA_signal_2922 ), .Q ( new_AGEMA_signal_3217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C ( clk ), .D ( new_AGEMA_signal_2924 ), .Q ( new_AGEMA_signal_3219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C ( clk ), .D ( new_AGEMA_signal_3222 ), .Q ( new_AGEMA_signal_3223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C ( clk ), .D ( new_AGEMA_signal_3226 ), .Q ( new_AGEMA_signal_3227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C ( clk ), .D ( new_AGEMA_signal_3058 ), .Q ( new_AGEMA_signal_3229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C ( clk ), .D ( new_AGEMA_signal_3060 ), .Q ( new_AGEMA_signal_3231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C ( clk ), .D ( n2498 ), .Q ( new_AGEMA_signal_3233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C ( clk ), .D ( new_AGEMA_signal_1077 ), .Q ( new_AGEMA_signal_3235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C ( clk ), .D ( n2178 ), .Q ( new_AGEMA_signal_3237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_3239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C ( clk ), .D ( new_AGEMA_signal_3242 ), .Q ( new_AGEMA_signal_3243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C ( clk ), .D ( new_AGEMA_signal_3246 ), .Q ( new_AGEMA_signal_3247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C ( clk ), .D ( n2505 ), .Q ( new_AGEMA_signal_3249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C ( clk ), .D ( new_AGEMA_signal_1146 ), .Q ( new_AGEMA_signal_3251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C ( clk ), .D ( n2540 ), .Q ( new_AGEMA_signal_3253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C ( clk ), .D ( new_AGEMA_signal_1221 ), .Q ( new_AGEMA_signal_3255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C ( clk ), .D ( n2266 ), .Q ( new_AGEMA_signal_3257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_3259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C ( clk ), .D ( n2278 ), .Q ( new_AGEMA_signal_3261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C ( clk ), .D ( new_AGEMA_signal_1225 ), .Q ( new_AGEMA_signal_3263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C ( clk ), .D ( new_AGEMA_signal_2970 ), .Q ( new_AGEMA_signal_3265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C ( clk ), .D ( new_AGEMA_signal_2972 ), .Q ( new_AGEMA_signal_3267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C ( clk ), .D ( new_AGEMA_signal_3014 ), .Q ( new_AGEMA_signal_3269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C ( clk ), .D ( new_AGEMA_signal_3016 ), .Q ( new_AGEMA_signal_3271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C ( clk ), .D ( new_AGEMA_signal_2878 ), .Q ( new_AGEMA_signal_3273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C ( clk ), .D ( new_AGEMA_signal_2880 ), .Q ( new_AGEMA_signal_3275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C ( clk ), .D ( new_AGEMA_signal_2870 ), .Q ( new_AGEMA_signal_3277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C ( clk ), .D ( new_AGEMA_signal_2872 ), .Q ( new_AGEMA_signal_3279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C ( clk ), .D ( n2318 ), .Q ( new_AGEMA_signal_3281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C ( clk ), .D ( new_AGEMA_signal_1098 ), .Q ( new_AGEMA_signal_3283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C ( clk ), .D ( n2325 ), .Q ( new_AGEMA_signal_3285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C ( clk ), .D ( new_AGEMA_signal_1235 ), .Q ( new_AGEMA_signal_3287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C ( clk ), .D ( n2677 ), .Q ( new_AGEMA_signal_3289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C ( clk ), .D ( new_AGEMA_signal_1047 ), .Q ( new_AGEMA_signal_3291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C ( clk ), .D ( new_AGEMA_signal_3050 ), .Q ( new_AGEMA_signal_3293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C ( clk ), .D ( new_AGEMA_signal_3052 ), .Q ( new_AGEMA_signal_3295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C ( clk ), .D ( new_AGEMA_signal_3066 ), .Q ( new_AGEMA_signal_3297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C ( clk ), .D ( new_AGEMA_signal_3068 ), .Q ( new_AGEMA_signal_3299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C ( clk ), .D ( new_AGEMA_signal_2914 ), .Q ( new_AGEMA_signal_3301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C ( clk ), .D ( new_AGEMA_signal_2916 ), .Q ( new_AGEMA_signal_3303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C ( clk ), .D ( new_AGEMA_signal_2814 ), .Q ( new_AGEMA_signal_3305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C ( clk ), .D ( new_AGEMA_signal_2816 ), .Q ( new_AGEMA_signal_3307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C ( clk ), .D ( n2625 ), .Q ( new_AGEMA_signal_3309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C ( clk ), .D ( new_AGEMA_signal_1148 ), .Q ( new_AGEMA_signal_3311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C ( clk ), .D ( n2431 ), .Q ( new_AGEMA_signal_3313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C ( clk ), .D ( new_AGEMA_signal_1256 ), .Q ( new_AGEMA_signal_3315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C ( clk ), .D ( new_AGEMA_signal_3320 ), .Q ( new_AGEMA_signal_3321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C ( clk ), .D ( new_AGEMA_signal_3326 ), .Q ( new_AGEMA_signal_3327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C ( clk ), .D ( n2453 ), .Q ( new_AGEMA_signal_3329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_3331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C ( clk ), .D ( n2475 ), .Q ( new_AGEMA_signal_3333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C ( clk ), .D ( new_AGEMA_signal_1113 ), .Q ( new_AGEMA_signal_3335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C ( clk ), .D ( n2487 ), .Q ( new_AGEMA_signal_3337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C ( clk ), .D ( new_AGEMA_signal_1264 ), .Q ( new_AGEMA_signal_3339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C ( clk ), .D ( new_AGEMA_signal_3342 ), .Q ( new_AGEMA_signal_3343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C ( clk ), .D ( new_AGEMA_signal_3346 ), .Q ( new_AGEMA_signal_3347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C ( clk ), .D ( new_AGEMA_signal_2954 ), .Q ( new_AGEMA_signal_3349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C ( clk ), .D ( new_AGEMA_signal_2956 ), .Q ( new_AGEMA_signal_3351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C ( clk ), .D ( new_AGEMA_signal_2962 ), .Q ( new_AGEMA_signal_3353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C ( clk ), .D ( new_AGEMA_signal_2964 ), .Q ( new_AGEMA_signal_3355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C ( clk ), .D ( n2564 ), .Q ( new_AGEMA_signal_3357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C ( clk ), .D ( new_AGEMA_signal_1275 ), .Q ( new_AGEMA_signal_3359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C ( clk ), .D ( new_AGEMA_signal_3362 ), .Q ( new_AGEMA_signal_3363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C ( clk ), .D ( new_AGEMA_signal_3366 ), .Q ( new_AGEMA_signal_3367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C ( clk ), .D ( n2617 ), .Q ( new_AGEMA_signal_3369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C ( clk ), .D ( new_AGEMA_signal_1119 ), .Q ( new_AGEMA_signal_3371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C ( clk ), .D ( n2647 ), .Q ( new_AGEMA_signal_3373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_3375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C ( clk ), .D ( n2674 ), .Q ( new_AGEMA_signal_3377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C ( clk ), .D ( new_AGEMA_signal_1375 ), .Q ( new_AGEMA_signal_3379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C ( clk ), .D ( n2683 ), .Q ( new_AGEMA_signal_3381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C ( clk ), .D ( new_AGEMA_signal_1022 ), .Q ( new_AGEMA_signal_3383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C ( clk ), .D ( n2714 ), .Q ( new_AGEMA_signal_3385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C ( clk ), .D ( new_AGEMA_signal_1122 ), .Q ( new_AGEMA_signal_3387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C ( clk ), .D ( n2726 ), .Q ( new_AGEMA_signal_3389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C ( clk ), .D ( new_AGEMA_signal_1297 ), .Q ( new_AGEMA_signal_3391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C ( clk ), .D ( n2734 ), .Q ( new_AGEMA_signal_3393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C ( clk ), .D ( new_AGEMA_signal_1133 ), .Q ( new_AGEMA_signal_3395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C ( clk ), .D ( new_AGEMA_signal_3398 ), .Q ( new_AGEMA_signal_3399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C ( clk ), .D ( new_AGEMA_signal_3402 ), .Q ( new_AGEMA_signal_3403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C ( clk ), .D ( n2763 ), .Q ( new_AGEMA_signal_3405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C ( clk ), .D ( new_AGEMA_signal_1134 ), .Q ( new_AGEMA_signal_3407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C ( clk ), .D ( n2784 ), .Q ( new_AGEMA_signal_3409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C ( clk ), .D ( new_AGEMA_signal_1287 ), .Q ( new_AGEMA_signal_3411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C ( clk ), .D ( new_AGEMA_signal_3414 ), .Q ( new_AGEMA_signal_3415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C ( clk ), .D ( new_AGEMA_signal_3418 ), .Q ( new_AGEMA_signal_3419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C ( clk ), .D ( n2820 ), .Q ( new_AGEMA_signal_3421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C ( clk ), .D ( new_AGEMA_signal_1126 ), .Q ( new_AGEMA_signal_3423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C ( clk ), .D ( new_AGEMA_signal_3042 ), .Q ( new_AGEMA_signal_3425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C ( clk ), .D ( new_AGEMA_signal_3044 ), .Q ( new_AGEMA_signal_3429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C ( clk ), .D ( n1930 ), .Q ( new_AGEMA_signal_3433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C ( clk ), .D ( new_AGEMA_signal_1036 ), .Q ( new_AGEMA_signal_3437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C ( clk ), .D ( n1976 ), .Q ( new_AGEMA_signal_3449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_3453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C ( clk ), .D ( new_AGEMA_signal_2874 ), .Q ( new_AGEMA_signal_3461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C ( clk ), .D ( new_AGEMA_signal_2876 ), .Q ( new_AGEMA_signal_3465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C ( clk ), .D ( n2008 ), .Q ( new_AGEMA_signal_3473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C ( clk ), .D ( new_AGEMA_signal_1159 ), .Q ( new_AGEMA_signal_3477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C ( clk ), .D ( n2022 ), .Q ( new_AGEMA_signal_3481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C ( clk ), .D ( new_AGEMA_signal_1164 ), .Q ( new_AGEMA_signal_3485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C ( clk ), .D ( n2057 ), .Q ( new_AGEMA_signal_3505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C ( clk ), .D ( new_AGEMA_signal_1177 ), .Q ( new_AGEMA_signal_3509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C ( clk ), .D ( n2062 ), .Q ( new_AGEMA_signal_3513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C ( clk ), .D ( new_AGEMA_signal_1179 ), .Q ( new_AGEMA_signal_3517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C ( clk ), .D ( n2075 ), .Q ( new_AGEMA_signal_3521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_3525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C ( clk ), .D ( n2121 ), .Q ( new_AGEMA_signal_3541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C ( clk ), .D ( new_AGEMA_signal_1191 ), .Q ( new_AGEMA_signal_3545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C ( clk ), .D ( new_AGEMA_signal_2854 ), .Q ( new_AGEMA_signal_3553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C ( clk ), .D ( new_AGEMA_signal_2856 ), .Q ( new_AGEMA_signal_3557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C ( clk ), .D ( new_AGEMA_signal_3562 ), .Q ( new_AGEMA_signal_3563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C ( clk ), .D ( new_AGEMA_signal_3568 ), .Q ( new_AGEMA_signal_3569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C ( clk ), .D ( new_AGEMA_signal_2998 ), .Q ( new_AGEMA_signal_3573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C ( clk ), .D ( new_AGEMA_signal_3000 ), .Q ( new_AGEMA_signal_3577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C ( clk ), .D ( new_AGEMA_signal_3026 ), .Q ( new_AGEMA_signal_3581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C ( clk ), .D ( new_AGEMA_signal_3028 ), .Q ( new_AGEMA_signal_3585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C ( clk ), .D ( n2245 ), .Q ( new_AGEMA_signal_3605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C ( clk ), .D ( new_AGEMA_signal_1220 ), .Q ( new_AGEMA_signal_3609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C ( clk ), .D ( new_AGEMA_signal_3614 ), .Q ( new_AGEMA_signal_3615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C ( clk ), .D ( new_AGEMA_signal_3620 ), .Q ( new_AGEMA_signal_3621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C ( clk ), .D ( n2262 ), .Q ( new_AGEMA_signal_3625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C ( clk ), .D ( new_AGEMA_signal_1091 ), .Q ( new_AGEMA_signal_3629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C ( clk ), .D ( n2343 ), .Q ( new_AGEMA_signal_3645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C ( clk ), .D ( new_AGEMA_signal_1237 ), .Q ( new_AGEMA_signal_3649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C ( clk ), .D ( new_AGEMA_signal_3002 ), .Q ( new_AGEMA_signal_3661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C ( clk ), .D ( new_AGEMA_signal_3004 ), .Q ( new_AGEMA_signal_3665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C ( clk ), .D ( new_AGEMA_signal_2986 ), .Q ( new_AGEMA_signal_3669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C ( clk ), .D ( new_AGEMA_signal_2988 ), .Q ( new_AGEMA_signal_3673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C ( clk ), .D ( new_AGEMA_signal_2846 ), .Q ( new_AGEMA_signal_3677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C ( clk ), .D ( new_AGEMA_signal_2848 ), .Q ( new_AGEMA_signal_3681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C ( clk ), .D ( new_AGEMA_signal_2898 ), .Q ( new_AGEMA_signal_3685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C ( clk ), .D ( new_AGEMA_signal_2900 ), .Q ( new_AGEMA_signal_3689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C ( clk ), .D ( n2417 ), .Q ( new_AGEMA_signal_3693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C ( clk ), .D ( new_AGEMA_signal_1324 ), .Q ( new_AGEMA_signal_3697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C ( clk ), .D ( new_AGEMA_signal_3038 ), .Q ( new_AGEMA_signal_3717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C ( clk ), .D ( new_AGEMA_signal_3040 ), .Q ( new_AGEMA_signal_3721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C ( clk ), .D ( n2483 ), .Q ( new_AGEMA_signal_3725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C ( clk ), .D ( new_AGEMA_signal_1107 ), .Q ( new_AGEMA_signal_3729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C ( clk ), .D ( n2629 ), .Q ( new_AGEMA_signal_3769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C ( clk ), .D ( new_AGEMA_signal_1120 ), .Q ( new_AGEMA_signal_3773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C ( clk ), .D ( n2736 ), .Q ( new_AGEMA_signal_3797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C ( clk ), .D ( new_AGEMA_signal_1051 ), .Q ( new_AGEMA_signal_3801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C ( clk ), .D ( new_AGEMA_signal_2950 ), .Q ( new_AGEMA_signal_3805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C ( clk ), .D ( new_AGEMA_signal_2952 ), .Q ( new_AGEMA_signal_3809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C ( clk ), .D ( new_AGEMA_signal_2894 ), .Q ( new_AGEMA_signal_3813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C ( clk ), .D ( new_AGEMA_signal_2896 ), .Q ( new_AGEMA_signal_3817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C ( clk ), .D ( n2787 ), .Q ( new_AGEMA_signal_3821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C ( clk ), .D ( new_AGEMA_signal_1303 ), .Q ( new_AGEMA_signal_3825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C ( clk ), .D ( new_AGEMA_signal_3846 ), .Q ( new_AGEMA_signal_3847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C ( clk ), .D ( new_AGEMA_signal_3854 ), .Q ( new_AGEMA_signal_3855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C ( clk ), .D ( new_AGEMA_signal_3866 ), .Q ( new_AGEMA_signal_3867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C ( clk ), .D ( new_AGEMA_signal_3874 ), .Q ( new_AGEMA_signal_3875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C ( clk ), .D ( n2009 ), .Q ( new_AGEMA_signal_3881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C ( clk ), .D ( new_AGEMA_signal_1162 ), .Q ( new_AGEMA_signal_3887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C ( clk ), .D ( n2034 ), .Q ( new_AGEMA_signal_3901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_3907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C ( clk ), .D ( new_AGEMA_signal_3034 ), .Q ( new_AGEMA_signal_3917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C ( clk ), .D ( new_AGEMA_signal_3036 ), .Q ( new_AGEMA_signal_3923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C ( clk ), .D ( new_AGEMA_signal_3062 ), .Q ( new_AGEMA_signal_3929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C ( clk ), .D ( new_AGEMA_signal_3064 ), .Q ( new_AGEMA_signal_3935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C ( clk ), .D ( new_AGEMA_signal_2810 ), .Q ( new_AGEMA_signal_3953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C ( clk ), .D ( new_AGEMA_signal_2812 ), .Q ( new_AGEMA_signal_3959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C ( clk ), .D ( n2122 ), .Q ( new_AGEMA_signal_3965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C ( clk ), .D ( new_AGEMA_signal_1193 ), .Q ( new_AGEMA_signal_3971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C ( clk ), .D ( n2220 ), .Q ( new_AGEMA_signal_3981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C ( clk ), .D ( new_AGEMA_signal_1199 ), .Q ( new_AGEMA_signal_3987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C ( clk ), .D ( new_AGEMA_signal_4018 ), .Q ( new_AGEMA_signal_4019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C ( clk ), .D ( new_AGEMA_signal_4026 ), .Q ( new_AGEMA_signal_4027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C ( clk ), .D ( new_AGEMA_signal_2910 ), .Q ( new_AGEMA_signal_4033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C ( clk ), .D ( new_AGEMA_signal_2912 ), .Q ( new_AGEMA_signal_4039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C ( clk ), .D ( n2344 ), .Q ( new_AGEMA_signal_4089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C ( clk ), .D ( new_AGEMA_signal_1239 ), .Q ( new_AGEMA_signal_4095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C ( clk ), .D ( n2468 ), .Q ( new_AGEMA_signal_4153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C ( clk ), .D ( new_AGEMA_signal_1110 ), .Q ( new_AGEMA_signal_4159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C ( clk ), .D ( n2761 ), .Q ( new_AGEMA_signal_4165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C ( clk ), .D ( new_AGEMA_signal_1144 ), .Q ( new_AGEMA_signal_4171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C ( clk ), .D ( new_AGEMA_signal_4190 ), .Q ( new_AGEMA_signal_4191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C ( clk ), .D ( new_AGEMA_signal_4198 ), .Q ( new_AGEMA_signal_4199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C ( clk ), .D ( new_AGEMA_signal_4250 ), .Q ( new_AGEMA_signal_4251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C ( clk ), .D ( new_AGEMA_signal_4258 ), .Q ( new_AGEMA_signal_4259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C ( clk ), .D ( n2825 ), .Q ( new_AGEMA_signal_4281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C ( clk ), .D ( new_AGEMA_signal_1308 ), .Q ( new_AGEMA_signal_4287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C ( clk ), .D ( n1957 ), .Q ( new_AGEMA_signal_4297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C ( clk ), .D ( new_AGEMA_signal_1049 ), .Q ( new_AGEMA_signal_4305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C ( clk ), .D ( n2026 ), .Q ( new_AGEMA_signal_4325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_4333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C ( clk ), .D ( n2811 ), .Q ( new_AGEMA_signal_4365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C ( clk ), .D ( new_AGEMA_signal_1194 ), .Q ( new_AGEMA_signal_4373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C ( clk ), .D ( new_AGEMA_signal_3074 ), .Q ( new_AGEMA_signal_4457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C ( clk ), .D ( new_AGEMA_signal_3076 ), .Q ( new_AGEMA_signal_4465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C ( clk ), .D ( n2363 ), .Q ( new_AGEMA_signal_4493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_4501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C ( clk ), .D ( new_AGEMA_signal_3030 ), .Q ( new_AGEMA_signal_4557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C ( clk ), .D ( new_AGEMA_signal_3032 ), .Q ( new_AGEMA_signal_4565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C ( clk ), .D ( new_AGEMA_signal_2830 ), .Q ( new_AGEMA_signal_4573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C ( clk ), .D ( new_AGEMA_signal_2832 ), .Q ( new_AGEMA_signal_4581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C ( clk ), .D ( n2544 ), .Q ( new_AGEMA_signal_4745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C ( clk ), .D ( new_AGEMA_signal_1079 ), .Q ( new_AGEMA_signal_4755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C ( clk ), .D ( n2364 ), .Q ( new_AGEMA_signal_4845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C ( clk ), .D ( new_AGEMA_signal_1245 ), .Q ( new_AGEMA_signal_4855 ) ) ;

    /* cells in depth 6 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1960 ( .a ({new_AGEMA_signal_1127, n2575}), .b ({new_AGEMA_signal_1128, n1962}), .clk ( clk ), .r ( Fresh[238] ), .c ({new_AGEMA_signal_1309, n1924}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1967 ( .a ({new_AGEMA_signal_1129, n1922}), .b ({new_AGEMA_signal_2808, new_AGEMA_signal_2806}), .clk ( clk ), .r ( Fresh[239] ), .c ({new_AGEMA_signal_1310, n1923}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1981 ( .a ({new_AGEMA_signal_1130, n1926}), .b ({new_AGEMA_signal_1131, n1925}), .clk ( clk ), .r ( Fresh[240] ), .c ({new_AGEMA_signal_1311, n1927}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1993 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_1134, n2763}), .clk ( clk ), .r ( Fresh[241] ), .c ({new_AGEMA_signal_1312, n1929}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2007 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[242] ), .c ({new_AGEMA_signal_1313, n2665}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2011 ( .a ({new_AGEMA_signal_2816, new_AGEMA_signal_2814}), .b ({new_AGEMA_signal_1136, n1937}), .clk ( clk ), .r ( Fresh[243] ), .c ({new_AGEMA_signal_1314, n1938}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2019 ( .a ({new_AGEMA_signal_2820, new_AGEMA_signal_2818}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[244] ), .c ({new_AGEMA_signal_1315, n2235}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2023 ( .a ({new_AGEMA_signal_2824, new_AGEMA_signal_2822}), .b ({new_AGEMA_signal_1042, n1942}), .clk ( clk ), .r ( Fresh[245] ), .c ({new_AGEMA_signal_1137, n1943}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2027 ( .a ({new_AGEMA_signal_1043, n2676}), .b ({new_AGEMA_signal_2828, new_AGEMA_signal_2826}), .clk ( clk ), .r ( Fresh[246] ), .c ({new_AGEMA_signal_1138, n1946}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2031 ( .a ({new_AGEMA_signal_2832, new_AGEMA_signal_2830}), .b ({new_AGEMA_signal_1139, n1944}), .clk ( clk ), .r ( Fresh[247] ), .c ({new_AGEMA_signal_1316, n1945}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2034 ( .a ({new_AGEMA_signal_2836, new_AGEMA_signal_2834}), .b ({new_AGEMA_signal_1133, n2734}), .clk ( clk ), .r ( Fresh[248] ), .c ({new_AGEMA_signal_1317, n1956}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2040 ( .a ({new_AGEMA_signal_1140, n1950}), .b ({new_AGEMA_signal_1046, n1949}), .clk ( clk ), .r ( Fresh[249] ), .c ({new_AGEMA_signal_1318, n1951}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2048 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ( Fresh[250] ), .c ({new_AGEMA_signal_1319, n1952}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2057 ( .a ({new_AGEMA_signal_2840, new_AGEMA_signal_2838}), .b ({new_AGEMA_signal_1142, n2088}), .clk ( clk ), .r ( Fresh[251] ), .c ({new_AGEMA_signal_1320, n2687}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) U2061 ( .a ({new_AGEMA_signal_1128, n1962}), .b ({new_AGEMA_signal_2844, new_AGEMA_signal_2842}), .clk ( clk ), .r ( Fresh[252] ), .c ({new_AGEMA_signal_1321, n1966}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2064 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_2848, new_AGEMA_signal_2846}), .clk ( clk ), .r ( Fresh[253] ), .c ({new_AGEMA_signal_1143, n1963}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2077 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ( Fresh[254] ), .c ({new_AGEMA_signal_1480, n1968}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2082 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[255] ), .c ({new_AGEMA_signal_1325, n2684}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2088 ( .a ({new_AGEMA_signal_2852, new_AGEMA_signal_2850}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ( Fresh[256] ), .c ({new_AGEMA_signal_1326, n1972}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2092 ( .a ({new_AGEMA_signal_2856, new_AGEMA_signal_2854}), .b ({new_AGEMA_signal_1059, n2190}), .clk ( clk ), .r ( Fresh[257] ), .c ({new_AGEMA_signal_1149, n1971}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2099 ( .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2858}), .b ({new_AGEMA_signal_1150, n2535}), .clk ( clk ), .r ( Fresh[258] ), .c ({new_AGEMA_signal_1327, n1974}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2106 ( .a ({new_AGEMA_signal_1135, n2732}), .b ({new_AGEMA_signal_2840, new_AGEMA_signal_2838}), .clk ( clk ), .r ( Fresh[259] ), .c ({new_AGEMA_signal_1328, n1979}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2112 ( .a ({new_AGEMA_signal_2864, new_AGEMA_signal_2862}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[260] ), .c ({new_AGEMA_signal_1152, n1985}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2121 ( .a ({new_AGEMA_signal_1154, n1992}), .b ({new_AGEMA_signal_1155, n1991}), .clk ( clk ), .r ( Fresh[261] ), .c ({new_AGEMA_signal_1330, n1994}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2126 ( .a ({new_AGEMA_signal_2868, new_AGEMA_signal_2866}), .b ({new_AGEMA_signal_1156, n1995}), .clk ( clk ), .r ( Fresh[262] ), .c ({new_AGEMA_signal_1331, n1996}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2136 ( .a ({new_AGEMA_signal_2872, new_AGEMA_signal_2870}), .b ({new_AGEMA_signal_1158, n2003}), .clk ( clk ), .r ( Fresh[263] ), .c ({new_AGEMA_signal_1332, n2137}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2142 ( .a ({new_AGEMA_signal_2876, new_AGEMA_signal_2874}), .b ({new_AGEMA_signal_1160, n2572}), .clk ( clk ), .r ( Fresh[264] ), .c ({new_AGEMA_signal_1333, n2006}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2144 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2878}), .b ({new_AGEMA_signal_1161, n2004}), .clk ( clk ), .r ( Fresh[265] ), .c ({new_AGEMA_signal_1334, n2005}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2152 ( .a ({new_AGEMA_signal_2884, new_AGEMA_signal_2882}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[266] ), .c ({new_AGEMA_signal_1335, n2013}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2160 ( .a ({new_AGEMA_signal_2888, new_AGEMA_signal_2886}), .b ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .r ( Fresh[267] ), .c ({new_AGEMA_signal_1165, n2020}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2164 ( .a ({new_AGEMA_signal_1062, n2817}), .b ({new_AGEMA_signal_2892, new_AGEMA_signal_2890}), .clk ( clk ), .r ( Fresh[268] ), .c ({new_AGEMA_signal_1166, n2023}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2168 ( .a ({new_AGEMA_signal_1009, n2027}), .b ({new_AGEMA_signal_2896, new_AGEMA_signal_2894}), .clk ( clk ), .r ( Fresh[269] ), .c ({new_AGEMA_signal_1071, n2028}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2172 ( .a ({new_AGEMA_signal_1167, n2214}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[270] ), .c ({new_AGEMA_signal_1337, n2033}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2175 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_2904, new_AGEMA_signal_2902}), .clk ( clk ), .r ( Fresh[271] ), .c ({new_AGEMA_signal_1338, n2031}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2184 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1170, n2039}), .clk ( clk ), .r ( Fresh[272] ), .c ({new_AGEMA_signal_1339, n2040}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2187 ( .a ({new_AGEMA_signal_2908, new_AGEMA_signal_2906}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[273] ), .c ({new_AGEMA_signal_1171, n2050}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2193 ( .a ({new_AGEMA_signal_2912, new_AGEMA_signal_2910}), .b ({new_AGEMA_signal_1174, n2044}), .clk ( clk ), .r ( Fresh[274] ), .c ({new_AGEMA_signal_1340, n2045}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2199 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_2840, new_AGEMA_signal_2838}), .clk ( clk ), .r ( Fresh[275] ), .c ({new_AGEMA_signal_1341, n2051}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2203 ( .a ({new_AGEMA_signal_2916, new_AGEMA_signal_2914}), .b ({new_AGEMA_signal_1176, n2055}), .clk ( clk ), .r ( Fresh[276] ), .c ({new_AGEMA_signal_1342, n2056}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2209 ( .a ({new_AGEMA_signal_1178, n2407}), .b ({new_AGEMA_signal_2920, new_AGEMA_signal_2918}), .clk ( clk ), .r ( Fresh[277] ), .c ({new_AGEMA_signal_1343, n2060}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2215 ( .a ({new_AGEMA_signal_2924, new_AGEMA_signal_2922}), .b ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .r ( Fresh[278] ), .c ({new_AGEMA_signal_1344, n2066}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2217 ( .a ({new_AGEMA_signal_2896, new_AGEMA_signal_2894}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ( Fresh[279] ), .c ({new_AGEMA_signal_1345, n2065}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2221 ( .a ({new_AGEMA_signal_1181, n2068}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[280] ), .c ({new_AGEMA_signal_1346, n2069}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2226 ( .a ({new_AGEMA_signal_2928, new_AGEMA_signal_2926}), .b ({new_AGEMA_signal_1182, n2252}), .clk ( clk ), .r ( Fresh[281] ), .c ({new_AGEMA_signal_1347, n2074}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2235 ( .a ({new_AGEMA_signal_1076, n2081}), .b ({new_AGEMA_signal_1183, n2080}), .clk ( clk ), .r ( Fresh[282] ), .c ({new_AGEMA_signal_1348, n2082}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2240 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2878}), .b ({new_AGEMA_signal_1185, n2083}), .clk ( clk ), .r ( Fresh[283] ), .c ({new_AGEMA_signal_1349, n2084}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2242 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .clk ( clk ), .r ( Fresh[284] ), .c ({new_AGEMA_signal_1350, n2085}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2245 ( .a ({new_AGEMA_signal_2932, new_AGEMA_signal_2930}), .b ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .r ( Fresh[285] ), .c ({new_AGEMA_signal_1351, n2131}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2248 ( .a ({new_AGEMA_signal_1142, n2088}), .b ({new_AGEMA_signal_1078, n2087}), .clk ( clk ), .r ( Fresh[286] ), .c ({new_AGEMA_signal_1352, n2089}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2252 ( .a ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .b ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .r ( Fresh[287] ), .c ({new_AGEMA_signal_1353, n2330}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2254 ( .a ({new_AGEMA_signal_2936, new_AGEMA_signal_2934}), .b ({new_AGEMA_signal_1132, n2151}), .clk ( clk ), .r ( Fresh[288] ), .c ({new_AGEMA_signal_1354, n2092}) ) ;
    or_HPC2 #(.security_order(1), .pipeline(1)) U2256 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1147, n2359}), .clk ( clk ), .r ( Fresh[289] ), .c ({new_AGEMA_signal_1355, n2094}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2261 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1188, n2100}), .clk ( clk ), .r ( Fresh[290] ), .c ({new_AGEMA_signal_1356, n2160}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2265 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[291] ), .c ({new_AGEMA_signal_1189, n2504}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2271 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[292] ), .c ({new_AGEMA_signal_1504, n2114}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2273 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_2880, new_AGEMA_signal_2878}), .clk ( clk ), .r ( Fresh[293] ), .c ({new_AGEMA_signal_1190, n2115}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2280 ( .a ({new_AGEMA_signal_2940, new_AGEMA_signal_2938}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ( Fresh[294] ), .c ({new_AGEMA_signal_1358, n2291}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2281 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[295] ), .c ({new_AGEMA_signal_1192, n2119}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2291 ( .a ({new_AGEMA_signal_2944, new_AGEMA_signal_2942}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[296] ), .c ({new_AGEMA_signal_1195, n2130}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2292 ( .a ({new_AGEMA_signal_1062, n2817}), .b ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .r ( Fresh[297] ), .c ({new_AGEMA_signal_1196, n2129}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2295 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .clk ( clk ), .r ( Fresh[298] ), .c ({new_AGEMA_signal_1197, n2150}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2298 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1082, n2132}), .clk ( clk ), .r ( Fresh[299] ), .c ({new_AGEMA_signal_1198, n2133}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2302 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_2952, new_AGEMA_signal_2950}), .clk ( clk ), .r ( Fresh[300] ), .c ({new_AGEMA_signal_1361, n2136}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2306 ( .a ({new_AGEMA_signal_1160, n2572}), .b ({new_AGEMA_signal_1200, n2138}), .clk ( clk ), .r ( Fresh[301] ), .c ({new_AGEMA_signal_1362, n2139}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2313 ( .a ({new_AGEMA_signal_2956, new_AGEMA_signal_2954}), .b ({new_AGEMA_signal_1201, n2555}), .clk ( clk ), .r ( Fresh[302] ), .c ({new_AGEMA_signal_1363, n2144}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2318 ( .a ({new_AGEMA_signal_1132, n2151}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[303] ), .c ({new_AGEMA_signal_1364, n2152}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2321 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .r ( Fresh[304] ), .c ({new_AGEMA_signal_1365, n2170}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2323 ( .a ({new_AGEMA_signal_1202, n2429}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[305] ), .c ({new_AGEMA_signal_1366, n2157}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2329 ( .a ({new_AGEMA_signal_2960, new_AGEMA_signal_2958}), .b ({new_AGEMA_signal_1083, n2162}), .clk ( clk ), .r ( Fresh[306] ), .c ({new_AGEMA_signal_1203, n2163}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2335 ( .a ({new_AGEMA_signal_1073, n2171}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ( Fresh[307] ), .c ({new_AGEMA_signal_1368, n2172}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2338 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .b ({new_AGEMA_signal_1014, n2545}), .clk ( clk ), .r ( Fresh[308] ), .c ({new_AGEMA_signal_1084, n2186}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2339 ( .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2858}), .b ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .r ( Fresh[309] ), .c ({new_AGEMA_signal_1369, n2181}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2344 ( .a ({new_AGEMA_signal_1204, n2176}), .b ({new_AGEMA_signal_1205, n2175}), .clk ( clk ), .r ( Fresh[310] ), .c ({new_AGEMA_signal_1370, n2177}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2349 ( .a ({new_AGEMA_signal_2840, new_AGEMA_signal_2838}), .b ({new_AGEMA_signal_1016, n2182}), .clk ( clk ), .r ( Fresh[311] ), .c ({new_AGEMA_signal_1086, n2183}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2354 ( .a ({new_AGEMA_signal_2964, new_AGEMA_signal_2962}), .b ({new_AGEMA_signal_1206, n2188}), .clk ( clk ), .r ( Fresh[312] ), .c ({new_AGEMA_signal_1371, n2195}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2356 ( .a ({new_AGEMA_signal_1059, n2190}), .b ({new_AGEMA_signal_1207, n2189}), .clk ( clk ), .r ( Fresh[313] ), .c ({new_AGEMA_signal_1372, n2193}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2358 ( .a ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .b ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .r ( Fresh[314] ), .c ({new_AGEMA_signal_1373, n2191}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2364 ( .a ({new_AGEMA_signal_1087, n2576}), .b ({new_AGEMA_signal_1088, n2748}), .clk ( clk ), .r ( Fresh[315] ), .c ({new_AGEMA_signal_1209, n2196}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2367 ( .a ({new_AGEMA_signal_2828, new_AGEMA_signal_2826}), .b ({new_AGEMA_signal_1146, n2505}), .clk ( clk ), .r ( Fresh[316] ), .c ({new_AGEMA_signal_1374, n2201}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2369 ( .a ({new_AGEMA_signal_1375, n2674}), .b ({new_AGEMA_signal_2972, new_AGEMA_signal_2970}), .clk ( clk ), .r ( Fresh[317] ), .c ({new_AGEMA_signal_1515, n2200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2371 ( .s ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .b ({new_AGEMA_signal_1133, n2734}), .a ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ( Fresh[318] ), .c ({new_AGEMA_signal_1516, n2202}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2379 ( .a ({new_AGEMA_signal_1167, n2214}), .b ({new_AGEMA_signal_1089, n2213}), .clk ( clk ), .r ( Fresh[319] ), .c ({new_AGEMA_signal_1376, n2217}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2381 ( .a ({new_AGEMA_signal_2976, new_AGEMA_signal_2974}), .b ({new_AGEMA_signal_1090, n2215}), .clk ( clk ), .r ( Fresh[320] ), .c ({new_AGEMA_signal_1210, n2216}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2385 ( .a ({new_AGEMA_signal_1211, n2218}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .clk ( clk ), .r ( Fresh[321] ), .c ({new_AGEMA_signal_1377, n2222}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2387 ( .a ({new_AGEMA_signal_1199, n2220}), .b ({new_AGEMA_signal_1212, n2219}), .clk ( clk ), .r ( Fresh[322] ), .c ({new_AGEMA_signal_1378, n2221}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2391 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_2980, new_AGEMA_signal_2978}), .clk ( clk ), .r ( Fresh[323] ), .c ({new_AGEMA_signal_1213, n2226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2393 ( .s ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .b ({new_AGEMA_signal_1056, n2651}), .a ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .r ( Fresh[324] ), .c ({new_AGEMA_signal_1214, n2228}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2397 ( .a ({new_AGEMA_signal_2888, new_AGEMA_signal_2886}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[325] ), .c ({new_AGEMA_signal_1215, n2237}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2398 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .clk ( clk ), .r ( Fresh[326] ), .c ({new_AGEMA_signal_1520, n2233}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2403 ( .a ({new_AGEMA_signal_2984, new_AGEMA_signal_2982}), .b ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .r ( Fresh[327] ), .c ({new_AGEMA_signal_1216, n2238}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2406 ( .a ({new_AGEMA_signal_1157, n2241}), .b ({new_AGEMA_signal_1217, n2240}), .clk ( clk ), .r ( Fresh[328] ), .c ({new_AGEMA_signal_1380, n2248}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2409 ( .a ({new_AGEMA_signal_1218, n2561}), .b ({new_AGEMA_signal_1219, n2243}), .clk ( clk ), .r ( Fresh[329] ), .c ({new_AGEMA_signal_1381, n2244}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2414 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_2808, new_AGEMA_signal_2806}), .clk ( clk ), .r ( Fresh[330] ), .c ({new_AGEMA_signal_1382, n2249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2417 ( .s ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .b ({new_AGEMA_signal_1182, n2252}), .a ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[331] ), .c ({new_AGEMA_signal_1383, n2253}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2424 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_1222, n2259}), .clk ( clk ), .r ( Fresh[332] ), .c ({new_AGEMA_signal_1384, n2260}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2429 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_2988, new_AGEMA_signal_2986}), .clk ( clk ), .r ( Fresh[333] ), .c ({new_AGEMA_signal_1524, n2273}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2430 ( .a ({new_AGEMA_signal_2992, new_AGEMA_signal_2990}), .b ({new_AGEMA_signal_1323, n2720}), .clk ( clk ), .r ( Fresh[334] ), .c ({new_AGEMA_signal_1525, n2752}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2433 ( .a ({new_AGEMA_signal_1093, n2645}), .b ({new_AGEMA_signal_2940, new_AGEMA_signal_2938}), .clk ( clk ), .r ( Fresh[335] ), .c ({new_AGEMA_signal_1223, n2265}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2437 ( .a ({new_AGEMA_signal_2996, new_AGEMA_signal_2994}), .b ({new_AGEMA_signal_1094, n2268}), .clk ( clk ), .r ( Fresh[336] ), .c ({new_AGEMA_signal_1224, n2269}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2444 ( .a ({new_AGEMA_signal_2848, new_AGEMA_signal_2846}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[337] ), .c ({new_AGEMA_signal_1226, n2277}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2449 ( .a ({new_AGEMA_signal_3000, new_AGEMA_signal_2998}), .b ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .r ( Fresh[338] ), .c ({new_AGEMA_signal_1227, n2282}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2452 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[339] ), .c ({new_AGEMA_signal_1389, n2284}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2456 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_3004, new_AGEMA_signal_3002}), .clk ( clk ), .r ( Fresh[340] ), .c ({new_AGEMA_signal_1390, n2459}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2459 ( .a ({new_AGEMA_signal_2816, new_AGEMA_signal_2814}), .b ({new_AGEMA_signal_1229, n2287}), .clk ( clk ), .r ( Fresh[341] ), .c ({new_AGEMA_signal_1391, n2288}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2462 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .b ({new_AGEMA_signal_1144, n2761}), .clk ( clk ), .r ( Fresh[342] ), .c ({new_AGEMA_signal_1392, n2458}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2464 ( .a ({new_AGEMA_signal_2960, new_AGEMA_signal_2958}), .b ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .r ( Fresh[343] ), .c ({new_AGEMA_signal_1393, n2293}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2467 ( .a ({new_AGEMA_signal_2936, new_AGEMA_signal_2934}), .b ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .r ( Fresh[344] ), .c ({new_AGEMA_signal_1230, n2294}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2472 ( .a ({new_AGEMA_signal_1231, n2438}), .b ({new_AGEMA_signal_1096, n2299}), .clk ( clk ), .r ( Fresh[345] ), .c ({new_AGEMA_signal_1394, n2300}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2480 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .clk ( clk ), .r ( Fresh[346] ), .c ({new_AGEMA_signal_1395, n2323}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) U2482 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1232, n2371}), .clk ( clk ), .r ( Fresh[347] ), .c ({new_AGEMA_signal_1396, n2314}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2485 ( .a ({new_AGEMA_signal_1018, n2316}), .b ({new_AGEMA_signal_3008, new_AGEMA_signal_3006}), .clk ( clk ), .r ( Fresh[348] ), .c ({new_AGEMA_signal_1097, n2319}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2491 ( .a ({new_AGEMA_signal_1074, n2642}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[349] ), .c ({new_AGEMA_signal_1234, n2326}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2496 ( .a ({new_AGEMA_signal_1236, n2328}), .b ({new_AGEMA_signal_1099, n2327}), .clk ( clk ), .r ( Fresh[350] ), .c ({new_AGEMA_signal_1398, n2329}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2501 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[351] ), .c ({new_AGEMA_signal_1537, n2335}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2506 ( .a ({new_AGEMA_signal_2884, new_AGEMA_signal_2882}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ( Fresh[352] ), .c ({new_AGEMA_signal_1399, n2341}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2507 ( .a ({new_AGEMA_signal_3012, new_AGEMA_signal_3010}), .b ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .r ( Fresh[353] ), .c ({new_AGEMA_signal_1238, n2340}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2514 ( .a ({new_AGEMA_signal_1100, n2348}), .b ({new_AGEMA_signal_1101, n2347}), .clk ( clk ), .r ( Fresh[354] ), .c ({new_AGEMA_signal_1240, n2349}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2517 ( .a ({new_AGEMA_signal_3016, new_AGEMA_signal_3014}), .b ({new_AGEMA_signal_1061, n2690}), .clk ( clk ), .r ( Fresh[355] ), .c ({new_AGEMA_signal_1241, n2375}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2518 ( .a ({new_AGEMA_signal_2956, new_AGEMA_signal_2954}), .b ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .r ( Fresh[356] ), .c ({new_AGEMA_signal_1242, n2352}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2522 ( .a ({new_AGEMA_signal_1243, n2353}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[357] ), .c ({new_AGEMA_signal_1401, n2354}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2525 ( .a ({new_AGEMA_signal_3020, new_AGEMA_signal_3018}), .b ({new_AGEMA_signal_1244, n2355}), .clk ( clk ), .r ( Fresh[358] ), .c ({new_AGEMA_signal_1402, n2357}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2527 ( .a ({new_AGEMA_signal_1147, n2359}), .b ({new_AGEMA_signal_3024, new_AGEMA_signal_3022}), .clk ( clk ), .r ( Fresh[359] ), .c ({new_AGEMA_signal_1403, n2360}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2534 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[360] ), .c ({new_AGEMA_signal_1540, n2369}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2536 ( .a ({new_AGEMA_signal_1232, n2371}), .b ({new_AGEMA_signal_2980, new_AGEMA_signal_2978}), .clk ( clk ), .r ( Fresh[361] ), .c ({new_AGEMA_signal_1404, n2372}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2539 ( .a ({new_AGEMA_signal_1087, n2576}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ( Fresh[362] ), .c ({new_AGEMA_signal_1405, n2377}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2544 ( .a ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .b ({new_AGEMA_signal_1103, n2415}), .clk ( clk ), .r ( Fresh[363] ), .c ({new_AGEMA_signal_1246, n2467}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2545 ( .a ({new_AGEMA_signal_3028, new_AGEMA_signal_3026}), .b ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .r ( Fresh[364] ), .c ({new_AGEMA_signal_1247, n2385}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2546 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[365] ), .c ({new_AGEMA_signal_1248, n2384}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2548 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2878}), .b ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .r ( Fresh[366] ), .c ({new_AGEMA_signal_1407, n2386}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2552 ( .a ({new_AGEMA_signal_2964, new_AGEMA_signal_2962}), .b ({new_AGEMA_signal_1081, n2647}), .clk ( clk ), .r ( Fresh[367] ), .c ({new_AGEMA_signal_1249, n2394}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2553 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .clk ( clk ), .r ( Fresh[368] ), .c ({new_AGEMA_signal_1250, n2391}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2554 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[369] ), .c ({new_AGEMA_signal_1408, n2390}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2559 ( .a ({new_AGEMA_signal_2936, new_AGEMA_signal_2934}), .b ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .r ( Fresh[370] ), .c ({new_AGEMA_signal_1251, n2396}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2562 ( .a ({new_AGEMA_signal_3032, new_AGEMA_signal_3030}), .b ({new_AGEMA_signal_1231, n2438}), .clk ( clk ), .r ( Fresh[371] ), .c ({new_AGEMA_signal_1409, n2406}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2565 ( .a ({new_AGEMA_signal_1105, n2594}), .b ({new_AGEMA_signal_1106, n2402}), .clk ( clk ), .r ( Fresh[372] ), .c ({new_AGEMA_signal_1252, n2403}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2569 ( .a ({new_AGEMA_signal_1178, n2407}), .b ({new_AGEMA_signal_2952, new_AGEMA_signal_2950}), .clk ( clk ), .r ( Fresh[373] ), .c ({new_AGEMA_signal_1411, n2408}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2573 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_2984, new_AGEMA_signal_2982}), .clk ( clk ), .r ( Fresh[374] ), .c ({new_AGEMA_signal_1412, n2574}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2574 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_2912, new_AGEMA_signal_2910}), .clk ( clk ), .r ( Fresh[375] ), .c ({new_AGEMA_signal_1253, n2413}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2577 ( .a ({new_AGEMA_signal_1103, n2415}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[376] ), .c ({new_AGEMA_signal_1254, n2416}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2586 ( .a ({new_AGEMA_signal_1255, n2428}), .b ({new_AGEMA_signal_3036, new_AGEMA_signal_3034}), .clk ( clk ), .r ( Fresh[377] ), .c ({new_AGEMA_signal_1414, n2433}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2587 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .b ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .r ( Fresh[378] ), .c ({new_AGEMA_signal_1415, n2689}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2591 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .r ( Fresh[379] ), .c ({new_AGEMA_signal_1257, n2434}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2595 ( .a ({new_AGEMA_signal_1231, n2438}), .b ({new_AGEMA_signal_1107, n2483}), .clk ( clk ), .r ( Fresh[380] ), .c ({new_AGEMA_signal_1417, n2439}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2598 ( .a ({new_AGEMA_signal_3028, new_AGEMA_signal_3026}), .b ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .r ( Fresh[381] ), .c ({new_AGEMA_signal_1418, n2445}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2600 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1258, n2443}), .clk ( clk ), .r ( Fresh[382] ), .c ({new_AGEMA_signal_1419, n2444}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2602 ( .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2858}), .b ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .r ( Fresh[383] ), .c ({new_AGEMA_signal_1420, n2447}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2607 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .r ( Fresh[384] ), .c ({new_AGEMA_signal_1421, n2454}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2617 ( .a ({new_AGEMA_signal_2940, new_AGEMA_signal_2938}), .b ({new_AGEMA_signal_1109, n2464}), .clk ( clk ), .r ( Fresh[385] ), .c ({new_AGEMA_signal_1260, n2465}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2622 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .b ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .r ( Fresh[386] ), .c ({new_AGEMA_signal_1261, n2470}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2626 ( .a ({new_AGEMA_signal_1111, n2473}), .b ({new_AGEMA_signal_1112, n2472}), .clk ( clk ), .r ( Fresh[387] ), .c ({new_AGEMA_signal_1262, n2476}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2633 ( .a ({new_AGEMA_signal_3040, new_AGEMA_signal_3038}), .b ({new_AGEMA_signal_1263, n2480}), .clk ( clk ), .r ( Fresh[388] ), .c ({new_AGEMA_signal_1424, n2481}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2639 ( .a ({new_AGEMA_signal_3044, new_AGEMA_signal_3042}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[389] ), .c ({new_AGEMA_signal_1265, n2486}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2642 ( .a ({new_AGEMA_signal_2992, new_AGEMA_signal_2990}), .b ({new_AGEMA_signal_1114, n2488}), .clk ( clk ), .r ( Fresh[390] ), .c ({new_AGEMA_signal_1266, n2489}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2645 ( .a ({new_AGEMA_signal_3048, new_AGEMA_signal_3046}), .b ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .r ( Fresh[391] ), .c ({new_AGEMA_signal_1267, n2497}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2646 ( .a ({new_AGEMA_signal_3052, new_AGEMA_signal_3050}), .b ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .r ( Fresh[392] ), .c ({new_AGEMA_signal_1268, n2495}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2647 ( .a ({new_AGEMA_signal_2944, new_AGEMA_signal_2942}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ( Fresh[393] ), .c ({new_AGEMA_signal_1426, n2494}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2650 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_2828, new_AGEMA_signal_2826}), .clk ( clk ), .r ( Fresh[394] ), .c ({new_AGEMA_signal_1269, n2499}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2653 ( .a ({new_AGEMA_signal_2828, new_AGEMA_signal_2826}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[395] ), .c ({new_AGEMA_signal_1557, n2503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2655 ( .s ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .b ({new_AGEMA_signal_1146, n2505}), .a ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[396] ), .c ({new_AGEMA_signal_1427, n2506}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2662 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_2872, new_AGEMA_signal_2870}), .clk ( clk ), .r ( Fresh[397] ), .c ({new_AGEMA_signal_1428, n2518}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2663 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[398] ), .c ({new_AGEMA_signal_1558, n2517}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2666 ( .a ({new_AGEMA_signal_1270, n2520}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .clk ( clk ), .r ( Fresh[399] ), .c ({new_AGEMA_signal_1429, n2523}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2668 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_1115, n2521}), .clk ( clk ), .r ( Fresh[400] ), .c ({new_AGEMA_signal_1430, n2522}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2675 ( .a ({new_AGEMA_signal_2872, new_AGEMA_signal_2870}), .b ({new_AGEMA_signal_1271, n2531}), .clk ( clk ), .r ( Fresh[401] ), .c ({new_AGEMA_signal_1431, n2532}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2677 ( .a ({new_AGEMA_signal_2808, new_AGEMA_signal_2806}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[402] ), .c ({new_AGEMA_signal_1432, n2534}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2681 ( .a ({new_AGEMA_signal_3056, new_AGEMA_signal_3054}), .b ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .r ( Fresh[403] ), .c ({new_AGEMA_signal_1433, n2542}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2683 ( .a ({new_AGEMA_signal_1014, n2545}), .b ({new_AGEMA_signal_1079, n2544}), .clk ( clk ), .r ( Fresh[404] ), .c ({new_AGEMA_signal_1272, n2546}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2687 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[405] ), .c ({new_AGEMA_signal_1435, n2551}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2690 ( .a ({new_AGEMA_signal_1273, n2553}), .b ({new_AGEMA_signal_3060, new_AGEMA_signal_3058}), .clk ( clk ), .r ( Fresh[406] ), .c ({new_AGEMA_signal_1436, n2558}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2692 ( .a ({new_AGEMA_signal_1201, n2555}), .b ({new_AGEMA_signal_1274, n2554}), .clk ( clk ), .r ( Fresh[407] ), .c ({new_AGEMA_signal_1437, n2556}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2696 ( .a ({new_AGEMA_signal_1218, n2561}), .b ({new_AGEMA_signal_1116, n2560}), .clk ( clk ), .r ( Fresh[408] ), .c ({new_AGEMA_signal_1438, n2566}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2697 ( .a ({new_AGEMA_signal_3064, new_AGEMA_signal_3062}), .b ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .r ( Fresh[409] ), .c ({new_AGEMA_signal_1439, n2715}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2703 ( .a ({new_AGEMA_signal_1160, n2572}), .b ({new_AGEMA_signal_1055, n2571}), .clk ( clk ), .r ( Fresh[410] ), .c ({new_AGEMA_signal_1440, n2573}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2705 ( .a ({new_AGEMA_signal_3032, new_AGEMA_signal_3030}), .b ({new_AGEMA_signal_1173, n2754}), .clk ( clk ), .r ( Fresh[411] ), .c ({new_AGEMA_signal_1441, n2585}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2706 ( .a ({new_AGEMA_signal_2988, new_AGEMA_signal_2986}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ( Fresh[412] ), .c ({new_AGEMA_signal_1276, n2581}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2707 ( .a ({new_AGEMA_signal_1127, n2575}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[413] ), .c ({new_AGEMA_signal_1442, n2579}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2708 ( .a ({new_AGEMA_signal_3052, new_AGEMA_signal_3050}), .b ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .r ( Fresh[414] ), .c ({new_AGEMA_signal_1277, n2578}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2711 ( .a ({new_AGEMA_signal_1148, n2625}), .b ({new_AGEMA_signal_2972, new_AGEMA_signal_2970}), .clk ( clk ), .r ( Fresh[415] ), .c ({new_AGEMA_signal_1443, n2582}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2715 ( .a ({new_AGEMA_signal_2844, new_AGEMA_signal_2842}), .b ({new_AGEMA_signal_1278, n2586}), .clk ( clk ), .r ( Fresh[416] ), .c ({new_AGEMA_signal_1444, n2588}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2719 ( .a ({new_AGEMA_signal_1105, n2594}), .b ({new_AGEMA_signal_3032, new_AGEMA_signal_3030}), .clk ( clk ), .r ( Fresh[417] ), .c ({new_AGEMA_signal_1279, n2607}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2722 ( .a ({new_AGEMA_signal_1117, n2597}), .b ({new_AGEMA_signal_1280, n2596}), .clk ( clk ), .r ( Fresh[418] ), .c ({new_AGEMA_signal_1445, n2605}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2724 ( .a ({new_AGEMA_signal_1281, n2598}), .b ({new_AGEMA_signal_3068, new_AGEMA_signal_3066}), .clk ( clk ), .r ( Fresh[419] ), .c ({new_AGEMA_signal_1446, n2603}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2726 ( .a ({new_AGEMA_signal_1021, n2599}), .b ({new_AGEMA_signal_2984, new_AGEMA_signal_2982}), .clk ( clk ), .r ( Fresh[420] ), .c ({new_AGEMA_signal_1118, n2601}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2733 ( .a ({new_AGEMA_signal_1283, n2610}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2966}), .clk ( clk ), .r ( Fresh[421] ), .c ({new_AGEMA_signal_1447, n2620}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2736 ( .a ({new_AGEMA_signal_1284, n2614}), .b ({new_AGEMA_signal_1285, n2613}), .clk ( clk ), .r ( Fresh[422] ), .c ({new_AGEMA_signal_1448, n2618}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2743 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ( Fresh[423] ), .c ({new_AGEMA_signal_1449, n2626}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2746 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2898}), .clk ( clk ), .r ( Fresh[424] ), .c ({new_AGEMA_signal_1286, n2632}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2752 ( .a ({new_AGEMA_signal_1287, n2784}), .b ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .r ( Fresh[425] ), .c ({new_AGEMA_signal_1450, n2644}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2754 ( .a ({new_AGEMA_signal_2824, new_AGEMA_signal_2822}), .b ({new_AGEMA_signal_1093, n2645}), .clk ( clk ), .r ( Fresh[426] ), .c ({new_AGEMA_signal_1288, n2646}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2758 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_1121, n2650}), .clk ( clk ), .r ( Fresh[427] ), .c ({new_AGEMA_signal_1289, n2653}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2760 ( .a ({new_AGEMA_signal_2984, new_AGEMA_signal_2982}), .b ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .r ( Fresh[428] ), .c ({new_AGEMA_signal_1452, n2655}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2764 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_2992, new_AGEMA_signal_2990}), .clk ( clk ), .r ( Fresh[429] ), .c ({new_AGEMA_signal_1453, n2663}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2770 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_2972, new_AGEMA_signal_2970}), .clk ( clk ), .r ( Fresh[430] ), .c ({new_AGEMA_signal_1290, n2675}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2772 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1043, n2676}), .clk ( clk ), .r ( Fresh[431] ), .c ({new_AGEMA_signal_1291, n2678}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2780 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_2988, new_AGEMA_signal_2986}), .clk ( clk ), .r ( Fresh[432] ), .c ({new_AGEMA_signal_1292, n2691}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2782 ( .a ({new_AGEMA_signal_3000, new_AGEMA_signal_2998}), .b ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .r ( Fresh[433] ), .c ({new_AGEMA_signal_1455, n2695}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2785 ( .a ({new_AGEMA_signal_1104, n2700}), .b ({new_AGEMA_signal_3064, new_AGEMA_signal_3062}), .clk ( clk ), .r ( Fresh[434] ), .c ({new_AGEMA_signal_1293, n2701}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2791 ( .a ({new_AGEMA_signal_1294, n2711}), .b ({new_AGEMA_signal_1295, n2710}), .clk ( clk ), .r ( Fresh[435] ), .c ({new_AGEMA_signal_1456, n2717}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2796 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_2948, new_AGEMA_signal_2946}), .clk ( clk ), .r ( Fresh[436] ), .c ({new_AGEMA_signal_1576, n2729}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2798 ( .a ({new_AGEMA_signal_2880, new_AGEMA_signal_2878}), .b ({new_AGEMA_signal_1123, n2722}), .clk ( clk ), .r ( Fresh[437] ), .c ({new_AGEMA_signal_1296, n2727}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2803 ( .a ({new_AGEMA_signal_1135, n2732}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ( Fresh[438] ), .c ({new_AGEMA_signal_1458, n2733}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2807 ( .a ({new_AGEMA_signal_3072, new_AGEMA_signal_3070}), .b ({new_AGEMA_signal_1298, n2738}), .clk ( clk ), .r ( Fresh[439] ), .c ({new_AGEMA_signal_1459, n2740}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2812 ( .a ({new_AGEMA_signal_1088, n2748}), .b ({new_AGEMA_signal_2808, new_AGEMA_signal_2806}), .clk ( clk ), .r ( Fresh[440] ), .c ({new_AGEMA_signal_1299, n2749}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2815 ( .a ({new_AGEMA_signal_1173, n2754}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2886}), .clk ( clk ), .r ( Fresh[441] ), .c ({new_AGEMA_signal_1461, n2757}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2816 ( .a ({new_AGEMA_signal_1030, n2755}), .b ({new_AGEMA_signal_3076, new_AGEMA_signal_3074}), .clk ( clk ), .r ( Fresh[442] ), .c ({new_AGEMA_signal_1300, n2756}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2819 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_3004, new_AGEMA_signal_3002}), .clk ( clk ), .r ( Fresh[443] ), .c ({new_AGEMA_signal_1462, n2762}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2823 ( .a ({new_AGEMA_signal_2808, new_AGEMA_signal_2806}), .b ({new_AGEMA_signal_1301, n2768}), .clk ( clk ), .r ( Fresh[444] ), .c ({new_AGEMA_signal_1463, n2770}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2825 ( .a ({new_AGEMA_signal_1184, n2773}), .b ({new_AGEMA_signal_3076, new_AGEMA_signal_3074}), .clk ( clk ), .r ( Fresh[445] ), .c ({new_AGEMA_signal_1464, n2776}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2826 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2810}), .clk ( clk ), .r ( Fresh[446] ), .c ({new_AGEMA_signal_1465, n2775}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2830 ( .a ({new_AGEMA_signal_1124, n2782}), .b ({new_AGEMA_signal_1125, n2781}), .clk ( clk ), .r ( Fresh[447] ), .c ({new_AGEMA_signal_1302, n2783}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2836 ( .a ({new_AGEMA_signal_1304, n2794}), .b ({new_AGEMA_signal_1305, n2793}), .clk ( clk ), .r ( Fresh[448] ), .c ({new_AGEMA_signal_1467, n2795}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2845 ( .a ({new_AGEMA_signal_1306, n2812}), .b ({new_AGEMA_signal_1194, n2811}), .clk ( clk ), .r ( Fresh[449] ), .c ({new_AGEMA_signal_1468, n2814}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2848 ( .a ({new_AGEMA_signal_2856, new_AGEMA_signal_2854}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[450] ), .c ({new_AGEMA_signal_1307, n2819}) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C ( clk ), .D ( new_AGEMA_signal_3077 ), .Q ( new_AGEMA_signal_3078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C ( clk ), .D ( new_AGEMA_signal_3079 ), .Q ( new_AGEMA_signal_3080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C ( clk ), .D ( new_AGEMA_signal_3081 ), .Q ( new_AGEMA_signal_3082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C ( clk ), .D ( new_AGEMA_signal_3083 ), .Q ( new_AGEMA_signal_3084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C ( clk ), .D ( new_AGEMA_signal_3087 ), .Q ( new_AGEMA_signal_3088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C ( clk ), .D ( new_AGEMA_signal_3091 ), .Q ( new_AGEMA_signal_3092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C ( clk ), .D ( new_AGEMA_signal_3093 ), .Q ( new_AGEMA_signal_3094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C ( clk ), .D ( new_AGEMA_signal_3095 ), .Q ( new_AGEMA_signal_3096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C ( clk ), .D ( new_AGEMA_signal_3097 ), .Q ( new_AGEMA_signal_3098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C ( clk ), .D ( new_AGEMA_signal_3099 ), .Q ( new_AGEMA_signal_3100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C ( clk ), .D ( new_AGEMA_signal_3101 ), .Q ( new_AGEMA_signal_3102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C ( clk ), .D ( new_AGEMA_signal_3103 ), .Q ( new_AGEMA_signal_3104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C ( clk ), .D ( new_AGEMA_signal_3105 ), .Q ( new_AGEMA_signal_3106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C ( clk ), .D ( new_AGEMA_signal_3107 ), .Q ( new_AGEMA_signal_3108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C ( clk ), .D ( new_AGEMA_signal_3109 ), .Q ( new_AGEMA_signal_3110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C ( clk ), .D ( new_AGEMA_signal_3111 ), .Q ( new_AGEMA_signal_3112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C ( clk ), .D ( new_AGEMA_signal_3113 ), .Q ( new_AGEMA_signal_3114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C ( clk ), .D ( new_AGEMA_signal_3115 ), .Q ( new_AGEMA_signal_3116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C ( clk ), .D ( new_AGEMA_signal_3117 ), .Q ( new_AGEMA_signal_3118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C ( clk ), .D ( new_AGEMA_signal_3119 ), .Q ( new_AGEMA_signal_3120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C ( clk ), .D ( new_AGEMA_signal_3121 ), .Q ( new_AGEMA_signal_3122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C ( clk ), .D ( new_AGEMA_signal_3123 ), .Q ( new_AGEMA_signal_3124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C ( clk ), .D ( new_AGEMA_signal_3125 ), .Q ( new_AGEMA_signal_3126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C ( clk ), .D ( new_AGEMA_signal_3127 ), .Q ( new_AGEMA_signal_3128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C ( clk ), .D ( new_AGEMA_signal_3129 ), .Q ( new_AGEMA_signal_3130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C ( clk ), .D ( new_AGEMA_signal_3131 ), .Q ( new_AGEMA_signal_3132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C ( clk ), .D ( new_AGEMA_signal_3133 ), .Q ( new_AGEMA_signal_3134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C ( clk ), .D ( new_AGEMA_signal_3135 ), .Q ( new_AGEMA_signal_3136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C ( clk ), .D ( new_AGEMA_signal_3139 ), .Q ( new_AGEMA_signal_3140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C ( clk ), .D ( new_AGEMA_signal_3143 ), .Q ( new_AGEMA_signal_3144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C ( clk ), .D ( new_AGEMA_signal_3145 ), .Q ( new_AGEMA_signal_3146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C ( clk ), .D ( new_AGEMA_signal_3147 ), .Q ( new_AGEMA_signal_3148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C ( clk ), .D ( new_AGEMA_signal_3149 ), .Q ( new_AGEMA_signal_3150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C ( clk ), .D ( new_AGEMA_signal_3151 ), .Q ( new_AGEMA_signal_3152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C ( clk ), .D ( new_AGEMA_signal_3153 ), .Q ( new_AGEMA_signal_3154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C ( clk ), .D ( new_AGEMA_signal_3155 ), .Q ( new_AGEMA_signal_3156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C ( clk ), .D ( new_AGEMA_signal_3157 ), .Q ( new_AGEMA_signal_3158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C ( clk ), .D ( new_AGEMA_signal_3159 ), .Q ( new_AGEMA_signal_3160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C ( clk ), .D ( new_AGEMA_signal_3161 ), .Q ( new_AGEMA_signal_3162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C ( clk ), .D ( new_AGEMA_signal_3163 ), .Q ( new_AGEMA_signal_3164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C ( clk ), .D ( new_AGEMA_signal_3165 ), .Q ( new_AGEMA_signal_3166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C ( clk ), .D ( new_AGEMA_signal_3167 ), .Q ( new_AGEMA_signal_3168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C ( clk ), .D ( new_AGEMA_signal_3169 ), .Q ( new_AGEMA_signal_3170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C ( clk ), .D ( new_AGEMA_signal_3171 ), .Q ( new_AGEMA_signal_3172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C ( clk ), .D ( new_AGEMA_signal_3175 ), .Q ( new_AGEMA_signal_3176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C ( clk ), .D ( new_AGEMA_signal_3179 ), .Q ( new_AGEMA_signal_3180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C ( clk ), .D ( new_AGEMA_signal_3181 ), .Q ( new_AGEMA_signal_3182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C ( clk ), .D ( new_AGEMA_signal_3183 ), .Q ( new_AGEMA_signal_3184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C ( clk ), .D ( new_AGEMA_signal_3185 ), .Q ( new_AGEMA_signal_3186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C ( clk ), .D ( new_AGEMA_signal_3187 ), .Q ( new_AGEMA_signal_3188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C ( clk ), .D ( new_AGEMA_signal_3189 ), .Q ( new_AGEMA_signal_3190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C ( clk ), .D ( new_AGEMA_signal_3191 ), .Q ( new_AGEMA_signal_3192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C ( clk ), .D ( new_AGEMA_signal_3193 ), .Q ( new_AGEMA_signal_3194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C ( clk ), .D ( new_AGEMA_signal_3195 ), .Q ( new_AGEMA_signal_3196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C ( clk ), .D ( new_AGEMA_signal_3197 ), .Q ( new_AGEMA_signal_3198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C ( clk ), .D ( new_AGEMA_signal_3199 ), .Q ( new_AGEMA_signal_3200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C ( clk ), .D ( new_AGEMA_signal_3203 ), .Q ( new_AGEMA_signal_3204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C ( clk ), .D ( new_AGEMA_signal_3207 ), .Q ( new_AGEMA_signal_3208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C ( clk ), .D ( new_AGEMA_signal_3209 ), .Q ( new_AGEMA_signal_3210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C ( clk ), .D ( new_AGEMA_signal_3211 ), .Q ( new_AGEMA_signal_3212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C ( clk ), .D ( new_AGEMA_signal_3213 ), .Q ( new_AGEMA_signal_3214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C ( clk ), .D ( new_AGEMA_signal_3215 ), .Q ( new_AGEMA_signal_3216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C ( clk ), .D ( new_AGEMA_signal_3217 ), .Q ( new_AGEMA_signal_3218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C ( clk ), .D ( new_AGEMA_signal_3219 ), .Q ( new_AGEMA_signal_3220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C ( clk ), .D ( new_AGEMA_signal_3223 ), .Q ( new_AGEMA_signal_3224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C ( clk ), .D ( new_AGEMA_signal_3227 ), .Q ( new_AGEMA_signal_3228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C ( clk ), .D ( new_AGEMA_signal_3229 ), .Q ( new_AGEMA_signal_3230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C ( clk ), .D ( new_AGEMA_signal_3231 ), .Q ( new_AGEMA_signal_3232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C ( clk ), .D ( new_AGEMA_signal_3233 ), .Q ( new_AGEMA_signal_3234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C ( clk ), .D ( new_AGEMA_signal_3235 ), .Q ( new_AGEMA_signal_3236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C ( clk ), .D ( new_AGEMA_signal_3237 ), .Q ( new_AGEMA_signal_3238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C ( clk ), .D ( new_AGEMA_signal_3239 ), .Q ( new_AGEMA_signal_3240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C ( clk ), .D ( new_AGEMA_signal_3243 ), .Q ( new_AGEMA_signal_3244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C ( clk ), .D ( new_AGEMA_signal_3247 ), .Q ( new_AGEMA_signal_3248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C ( clk ), .D ( new_AGEMA_signal_3249 ), .Q ( new_AGEMA_signal_3250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C ( clk ), .D ( new_AGEMA_signal_3251 ), .Q ( new_AGEMA_signal_3252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C ( clk ), .D ( new_AGEMA_signal_3253 ), .Q ( new_AGEMA_signal_3254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C ( clk ), .D ( new_AGEMA_signal_3255 ), .Q ( new_AGEMA_signal_3256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C ( clk ), .D ( new_AGEMA_signal_3257 ), .Q ( new_AGEMA_signal_3258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C ( clk ), .D ( new_AGEMA_signal_3259 ), .Q ( new_AGEMA_signal_3260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C ( clk ), .D ( new_AGEMA_signal_3261 ), .Q ( new_AGEMA_signal_3262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C ( clk ), .D ( new_AGEMA_signal_3263 ), .Q ( new_AGEMA_signal_3264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C ( clk ), .D ( new_AGEMA_signal_3265 ), .Q ( new_AGEMA_signal_3266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C ( clk ), .D ( new_AGEMA_signal_3267 ), .Q ( new_AGEMA_signal_3268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C ( clk ), .D ( new_AGEMA_signal_3269 ), .Q ( new_AGEMA_signal_3270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C ( clk ), .D ( new_AGEMA_signal_3271 ), .Q ( new_AGEMA_signal_3272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C ( clk ), .D ( new_AGEMA_signal_3273 ), .Q ( new_AGEMA_signal_3274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C ( clk ), .D ( new_AGEMA_signal_3275 ), .Q ( new_AGEMA_signal_3276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C ( clk ), .D ( new_AGEMA_signal_3277 ), .Q ( new_AGEMA_signal_3278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C ( clk ), .D ( new_AGEMA_signal_3279 ), .Q ( new_AGEMA_signal_3280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C ( clk ), .D ( new_AGEMA_signal_3281 ), .Q ( new_AGEMA_signal_3282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C ( clk ), .D ( new_AGEMA_signal_3283 ), .Q ( new_AGEMA_signal_3284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C ( clk ), .D ( new_AGEMA_signal_3285 ), .Q ( new_AGEMA_signal_3286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C ( clk ), .D ( new_AGEMA_signal_3287 ), .Q ( new_AGEMA_signal_3288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C ( clk ), .D ( new_AGEMA_signal_3289 ), .Q ( new_AGEMA_signal_3290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C ( clk ), .D ( new_AGEMA_signal_3291 ), .Q ( new_AGEMA_signal_3292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C ( clk ), .D ( new_AGEMA_signal_3293 ), .Q ( new_AGEMA_signal_3294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C ( clk ), .D ( new_AGEMA_signal_3295 ), .Q ( new_AGEMA_signal_3296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C ( clk ), .D ( new_AGEMA_signal_3297 ), .Q ( new_AGEMA_signal_3298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C ( clk ), .D ( new_AGEMA_signal_3299 ), .Q ( new_AGEMA_signal_3300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C ( clk ), .D ( new_AGEMA_signal_3301 ), .Q ( new_AGEMA_signal_3302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C ( clk ), .D ( new_AGEMA_signal_3303 ), .Q ( new_AGEMA_signal_3304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C ( clk ), .D ( new_AGEMA_signal_3305 ), .Q ( new_AGEMA_signal_3306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C ( clk ), .D ( new_AGEMA_signal_3307 ), .Q ( new_AGEMA_signal_3308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C ( clk ), .D ( new_AGEMA_signal_3309 ), .Q ( new_AGEMA_signal_3310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C ( clk ), .D ( new_AGEMA_signal_3311 ), .Q ( new_AGEMA_signal_3312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C ( clk ), .D ( new_AGEMA_signal_3313 ), .Q ( new_AGEMA_signal_3314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C ( clk ), .D ( new_AGEMA_signal_3315 ), .Q ( new_AGEMA_signal_3316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C ( clk ), .D ( new_AGEMA_signal_3321 ), .Q ( new_AGEMA_signal_3322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C ( clk ), .D ( new_AGEMA_signal_3327 ), .Q ( new_AGEMA_signal_3328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C ( clk ), .D ( new_AGEMA_signal_3329 ), .Q ( new_AGEMA_signal_3330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C ( clk ), .D ( new_AGEMA_signal_3331 ), .Q ( new_AGEMA_signal_3332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C ( clk ), .D ( new_AGEMA_signal_3333 ), .Q ( new_AGEMA_signal_3334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C ( clk ), .D ( new_AGEMA_signal_3335 ), .Q ( new_AGEMA_signal_3336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C ( clk ), .D ( new_AGEMA_signal_3337 ), .Q ( new_AGEMA_signal_3338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C ( clk ), .D ( new_AGEMA_signal_3339 ), .Q ( new_AGEMA_signal_3340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C ( clk ), .D ( new_AGEMA_signal_3343 ), .Q ( new_AGEMA_signal_3344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C ( clk ), .D ( new_AGEMA_signal_3347 ), .Q ( new_AGEMA_signal_3348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C ( clk ), .D ( new_AGEMA_signal_3349 ), .Q ( new_AGEMA_signal_3350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C ( clk ), .D ( new_AGEMA_signal_3351 ), .Q ( new_AGEMA_signal_3352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C ( clk ), .D ( new_AGEMA_signal_3353 ), .Q ( new_AGEMA_signal_3354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C ( clk ), .D ( new_AGEMA_signal_3355 ), .Q ( new_AGEMA_signal_3356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C ( clk ), .D ( new_AGEMA_signal_3357 ), .Q ( new_AGEMA_signal_3358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C ( clk ), .D ( new_AGEMA_signal_3359 ), .Q ( new_AGEMA_signal_3360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C ( clk ), .D ( new_AGEMA_signal_3363 ), .Q ( new_AGEMA_signal_3364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C ( clk ), .D ( new_AGEMA_signal_3367 ), .Q ( new_AGEMA_signal_3368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C ( clk ), .D ( new_AGEMA_signal_3369 ), .Q ( new_AGEMA_signal_3370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C ( clk ), .D ( new_AGEMA_signal_3371 ), .Q ( new_AGEMA_signal_3372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C ( clk ), .D ( new_AGEMA_signal_3373 ), .Q ( new_AGEMA_signal_3374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C ( clk ), .D ( new_AGEMA_signal_3375 ), .Q ( new_AGEMA_signal_3376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C ( clk ), .D ( new_AGEMA_signal_3377 ), .Q ( new_AGEMA_signal_3378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C ( clk ), .D ( new_AGEMA_signal_3379 ), .Q ( new_AGEMA_signal_3380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C ( clk ), .D ( new_AGEMA_signal_3381 ), .Q ( new_AGEMA_signal_3382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C ( clk ), .D ( new_AGEMA_signal_3383 ), .Q ( new_AGEMA_signal_3384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C ( clk ), .D ( new_AGEMA_signal_3385 ), .Q ( new_AGEMA_signal_3386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C ( clk ), .D ( new_AGEMA_signal_3387 ), .Q ( new_AGEMA_signal_3388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C ( clk ), .D ( new_AGEMA_signal_3389 ), .Q ( new_AGEMA_signal_3390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C ( clk ), .D ( new_AGEMA_signal_3391 ), .Q ( new_AGEMA_signal_3392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C ( clk ), .D ( new_AGEMA_signal_3393 ), .Q ( new_AGEMA_signal_3394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C ( clk ), .D ( new_AGEMA_signal_3395 ), .Q ( new_AGEMA_signal_3396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C ( clk ), .D ( new_AGEMA_signal_3399 ), .Q ( new_AGEMA_signal_3400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C ( clk ), .D ( new_AGEMA_signal_3403 ), .Q ( new_AGEMA_signal_3404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C ( clk ), .D ( new_AGEMA_signal_3405 ), .Q ( new_AGEMA_signal_3406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C ( clk ), .D ( new_AGEMA_signal_3407 ), .Q ( new_AGEMA_signal_3408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C ( clk ), .D ( new_AGEMA_signal_3409 ), .Q ( new_AGEMA_signal_3410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C ( clk ), .D ( new_AGEMA_signal_3411 ), .Q ( new_AGEMA_signal_3412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C ( clk ), .D ( new_AGEMA_signal_3415 ), .Q ( new_AGEMA_signal_3416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C ( clk ), .D ( new_AGEMA_signal_3419 ), .Q ( new_AGEMA_signal_3420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C ( clk ), .D ( new_AGEMA_signal_3421 ), .Q ( new_AGEMA_signal_3422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C ( clk ), .D ( new_AGEMA_signal_3423 ), .Q ( new_AGEMA_signal_3424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C ( clk ), .D ( new_AGEMA_signal_3425 ), .Q ( new_AGEMA_signal_3426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C ( clk ), .D ( new_AGEMA_signal_3429 ), .Q ( new_AGEMA_signal_3430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C ( clk ), .D ( new_AGEMA_signal_3433 ), .Q ( new_AGEMA_signal_3434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C ( clk ), .D ( new_AGEMA_signal_3437 ), .Q ( new_AGEMA_signal_3438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C ( clk ), .D ( new_AGEMA_signal_3449 ), .Q ( new_AGEMA_signal_3450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C ( clk ), .D ( new_AGEMA_signal_3453 ), .Q ( new_AGEMA_signal_3454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C ( clk ), .D ( new_AGEMA_signal_3461 ), .Q ( new_AGEMA_signal_3462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C ( clk ), .D ( new_AGEMA_signal_3465 ), .Q ( new_AGEMA_signal_3466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C ( clk ), .D ( new_AGEMA_signal_3473 ), .Q ( new_AGEMA_signal_3474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C ( clk ), .D ( new_AGEMA_signal_3477 ), .Q ( new_AGEMA_signal_3478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C ( clk ), .D ( new_AGEMA_signal_3481 ), .Q ( new_AGEMA_signal_3482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C ( clk ), .D ( new_AGEMA_signal_3485 ), .Q ( new_AGEMA_signal_3486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C ( clk ), .D ( new_AGEMA_signal_3505 ), .Q ( new_AGEMA_signal_3506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C ( clk ), .D ( new_AGEMA_signal_3509 ), .Q ( new_AGEMA_signal_3510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C ( clk ), .D ( new_AGEMA_signal_3513 ), .Q ( new_AGEMA_signal_3514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C ( clk ), .D ( new_AGEMA_signal_3517 ), .Q ( new_AGEMA_signal_3518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C ( clk ), .D ( new_AGEMA_signal_3521 ), .Q ( new_AGEMA_signal_3522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C ( clk ), .D ( new_AGEMA_signal_3525 ), .Q ( new_AGEMA_signal_3526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C ( clk ), .D ( new_AGEMA_signal_3541 ), .Q ( new_AGEMA_signal_3542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C ( clk ), .D ( new_AGEMA_signal_3545 ), .Q ( new_AGEMA_signal_3546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C ( clk ), .D ( new_AGEMA_signal_3553 ), .Q ( new_AGEMA_signal_3554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C ( clk ), .D ( new_AGEMA_signal_3557 ), .Q ( new_AGEMA_signal_3558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C ( clk ), .D ( new_AGEMA_signal_3563 ), .Q ( new_AGEMA_signal_3564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C ( clk ), .D ( new_AGEMA_signal_3569 ), .Q ( new_AGEMA_signal_3570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C ( clk ), .D ( new_AGEMA_signal_3573 ), .Q ( new_AGEMA_signal_3574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C ( clk ), .D ( new_AGEMA_signal_3577 ), .Q ( new_AGEMA_signal_3578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C ( clk ), .D ( new_AGEMA_signal_3581 ), .Q ( new_AGEMA_signal_3582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C ( clk ), .D ( new_AGEMA_signal_3585 ), .Q ( new_AGEMA_signal_3586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C ( clk ), .D ( new_AGEMA_signal_3605 ), .Q ( new_AGEMA_signal_3606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C ( clk ), .D ( new_AGEMA_signal_3609 ), .Q ( new_AGEMA_signal_3610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C ( clk ), .D ( new_AGEMA_signal_3615 ), .Q ( new_AGEMA_signal_3616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C ( clk ), .D ( new_AGEMA_signal_3621 ), .Q ( new_AGEMA_signal_3622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C ( clk ), .D ( new_AGEMA_signal_3625 ), .Q ( new_AGEMA_signal_3626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C ( clk ), .D ( new_AGEMA_signal_3629 ), .Q ( new_AGEMA_signal_3630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C ( clk ), .D ( new_AGEMA_signal_3645 ), .Q ( new_AGEMA_signal_3646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C ( clk ), .D ( new_AGEMA_signal_3649 ), .Q ( new_AGEMA_signal_3650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C ( clk ), .D ( new_AGEMA_signal_3661 ), .Q ( new_AGEMA_signal_3662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C ( clk ), .D ( new_AGEMA_signal_3665 ), .Q ( new_AGEMA_signal_3666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C ( clk ), .D ( new_AGEMA_signal_3669 ), .Q ( new_AGEMA_signal_3670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C ( clk ), .D ( new_AGEMA_signal_3673 ), .Q ( new_AGEMA_signal_3674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C ( clk ), .D ( new_AGEMA_signal_3677 ), .Q ( new_AGEMA_signal_3678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C ( clk ), .D ( new_AGEMA_signal_3681 ), .Q ( new_AGEMA_signal_3682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C ( clk ), .D ( new_AGEMA_signal_3685 ), .Q ( new_AGEMA_signal_3686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C ( clk ), .D ( new_AGEMA_signal_3689 ), .Q ( new_AGEMA_signal_3690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C ( clk ), .D ( new_AGEMA_signal_3693 ), .Q ( new_AGEMA_signal_3694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C ( clk ), .D ( new_AGEMA_signal_3697 ), .Q ( new_AGEMA_signal_3698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C ( clk ), .D ( new_AGEMA_signal_3717 ), .Q ( new_AGEMA_signal_3718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C ( clk ), .D ( new_AGEMA_signal_3721 ), .Q ( new_AGEMA_signal_3722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C ( clk ), .D ( new_AGEMA_signal_3725 ), .Q ( new_AGEMA_signal_3726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C ( clk ), .D ( new_AGEMA_signal_3729 ), .Q ( new_AGEMA_signal_3730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C ( clk ), .D ( new_AGEMA_signal_3769 ), .Q ( new_AGEMA_signal_3770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C ( clk ), .D ( new_AGEMA_signal_3773 ), .Q ( new_AGEMA_signal_3774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C ( clk ), .D ( new_AGEMA_signal_3797 ), .Q ( new_AGEMA_signal_3798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C ( clk ), .D ( new_AGEMA_signal_3801 ), .Q ( new_AGEMA_signal_3802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C ( clk ), .D ( new_AGEMA_signal_3805 ), .Q ( new_AGEMA_signal_3806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C ( clk ), .D ( new_AGEMA_signal_3809 ), .Q ( new_AGEMA_signal_3810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C ( clk ), .D ( new_AGEMA_signal_3813 ), .Q ( new_AGEMA_signal_3814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C ( clk ), .D ( new_AGEMA_signal_3817 ), .Q ( new_AGEMA_signal_3818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C ( clk ), .D ( new_AGEMA_signal_3821 ), .Q ( new_AGEMA_signal_3822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C ( clk ), .D ( new_AGEMA_signal_3825 ), .Q ( new_AGEMA_signal_3826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C ( clk ), .D ( new_AGEMA_signal_3847 ), .Q ( new_AGEMA_signal_3848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C ( clk ), .D ( new_AGEMA_signal_3855 ), .Q ( new_AGEMA_signal_3856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C ( clk ), .D ( new_AGEMA_signal_3867 ), .Q ( new_AGEMA_signal_3868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C ( clk ), .D ( new_AGEMA_signal_3875 ), .Q ( new_AGEMA_signal_3876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C ( clk ), .D ( new_AGEMA_signal_3881 ), .Q ( new_AGEMA_signal_3882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C ( clk ), .D ( new_AGEMA_signal_3887 ), .Q ( new_AGEMA_signal_3888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C ( clk ), .D ( new_AGEMA_signal_3901 ), .Q ( new_AGEMA_signal_3902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C ( clk ), .D ( new_AGEMA_signal_3907 ), .Q ( new_AGEMA_signal_3908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C ( clk ), .D ( new_AGEMA_signal_3917 ), .Q ( new_AGEMA_signal_3918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C ( clk ), .D ( new_AGEMA_signal_3923 ), .Q ( new_AGEMA_signal_3924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C ( clk ), .D ( new_AGEMA_signal_3929 ), .Q ( new_AGEMA_signal_3930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C ( clk ), .D ( new_AGEMA_signal_3935 ), .Q ( new_AGEMA_signal_3936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C ( clk ), .D ( new_AGEMA_signal_3953 ), .Q ( new_AGEMA_signal_3954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C ( clk ), .D ( new_AGEMA_signal_3959 ), .Q ( new_AGEMA_signal_3960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C ( clk ), .D ( new_AGEMA_signal_3965 ), .Q ( new_AGEMA_signal_3966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C ( clk ), .D ( new_AGEMA_signal_3971 ), .Q ( new_AGEMA_signal_3972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C ( clk ), .D ( new_AGEMA_signal_3981 ), .Q ( new_AGEMA_signal_3982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C ( clk ), .D ( new_AGEMA_signal_3987 ), .Q ( new_AGEMA_signal_3988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C ( clk ), .D ( new_AGEMA_signal_4019 ), .Q ( new_AGEMA_signal_4020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C ( clk ), .D ( new_AGEMA_signal_4027 ), .Q ( new_AGEMA_signal_4028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C ( clk ), .D ( new_AGEMA_signal_4033 ), .Q ( new_AGEMA_signal_4034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C ( clk ), .D ( new_AGEMA_signal_4039 ), .Q ( new_AGEMA_signal_4040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C ( clk ), .D ( new_AGEMA_signal_4089 ), .Q ( new_AGEMA_signal_4090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C ( clk ), .D ( new_AGEMA_signal_4095 ), .Q ( new_AGEMA_signal_4096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C ( clk ), .D ( new_AGEMA_signal_4153 ), .Q ( new_AGEMA_signal_4154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C ( clk ), .D ( new_AGEMA_signal_4159 ), .Q ( new_AGEMA_signal_4160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C ( clk ), .D ( new_AGEMA_signal_4165 ), .Q ( new_AGEMA_signal_4166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C ( clk ), .D ( new_AGEMA_signal_4171 ), .Q ( new_AGEMA_signal_4172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C ( clk ), .D ( new_AGEMA_signal_4191 ), .Q ( new_AGEMA_signal_4192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C ( clk ), .D ( new_AGEMA_signal_4199 ), .Q ( new_AGEMA_signal_4200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C ( clk ), .D ( new_AGEMA_signal_4251 ), .Q ( new_AGEMA_signal_4252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C ( clk ), .D ( new_AGEMA_signal_4259 ), .Q ( new_AGEMA_signal_4260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C ( clk ), .D ( new_AGEMA_signal_4281 ), .Q ( new_AGEMA_signal_4282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C ( clk ), .D ( new_AGEMA_signal_4287 ), .Q ( new_AGEMA_signal_4288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C ( clk ), .D ( new_AGEMA_signal_4297 ), .Q ( new_AGEMA_signal_4298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C ( clk ), .D ( new_AGEMA_signal_4305 ), .Q ( new_AGEMA_signal_4306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C ( clk ), .D ( new_AGEMA_signal_4325 ), .Q ( new_AGEMA_signal_4326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C ( clk ), .D ( new_AGEMA_signal_4333 ), .Q ( new_AGEMA_signal_4334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C ( clk ), .D ( new_AGEMA_signal_4365 ), .Q ( new_AGEMA_signal_4366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C ( clk ), .D ( new_AGEMA_signal_4373 ), .Q ( new_AGEMA_signal_4374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C ( clk ), .D ( new_AGEMA_signal_4457 ), .Q ( new_AGEMA_signal_4458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C ( clk ), .D ( new_AGEMA_signal_4465 ), .Q ( new_AGEMA_signal_4466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C ( clk ), .D ( new_AGEMA_signal_4493 ), .Q ( new_AGEMA_signal_4494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C ( clk ), .D ( new_AGEMA_signal_4501 ), .Q ( new_AGEMA_signal_4502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C ( clk ), .D ( new_AGEMA_signal_4557 ), .Q ( new_AGEMA_signal_4558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C ( clk ), .D ( new_AGEMA_signal_4565 ), .Q ( new_AGEMA_signal_4566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C ( clk ), .D ( new_AGEMA_signal_4573 ), .Q ( new_AGEMA_signal_4574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C ( clk ), .D ( new_AGEMA_signal_4581 ), .Q ( new_AGEMA_signal_4582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C ( clk ), .D ( new_AGEMA_signal_4745 ), .Q ( new_AGEMA_signal_4746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C ( clk ), .D ( new_AGEMA_signal_4755 ), .Q ( new_AGEMA_signal_4756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C ( clk ), .D ( new_AGEMA_signal_4845 ), .Q ( new_AGEMA_signal_4846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C ( clk ), .D ( new_AGEMA_signal_4855 ), .Q ( new_AGEMA_signal_4856 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_1609 ( .C ( clk ), .D ( new_AGEMA_signal_3426 ), .Q ( new_AGEMA_signal_3427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C ( clk ), .D ( new_AGEMA_signal_3430 ), .Q ( new_AGEMA_signal_3431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C ( clk ), .D ( new_AGEMA_signal_3434 ), .Q ( new_AGEMA_signal_3435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C ( clk ), .D ( new_AGEMA_signal_3438 ), .Q ( new_AGEMA_signal_3439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C ( clk ), .D ( new_AGEMA_signal_3350 ), .Q ( new_AGEMA_signal_3441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C ( clk ), .D ( new_AGEMA_signal_3352 ), .Q ( new_AGEMA_signal_3443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C ( clk ), .D ( n1966 ), .Q ( new_AGEMA_signal_3445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C ( clk ), .D ( new_AGEMA_signal_1321 ), .Q ( new_AGEMA_signal_3447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C ( clk ), .D ( new_AGEMA_signal_3450 ), .Q ( new_AGEMA_signal_3451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C ( clk ), .D ( new_AGEMA_signal_3454 ), .Q ( new_AGEMA_signal_3455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C ( clk ), .D ( new_AGEMA_signal_3278 ), .Q ( new_AGEMA_signal_3457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C ( clk ), .D ( new_AGEMA_signal_3280 ), .Q ( new_AGEMA_signal_3459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C ( clk ), .D ( new_AGEMA_signal_3462 ), .Q ( new_AGEMA_signal_3463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C ( clk ), .D ( new_AGEMA_signal_3466 ), .Q ( new_AGEMA_signal_3467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C ( clk ), .D ( n1996 ), .Q ( new_AGEMA_signal_3469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C ( clk ), .D ( new_AGEMA_signal_1331 ), .Q ( new_AGEMA_signal_3471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C ( clk ), .D ( new_AGEMA_signal_3474 ), .Q ( new_AGEMA_signal_3475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C ( clk ), .D ( new_AGEMA_signal_3478 ), .Q ( new_AGEMA_signal_3479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C ( clk ), .D ( new_AGEMA_signal_3482 ), .Q ( new_AGEMA_signal_3483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C ( clk ), .D ( new_AGEMA_signal_3486 ), .Q ( new_AGEMA_signal_3487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C ( clk ), .D ( n2033 ), .Q ( new_AGEMA_signal_3489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C ( clk ), .D ( new_AGEMA_signal_1337 ), .Q ( new_AGEMA_signal_3491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C ( clk ), .D ( new_AGEMA_signal_3190 ), .Q ( new_AGEMA_signal_3493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C ( clk ), .D ( new_AGEMA_signal_3192 ), .Q ( new_AGEMA_signal_3495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C ( clk ), .D ( new_AGEMA_signal_3210 ), .Q ( new_AGEMA_signal_3497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C ( clk ), .D ( new_AGEMA_signal_3212 ), .Q ( new_AGEMA_signal_3499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C ( clk ), .D ( new_AGEMA_signal_3266 ), .Q ( new_AGEMA_signal_3501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C ( clk ), .D ( new_AGEMA_signal_3268 ), .Q ( new_AGEMA_signal_3503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C ( clk ), .D ( new_AGEMA_signal_3506 ), .Q ( new_AGEMA_signal_3507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C ( clk ), .D ( new_AGEMA_signal_3510 ), .Q ( new_AGEMA_signal_3511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C ( clk ), .D ( new_AGEMA_signal_3514 ), .Q ( new_AGEMA_signal_3515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C ( clk ), .D ( new_AGEMA_signal_3518 ), .Q ( new_AGEMA_signal_3519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C ( clk ), .D ( new_AGEMA_signal_3522 ), .Q ( new_AGEMA_signal_3523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C ( clk ), .D ( new_AGEMA_signal_3526 ), .Q ( new_AGEMA_signal_3527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C ( clk ), .D ( n2089 ), .Q ( new_AGEMA_signal_3529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C ( clk ), .D ( new_AGEMA_signal_1352 ), .Q ( new_AGEMA_signal_3531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C ( clk ), .D ( n2092 ), .Q ( new_AGEMA_signal_3533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_3535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C ( clk ), .D ( n2115 ), .Q ( new_AGEMA_signal_3537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C ( clk ), .D ( new_AGEMA_signal_1190 ), .Q ( new_AGEMA_signal_3539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C ( clk ), .D ( new_AGEMA_signal_3542 ), .Q ( new_AGEMA_signal_3543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C ( clk ), .D ( new_AGEMA_signal_3546 ), .Q ( new_AGEMA_signal_3547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C ( clk ), .D ( n2687 ), .Q ( new_AGEMA_signal_3549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C ( clk ), .D ( new_AGEMA_signal_1320 ), .Q ( new_AGEMA_signal_3551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C ( clk ), .D ( new_AGEMA_signal_3554 ), .Q ( new_AGEMA_signal_3555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C ( clk ), .D ( new_AGEMA_signal_3558 ), .Q ( new_AGEMA_signal_3559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C ( clk ), .D ( new_AGEMA_signal_3564 ), .Q ( new_AGEMA_signal_3565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C ( clk ), .D ( new_AGEMA_signal_3570 ), .Q ( new_AGEMA_signal_3571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C ( clk ), .D ( new_AGEMA_signal_3574 ), .Q ( new_AGEMA_signal_3575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C ( clk ), .D ( new_AGEMA_signal_3578 ), .Q ( new_AGEMA_signal_3579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C ( clk ), .D ( new_AGEMA_signal_3582 ), .Q ( new_AGEMA_signal_3583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C ( clk ), .D ( new_AGEMA_signal_3586 ), .Q ( new_AGEMA_signal_3587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C ( clk ), .D ( n2193 ), .Q ( new_AGEMA_signal_3589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_3591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C ( clk ), .D ( n2202 ), .Q ( new_AGEMA_signal_3593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C ( clk ), .D ( new_AGEMA_signal_1516 ), .Q ( new_AGEMA_signal_3595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C ( clk ), .D ( n2228 ), .Q ( new_AGEMA_signal_3597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C ( clk ), .D ( new_AGEMA_signal_1214 ), .Q ( new_AGEMA_signal_3599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C ( clk ), .D ( n2235 ), .Q ( new_AGEMA_signal_3601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C ( clk ), .D ( new_AGEMA_signal_1315 ), .Q ( new_AGEMA_signal_3603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C ( clk ), .D ( new_AGEMA_signal_3606 ), .Q ( new_AGEMA_signal_3607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C ( clk ), .D ( new_AGEMA_signal_3610 ), .Q ( new_AGEMA_signal_3611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C ( clk ), .D ( new_AGEMA_signal_3616 ), .Q ( new_AGEMA_signal_3617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C ( clk ), .D ( new_AGEMA_signal_3622 ), .Q ( new_AGEMA_signal_3623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C ( clk ), .D ( new_AGEMA_signal_3626 ), .Q ( new_AGEMA_signal_3627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C ( clk ), .D ( new_AGEMA_signal_3630 ), .Q ( new_AGEMA_signal_3631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C ( clk ), .D ( n2752 ), .Q ( new_AGEMA_signal_3633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C ( clk ), .D ( new_AGEMA_signal_1525 ), .Q ( new_AGEMA_signal_3635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C ( clk ), .D ( new_AGEMA_signal_3322 ), .Q ( new_AGEMA_signal_3637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C ( clk ), .D ( new_AGEMA_signal_3328 ), .Q ( new_AGEMA_signal_3639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C ( clk ), .D ( n2293 ), .Q ( new_AGEMA_signal_3641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C ( clk ), .D ( new_AGEMA_signal_1393 ), .Q ( new_AGEMA_signal_3643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C ( clk ), .D ( new_AGEMA_signal_3646 ), .Q ( new_AGEMA_signal_3647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C ( clk ), .D ( new_AGEMA_signal_3650 ), .Q ( new_AGEMA_signal_3651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C ( clk ), .D ( n2357 ), .Q ( new_AGEMA_signal_3653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C ( clk ), .D ( new_AGEMA_signal_1402 ), .Q ( new_AGEMA_signal_3655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C ( clk ), .D ( n2386 ), .Q ( new_AGEMA_signal_3657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C ( clk ), .D ( new_AGEMA_signal_1407 ), .Q ( new_AGEMA_signal_3659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C ( clk ), .D ( new_AGEMA_signal_3662 ), .Q ( new_AGEMA_signal_3663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C ( clk ), .D ( new_AGEMA_signal_3666 ), .Q ( new_AGEMA_signal_3667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C ( clk ), .D ( new_AGEMA_signal_3670 ), .Q ( new_AGEMA_signal_3671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C ( clk ), .D ( new_AGEMA_signal_3674 ), .Q ( new_AGEMA_signal_3675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C ( clk ), .D ( new_AGEMA_signal_3678 ), .Q ( new_AGEMA_signal_3679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C ( clk ), .D ( new_AGEMA_signal_3682 ), .Q ( new_AGEMA_signal_3683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C ( clk ), .D ( new_AGEMA_signal_3686 ), .Q ( new_AGEMA_signal_3687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C ( clk ), .D ( new_AGEMA_signal_3690 ), .Q ( new_AGEMA_signal_3691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C ( clk ), .D ( new_AGEMA_signal_3694 ), .Q ( new_AGEMA_signal_3695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C ( clk ), .D ( new_AGEMA_signal_3698 ), .Q ( new_AGEMA_signal_3699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C ( clk ), .D ( n2433 ), .Q ( new_AGEMA_signal_3701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C ( clk ), .D ( new_AGEMA_signal_1414 ), .Q ( new_AGEMA_signal_3703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C ( clk ), .D ( new_AGEMA_signal_3204 ), .Q ( new_AGEMA_signal_3705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C ( clk ), .D ( new_AGEMA_signal_3208 ), .Q ( new_AGEMA_signal_3707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C ( clk ), .D ( n2459 ), .Q ( new_AGEMA_signal_3709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C ( clk ), .D ( new_AGEMA_signal_1390 ), .Q ( new_AGEMA_signal_3711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C ( clk ), .D ( n2467 ), .Q ( new_AGEMA_signal_3713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C ( clk ), .D ( new_AGEMA_signal_1246 ), .Q ( new_AGEMA_signal_3715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C ( clk ), .D ( new_AGEMA_signal_3718 ), .Q ( new_AGEMA_signal_3719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C ( clk ), .D ( new_AGEMA_signal_3722 ), .Q ( new_AGEMA_signal_3723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C ( clk ), .D ( new_AGEMA_signal_3726 ), .Q ( new_AGEMA_signal_3727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C ( clk ), .D ( new_AGEMA_signal_3730 ), .Q ( new_AGEMA_signal_3731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C ( clk ), .D ( n2489 ), .Q ( new_AGEMA_signal_3733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C ( clk ), .D ( new_AGEMA_signal_1266 ), .Q ( new_AGEMA_signal_3735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C ( clk ), .D ( n2497 ), .Q ( new_AGEMA_signal_3737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C ( clk ), .D ( new_AGEMA_signal_1267 ), .Q ( new_AGEMA_signal_3739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C ( clk ), .D ( n2506 ), .Q ( new_AGEMA_signal_3741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C ( clk ), .D ( new_AGEMA_signal_1427 ), .Q ( new_AGEMA_signal_3743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C ( clk ), .D ( n2542 ), .Q ( new_AGEMA_signal_3745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C ( clk ), .D ( new_AGEMA_signal_1433 ), .Q ( new_AGEMA_signal_3747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C ( clk ), .D ( n2558 ), .Q ( new_AGEMA_signal_3749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C ( clk ), .D ( new_AGEMA_signal_1436 ), .Q ( new_AGEMA_signal_3751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C ( clk ), .D ( n2566 ), .Q ( new_AGEMA_signal_3753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_3755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C ( clk ), .D ( n2581 ), .Q ( new_AGEMA_signal_3757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C ( clk ), .D ( new_AGEMA_signal_1276 ), .Q ( new_AGEMA_signal_3759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C ( clk ), .D ( n2603 ), .Q ( new_AGEMA_signal_3761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_3763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C ( clk ), .D ( n2620 ), .Q ( new_AGEMA_signal_3765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C ( clk ), .D ( new_AGEMA_signal_1447 ), .Q ( new_AGEMA_signal_3767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C ( clk ), .D ( new_AGEMA_signal_3770 ), .Q ( new_AGEMA_signal_3771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C ( clk ), .D ( new_AGEMA_signal_3774 ), .Q ( new_AGEMA_signal_3775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C ( clk ), .D ( n2653 ), .Q ( new_AGEMA_signal_3777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C ( clk ), .D ( new_AGEMA_signal_1289 ), .Q ( new_AGEMA_signal_3779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C ( clk ), .D ( n2665 ), .Q ( new_AGEMA_signal_3781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C ( clk ), .D ( new_AGEMA_signal_1313 ), .Q ( new_AGEMA_signal_3783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C ( clk ), .D ( n2691 ), .Q ( new_AGEMA_signal_3785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C ( clk ), .D ( new_AGEMA_signal_1292 ), .Q ( new_AGEMA_signal_3787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C ( clk ), .D ( n2717 ), .Q ( new_AGEMA_signal_3789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C ( clk ), .D ( new_AGEMA_signal_1456 ), .Q ( new_AGEMA_signal_3791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C ( clk ), .D ( n2729 ), .Q ( new_AGEMA_signal_3793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C ( clk ), .D ( new_AGEMA_signal_1576 ), .Q ( new_AGEMA_signal_3795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C ( clk ), .D ( new_AGEMA_signal_3798 ), .Q ( new_AGEMA_signal_3799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C ( clk ), .D ( new_AGEMA_signal_3802 ), .Q ( new_AGEMA_signal_3803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C ( clk ), .D ( new_AGEMA_signal_3806 ), .Q ( new_AGEMA_signal_3807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C ( clk ), .D ( new_AGEMA_signal_3810 ), .Q ( new_AGEMA_signal_3811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C ( clk ), .D ( new_AGEMA_signal_3814 ), .Q ( new_AGEMA_signal_3815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C ( clk ), .D ( new_AGEMA_signal_3818 ), .Q ( new_AGEMA_signal_3819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C ( clk ), .D ( new_AGEMA_signal_3822 ), .Q ( new_AGEMA_signal_3823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C ( clk ), .D ( new_AGEMA_signal_3826 ), .Q ( new_AGEMA_signal_3827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C ( clk ), .D ( new_AGEMA_signal_3294 ), .Q ( new_AGEMA_signal_3829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C ( clk ), .D ( new_AGEMA_signal_3296 ), .Q ( new_AGEMA_signal_3833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C ( clk ), .D ( n1956 ), .Q ( new_AGEMA_signal_3837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C ( clk ), .D ( new_AGEMA_signal_1317 ), .Q ( new_AGEMA_signal_3841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C ( clk ), .D ( new_AGEMA_signal_3848 ), .Q ( new_AGEMA_signal_3849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C ( clk ), .D ( new_AGEMA_signal_3856 ), .Q ( new_AGEMA_signal_3857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C ( clk ), .D ( new_AGEMA_signal_3868 ), .Q ( new_AGEMA_signal_3869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C ( clk ), .D ( new_AGEMA_signal_3876 ), .Q ( new_AGEMA_signal_3877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C ( clk ), .D ( new_AGEMA_signal_3882 ), .Q ( new_AGEMA_signal_3883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C ( clk ), .D ( new_AGEMA_signal_3888 ), .Q ( new_AGEMA_signal_3889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C ( clk ), .D ( n2023 ), .Q ( new_AGEMA_signal_3893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C ( clk ), .D ( new_AGEMA_signal_1166 ), .Q ( new_AGEMA_signal_3897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C ( clk ), .D ( new_AGEMA_signal_3902 ), .Q ( new_AGEMA_signal_3903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C ( clk ), .D ( new_AGEMA_signal_3908 ), .Q ( new_AGEMA_signal_3909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C ( clk ), .D ( new_AGEMA_signal_3918 ), .Q ( new_AGEMA_signal_3919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C ( clk ), .D ( new_AGEMA_signal_3924 ), .Q ( new_AGEMA_signal_3925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C ( clk ), .D ( new_AGEMA_signal_3930 ), .Q ( new_AGEMA_signal_3931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C ( clk ), .D ( new_AGEMA_signal_3936 ), .Q ( new_AGEMA_signal_3937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C ( clk ), .D ( n2094 ), .Q ( new_AGEMA_signal_3945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C ( clk ), .D ( new_AGEMA_signal_1355 ), .Q ( new_AGEMA_signal_3949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C ( clk ), .D ( new_AGEMA_signal_3954 ), .Q ( new_AGEMA_signal_3955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C ( clk ), .D ( new_AGEMA_signal_3960 ), .Q ( new_AGEMA_signal_3961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C ( clk ), .D ( new_AGEMA_signal_3966 ), .Q ( new_AGEMA_signal_3967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C ( clk ), .D ( new_AGEMA_signal_3972 ), .Q ( new_AGEMA_signal_3973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C ( clk ), .D ( new_AGEMA_signal_3982 ), .Q ( new_AGEMA_signal_3983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C ( clk ), .D ( new_AGEMA_signal_3988 ), .Q ( new_AGEMA_signal_3989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C ( clk ), .D ( n2181 ), .Q ( new_AGEMA_signal_3997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C ( clk ), .D ( new_AGEMA_signal_1369 ), .Q ( new_AGEMA_signal_4001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C ( clk ), .D ( n2195 ), .Q ( new_AGEMA_signal_4005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C ( clk ), .D ( new_AGEMA_signal_1371 ), .Q ( new_AGEMA_signal_4009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C ( clk ), .D ( new_AGEMA_signal_4020 ), .Q ( new_AGEMA_signal_4021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C ( clk ), .D ( new_AGEMA_signal_4028 ), .Q ( new_AGEMA_signal_4029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C ( clk ), .D ( new_AGEMA_signal_4034 ), .Q ( new_AGEMA_signal_4035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C ( clk ), .D ( new_AGEMA_signal_4040 ), .Q ( new_AGEMA_signal_4041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C ( clk ), .D ( n2237 ), .Q ( new_AGEMA_signal_4045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C ( clk ), .D ( new_AGEMA_signal_1215 ), .Q ( new_AGEMA_signal_4049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C ( clk ), .D ( n2248 ), .Q ( new_AGEMA_signal_4053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C ( clk ), .D ( new_AGEMA_signal_1380 ), .Q ( new_AGEMA_signal_4057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C ( clk ), .D ( n2294 ), .Q ( new_AGEMA_signal_4069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C ( clk ), .D ( new_AGEMA_signal_1230 ), .Q ( new_AGEMA_signal_4073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C ( clk ), .D ( n2323 ), .Q ( new_AGEMA_signal_4077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C ( clk ), .D ( new_AGEMA_signal_1395 ), .Q ( new_AGEMA_signal_4081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C ( clk ), .D ( new_AGEMA_signal_4090 ), .Q ( new_AGEMA_signal_4091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C ( clk ), .D ( new_AGEMA_signal_4096 ), .Q ( new_AGEMA_signal_4097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C ( clk ), .D ( n2360 ), .Q ( new_AGEMA_signal_4101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C ( clk ), .D ( new_AGEMA_signal_1403 ), .Q ( new_AGEMA_signal_4105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C ( clk ), .D ( n2394 ), .Q ( new_AGEMA_signal_4113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C ( clk ), .D ( new_AGEMA_signal_1249 ), .Q ( new_AGEMA_signal_4117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C ( clk ), .D ( n2406 ), .Q ( new_AGEMA_signal_4121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C ( clk ), .D ( new_AGEMA_signal_1409 ), .Q ( new_AGEMA_signal_4125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C ( clk ), .D ( new_AGEMA_signal_3094 ), .Q ( new_AGEMA_signal_4129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C ( clk ), .D ( new_AGEMA_signal_3096 ), .Q ( new_AGEMA_signal_4133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C ( clk ), .D ( new_AGEMA_signal_3098 ), .Q ( new_AGEMA_signal_4141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C ( clk ), .D ( new_AGEMA_signal_3100 ), .Q ( new_AGEMA_signal_4145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C ( clk ), .D ( new_AGEMA_signal_4154 ), .Q ( new_AGEMA_signal_4155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C ( clk ), .D ( new_AGEMA_signal_4160 ), .Q ( new_AGEMA_signal_4161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C ( clk ), .D ( new_AGEMA_signal_4166 ), .Q ( new_AGEMA_signal_4167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C ( clk ), .D ( new_AGEMA_signal_4172 ), .Q ( new_AGEMA_signal_4173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C ( clk ), .D ( n2499 ), .Q ( new_AGEMA_signal_4177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C ( clk ), .D ( new_AGEMA_signal_1269 ), .Q ( new_AGEMA_signal_4181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C ( clk ), .D ( new_AGEMA_signal_4192 ), .Q ( new_AGEMA_signal_4193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C ( clk ), .D ( new_AGEMA_signal_4200 ), .Q ( new_AGEMA_signal_4201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C ( clk ), .D ( n2582 ), .Q ( new_AGEMA_signal_4209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C ( clk ), .D ( new_AGEMA_signal_1443 ), .Q ( new_AGEMA_signal_4213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C ( clk ), .D ( n2605 ), .Q ( new_AGEMA_signal_4217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C ( clk ), .D ( new_AGEMA_signal_1445 ), .Q ( new_AGEMA_signal_4221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C ( clk ), .D ( n2632 ), .Q ( new_AGEMA_signal_4225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C ( clk ), .D ( new_AGEMA_signal_1286 ), .Q ( new_AGEMA_signal_4229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C ( clk ), .D ( n2655 ), .Q ( new_AGEMA_signal_4233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C ( clk ), .D ( new_AGEMA_signal_1452 ), .Q ( new_AGEMA_signal_4237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C ( clk ), .D ( n2695 ), .Q ( new_AGEMA_signal_4241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C ( clk ), .D ( new_AGEMA_signal_1455 ), .Q ( new_AGEMA_signal_4245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C ( clk ), .D ( new_AGEMA_signal_4252 ), .Q ( new_AGEMA_signal_4253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C ( clk ), .D ( new_AGEMA_signal_4260 ), .Q ( new_AGEMA_signal_4261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C ( clk ), .D ( n2770 ), .Q ( new_AGEMA_signal_4269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C ( clk ), .D ( new_AGEMA_signal_1463 ), .Q ( new_AGEMA_signal_4273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C ( clk ), .D ( new_AGEMA_signal_4282 ), .Q ( new_AGEMA_signal_4283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C ( clk ), .D ( new_AGEMA_signal_4288 ), .Q ( new_AGEMA_signal_4289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C ( clk ), .D ( new_AGEMA_signal_4298 ), .Q ( new_AGEMA_signal_4299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C ( clk ), .D ( new_AGEMA_signal_4306 ), .Q ( new_AGEMA_signal_4307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C ( clk ), .D ( new_AGEMA_signal_4326 ), .Q ( new_AGEMA_signal_4327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C ( clk ), .D ( new_AGEMA_signal_4334 ), .Q ( new_AGEMA_signal_4335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C ( clk ), .D ( n2050 ), .Q ( new_AGEMA_signal_4345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C ( clk ), .D ( new_AGEMA_signal_1171 ), .Q ( new_AGEMA_signal_4351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C ( clk ), .D ( new_AGEMA_signal_4366 ), .Q ( new_AGEMA_signal_4367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C ( clk ), .D ( new_AGEMA_signal_4374 ), .Q ( new_AGEMA_signal_4375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C ( clk ), .D ( n2183 ), .Q ( new_AGEMA_signal_4389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C ( clk ), .D ( new_AGEMA_signal_1086 ), .Q ( new_AGEMA_signal_4395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C ( clk ), .D ( n2196 ), .Q ( new_AGEMA_signal_4401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C ( clk ), .D ( new_AGEMA_signal_1209 ), .Q ( new_AGEMA_signal_4407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C ( clk ), .D ( n2238 ), .Q ( new_AGEMA_signal_4413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C ( clk ), .D ( new_AGEMA_signal_1216 ), .Q ( new_AGEMA_signal_4419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C ( clk ), .D ( n2249 ), .Q ( new_AGEMA_signal_4425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C ( clk ), .D ( new_AGEMA_signal_1382 ), .Q ( new_AGEMA_signal_4431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C ( clk ), .D ( n2273 ), .Q ( new_AGEMA_signal_4437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C ( clk ), .D ( new_AGEMA_signal_1524 ), .Q ( new_AGEMA_signal_4443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C ( clk ), .D ( new_AGEMA_signal_4458 ), .Q ( new_AGEMA_signal_4459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C ( clk ), .D ( new_AGEMA_signal_4466 ), .Q ( new_AGEMA_signal_4467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C ( clk ), .D ( n2349 ), .Q ( new_AGEMA_signal_4481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C ( clk ), .D ( new_AGEMA_signal_1240 ), .Q ( new_AGEMA_signal_4487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C ( clk ), .D ( new_AGEMA_signal_4494 ), .Q ( new_AGEMA_signal_4495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C ( clk ), .D ( new_AGEMA_signal_4502 ), .Q ( new_AGEMA_signal_4503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C ( clk ), .D ( n2396 ), .Q ( new_AGEMA_signal_4513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C ( clk ), .D ( new_AGEMA_signal_1251 ), .Q ( new_AGEMA_signal_4519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C ( clk ), .D ( n2439 ), .Q ( new_AGEMA_signal_4533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C ( clk ), .D ( new_AGEMA_signal_1417 ), .Q ( new_AGEMA_signal_4539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C ( clk ), .D ( n2470 ), .Q ( new_AGEMA_signal_4545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C ( clk ), .D ( new_AGEMA_signal_1261 ), .Q ( new_AGEMA_signal_4551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C ( clk ), .D ( new_AGEMA_signal_4558 ), .Q ( new_AGEMA_signal_4559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C ( clk ), .D ( new_AGEMA_signal_4566 ), .Q ( new_AGEMA_signal_4567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C ( clk ), .D ( new_AGEMA_signal_4574 ), .Q ( new_AGEMA_signal_4575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C ( clk ), .D ( new_AGEMA_signal_4582 ), .Q ( new_AGEMA_signal_4583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C ( clk ), .D ( n2585 ), .Q ( new_AGEMA_signal_4589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C ( clk ), .D ( new_AGEMA_signal_1441 ), .Q ( new_AGEMA_signal_4595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C ( clk ), .D ( n2607 ), .Q ( new_AGEMA_signal_4601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C ( clk ), .D ( new_AGEMA_signal_1279 ), .Q ( new_AGEMA_signal_4607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C ( clk ), .D ( n2013 ), .Q ( new_AGEMA_signal_4669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C ( clk ), .D ( new_AGEMA_signal_1335 ), .Q ( new_AGEMA_signal_4677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C ( clk ), .D ( n2028 ), .Q ( new_AGEMA_signal_4685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C ( clk ), .D ( new_AGEMA_signal_1071 ), .Q ( new_AGEMA_signal_4693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C ( clk ), .D ( n2051 ), .Q ( new_AGEMA_signal_4701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C ( clk ), .D ( new_AGEMA_signal_1341 ), .Q ( new_AGEMA_signal_4709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C ( clk ), .D ( n2069 ), .Q ( new_AGEMA_signal_4717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C ( clk ), .D ( new_AGEMA_signal_1346 ), .Q ( new_AGEMA_signal_4725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C ( clk ), .D ( new_AGEMA_signal_4746 ), .Q ( new_AGEMA_signal_4747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C ( clk ), .D ( new_AGEMA_signal_4756 ), .Q ( new_AGEMA_signal_4757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C ( clk ), .D ( n2144 ), .Q ( new_AGEMA_signal_4765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C ( clk ), .D ( new_AGEMA_signal_1363 ), .Q ( new_AGEMA_signal_4773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C ( clk ), .D ( n2170 ), .Q ( new_AGEMA_signal_4781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C ( clk ), .D ( new_AGEMA_signal_1365 ), .Q ( new_AGEMA_signal_4789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C ( clk ), .D ( n2186 ), .Q ( new_AGEMA_signal_4797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_4805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C ( clk ), .D ( new_AGEMA_signal_4846 ), .Q ( new_AGEMA_signal_4847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C ( clk ), .D ( new_AGEMA_signal_4856 ), .Q ( new_AGEMA_signal_4857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C ( clk ), .D ( new_AGEMA_signal_3354 ), .Q ( new_AGEMA_signal_4865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C ( clk ), .D ( new_AGEMA_signal_3356 ), .Q ( new_AGEMA_signal_4873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C ( clk ), .D ( n2551 ), .Q ( new_AGEMA_signal_4893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C ( clk ), .D ( new_AGEMA_signal_1435 ), .Q ( new_AGEMA_signal_4901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C ( clk ), .D ( n2588 ), .Q ( new_AGEMA_signal_4909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C ( clk ), .D ( new_AGEMA_signal_1444 ), .Q ( new_AGEMA_signal_4917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C ( clk ), .D ( n2701 ), .Q ( new_AGEMA_signal_4945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C ( clk ), .D ( new_AGEMA_signal_1293 ), .Q ( new_AGEMA_signal_4953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C ( clk ), .D ( n2172 ), .Q ( new_AGEMA_signal_5077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C ( clk ), .D ( new_AGEMA_signal_1368 ), .Q ( new_AGEMA_signal_5087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C ( clk ), .D ( n2150 ), .Q ( new_AGEMA_signal_5469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C ( clk ), .D ( new_AGEMA_signal_1197 ), .Q ( new_AGEMA_signal_5483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C ( clk ), .D ( n2369 ), .Q ( new_AGEMA_signal_5513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C ( clk ), .D ( new_AGEMA_signal_1540 ), .Q ( new_AGEMA_signal_5527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C ( clk ), .D ( n2152 ), .Q ( new_AGEMA_signal_5585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C ( clk ), .D ( new_AGEMA_signal_1364 ), .Q ( new_AGEMA_signal_5601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C ( clk ), .D ( n2372 ), .Q ( new_AGEMA_signal_5629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C ( clk ), .D ( new_AGEMA_signal_1404 ), .Q ( new_AGEMA_signal_5645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C ( clk ), .D ( n2375 ), .Q ( new_AGEMA_signal_5781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C ( clk ), .D ( new_AGEMA_signal_1241 ), .Q ( new_AGEMA_signal_5799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C ( clk ), .D ( n2377 ), .Q ( new_AGEMA_signal_5881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C ( clk ), .D ( new_AGEMA_signal_1405 ), .Q ( new_AGEMA_signal_5901 ) ) ;

    /* cells in depth 8 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1968 ( .a ({new_AGEMA_signal_1309, n1924}), .b ({new_AGEMA_signal_1310, n1923}), .clk ( clk ), .r ( Fresh[451] ), .c ({new_AGEMA_signal_1470, n1936}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1982 ( .a ({new_AGEMA_signal_3080, new_AGEMA_signal_3078}), .b ({new_AGEMA_signal_1311, n1927}), .clk ( clk ), .r ( Fresh[452] ), .c ({new_AGEMA_signal_1471, n1928}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U1994 ( .a ({new_AGEMA_signal_3084, new_AGEMA_signal_3082}), .b ({new_AGEMA_signal_1312, n1929}), .clk ( clk ), .r ( Fresh[453] ), .c ({new_AGEMA_signal_1472, n1931}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2012 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_1314, n1938}), .clk ( clk ), .r ( Fresh[454] ), .c ({new_AGEMA_signal_1473, n1939}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2024 ( .a ({new_AGEMA_signal_1315, n2235}), .b ({new_AGEMA_signal_1137, n1943}), .clk ( clk ), .r ( Fresh[455] ), .c ({new_AGEMA_signal_1474, n1948}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2032 ( .a ({new_AGEMA_signal_1138, n1946}), .b ({new_AGEMA_signal_1316, n1945}), .clk ( clk ), .r ( Fresh[456] ), .c ({new_AGEMA_signal_1475, n1947}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2041 ( .a ({new_AGEMA_signal_3092, new_AGEMA_signal_3088}), .b ({new_AGEMA_signal_1318, n1951}), .clk ( clk ), .r ( Fresh[457] ), .c ({new_AGEMA_signal_1476, n1954}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2049 ( .a ({new_AGEMA_signal_3096, new_AGEMA_signal_3094}), .b ({new_AGEMA_signal_1319, n1952}), .clk ( clk ), .r ( Fresh[458] ), .c ({new_AGEMA_signal_1477, n1953}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2058 ( .a ({new_AGEMA_signal_3100, new_AGEMA_signal_3098}), .b ({new_AGEMA_signal_1320, n2687}), .clk ( clk ), .r ( Fresh[459] ), .c ({new_AGEMA_signal_1478, n2658}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2065 ( .a ({new_AGEMA_signal_3104, new_AGEMA_signal_3102}), .b ({new_AGEMA_signal_1143, n1963}), .clk ( clk ), .r ( Fresh[460] ), .c ({new_AGEMA_signal_1322, n1965}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2078 ( .a ({new_AGEMA_signal_3108, new_AGEMA_signal_3106}), .b ({new_AGEMA_signal_1480, n1968}), .clk ( clk ), .r ( Fresh[461] ), .c ({new_AGEMA_signal_1591, n1970}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2084 ( .a ({new_AGEMA_signal_1325, n2684}), .b ({new_AGEMA_signal_3112, new_AGEMA_signal_3110}), .clk ( clk ), .r ( Fresh[462] ), .c ({new_AGEMA_signal_1481, n1969}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2093 ( .a ({new_AGEMA_signal_1326, n1972}), .b ({new_AGEMA_signal_1149, n1971}), .clk ( clk ), .r ( Fresh[463] ), .c ({new_AGEMA_signal_1482, n1978}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2102 ( .a ({new_AGEMA_signal_1327, n1974}), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3114}), .clk ( clk ), .r ( Fresh[464] ), .c ({new_AGEMA_signal_1483, n1975}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2107 ( .a ({new_AGEMA_signal_3120, new_AGEMA_signal_3118}), .b ({new_AGEMA_signal_1328, n1979}), .clk ( clk ), .r ( Fresh[465] ), .c ({new_AGEMA_signal_1484, n1980}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2114 ( .a ({new_AGEMA_signal_1152, n1985}), .b ({new_AGEMA_signal_3124, new_AGEMA_signal_3122}), .clk ( clk ), .r ( Fresh[466] ), .c ({new_AGEMA_signal_1329, n1986}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2124 ( .a ({new_AGEMA_signal_1330, n1994}), .b ({new_AGEMA_signal_3128, new_AGEMA_signal_3126}), .clk ( clk ), .r ( Fresh[467] ), .c ({new_AGEMA_signal_1486, n1997}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2137 ( .a ({new_AGEMA_signal_3132, new_AGEMA_signal_3130}), .b ({new_AGEMA_signal_1332, n2137}), .clk ( clk ), .r ( Fresh[468] ), .c ({new_AGEMA_signal_1487, n2012}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2145 ( .a ({new_AGEMA_signal_1333, n2006}), .b ({new_AGEMA_signal_1334, n2005}), .clk ( clk ), .r ( Fresh[469] ), .c ({new_AGEMA_signal_1488, n2007}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2161 ( .s ({new_AGEMA_signal_3136, new_AGEMA_signal_3134}), .b ({new_AGEMA_signal_1165, n2020}), .a ({new_AGEMA_signal_3144, new_AGEMA_signal_3140}), .clk ( clk ), .r ( Fresh[470] ), .c ({new_AGEMA_signal_1336, n2021}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2176 ( .a ({new_AGEMA_signal_3148, new_AGEMA_signal_3146}), .b ({new_AGEMA_signal_1338, n2031}), .clk ( clk ), .r ( Fresh[471] ), .c ({new_AGEMA_signal_1490, n2032}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2185 ( .a ({new_AGEMA_signal_3152, new_AGEMA_signal_3150}), .b ({new_AGEMA_signal_1339, n2040}), .clk ( clk ), .r ( Fresh[472] ), .c ({new_AGEMA_signal_1491, n2041}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2189 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_3156, new_AGEMA_signal_3154}), .clk ( clk ), .r ( Fresh[473] ), .c ({new_AGEMA_signal_1492, n2043}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2194 ( .a ({new_AGEMA_signal_3160, new_AGEMA_signal_3158}), .b ({new_AGEMA_signal_1340, n2045}), .clk ( clk ), .r ( Fresh[474] ), .c ({new_AGEMA_signal_1493, n2046}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2204 ( .s ({new_AGEMA_signal_3136, new_AGEMA_signal_3134}), .b ({new_AGEMA_signal_1342, n2056}), .a ({new_AGEMA_signal_3164, new_AGEMA_signal_3162}), .clk ( clk ), .r ( Fresh[475] ), .c ({new_AGEMA_signal_1494, n2058}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2210 ( .a ({new_AGEMA_signal_3168, new_AGEMA_signal_3166}), .b ({new_AGEMA_signal_1343, n2060}), .clk ( clk ), .r ( Fresh[476] ), .c ({new_AGEMA_signal_1495, n2063}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2218 ( .a ({new_AGEMA_signal_1344, n2066}), .b ({new_AGEMA_signal_1345, n2065}), .clk ( clk ), .r ( Fresh[477] ), .c ({new_AGEMA_signal_1496, n2652}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2227 ( .a ({new_AGEMA_signal_3172, new_AGEMA_signal_3170}), .b ({new_AGEMA_signal_1347, n2074}), .clk ( clk ), .r ( Fresh[478] ), .c ({new_AGEMA_signal_1497, n2076}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2236 ( .a ({new_AGEMA_signal_3180, new_AGEMA_signal_3176}), .b ({new_AGEMA_signal_1348, n2082}), .clk ( clk ), .r ( Fresh[479] ), .c ({new_AGEMA_signal_1498, n2105}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2241 ( .a ({new_AGEMA_signal_3184, new_AGEMA_signal_3182}), .b ({new_AGEMA_signal_1349, n2084}), .clk ( clk ), .r ( Fresh[480] ), .c ({new_AGEMA_signal_1499, n2099}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2243 ( .a ({new_AGEMA_signal_1350, n2085}), .b ({new_AGEMA_signal_3188, new_AGEMA_signal_3186}), .clk ( clk ), .r ( Fresh[481] ), .c ({new_AGEMA_signal_1500, n2091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) U2246 ( .a ({new_AGEMA_signal_3192, new_AGEMA_signal_3190}), .b ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .r ( Fresh[482] ), .c ({new_AGEMA_signal_1501, n2090}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2253 ( .a ({new_AGEMA_signal_3196, new_AGEMA_signal_3194}), .b ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .r ( Fresh[483] ), .c ({new_AGEMA_signal_1502, n2093}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2262 ( .a ({new_AGEMA_signal_3200, new_AGEMA_signal_3198}), .b ({new_AGEMA_signal_1356, n2160}), .clk ( clk ), .r ( Fresh[484] ), .c ({new_AGEMA_signal_1503, n2102}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2266 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_3208, new_AGEMA_signal_3204}), .clk ( clk ), .r ( Fresh[485] ), .c ({new_AGEMA_signal_1357, n2106}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2272 ( .a ({new_AGEMA_signal_3212, new_AGEMA_signal_3210}), .b ({new_AGEMA_signal_1504, n2114}), .clk ( clk ), .r ( Fresh[486] ), .c ({new_AGEMA_signal_1606, n2116}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2282 ( .a ({new_AGEMA_signal_1358, n2291}), .b ({new_AGEMA_signal_1192, n2119}), .clk ( clk ), .r ( Fresh[487] ), .c ({new_AGEMA_signal_1505, n2120}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2293 ( .a ({new_AGEMA_signal_1195, n2130}), .b ({new_AGEMA_signal_1196, n2129}), .clk ( clk ), .r ( Fresh[488] ), .c ({new_AGEMA_signal_1359, n2155}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2296 ( .a ({new_AGEMA_signal_3216, new_AGEMA_signal_3214}), .b ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .r ( Fresh[489] ), .c ({new_AGEMA_signal_1506, n2543}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2299 ( .a ({new_AGEMA_signal_1198, n2133}), .b ({new_AGEMA_signal_3220, new_AGEMA_signal_3218}), .clk ( clk ), .r ( Fresh[490] ), .c ({new_AGEMA_signal_1360, n2134}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2303 ( .a ({new_AGEMA_signal_1332, n2137}), .b ({new_AGEMA_signal_1361, n2136}), .clk ( clk ), .r ( Fresh[491] ), .c ({new_AGEMA_signal_1508, n2143}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2308 ( .a ({new_AGEMA_signal_1362, n2139}), .b ({new_AGEMA_signal_3228, new_AGEMA_signal_3224}), .clk ( clk ), .r ( Fresh[492] ), .c ({new_AGEMA_signal_1509, n2140}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2324 ( .a ({new_AGEMA_signal_1366, n2157}), .b ({new_AGEMA_signal_3232, new_AGEMA_signal_3230}), .clk ( clk ), .r ( Fresh[493] ), .c ({new_AGEMA_signal_1510, n2159}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2326 ( .a ({new_AGEMA_signal_1356, n2160}), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3234}), .clk ( clk ), .r ( Fresh[494] ), .c ({new_AGEMA_signal_1511, n2161}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2330 ( .a ({new_AGEMA_signal_3092, new_AGEMA_signal_3088}), .b ({new_AGEMA_signal_1203, n2163}), .clk ( clk ), .r ( Fresh[495] ), .c ({new_AGEMA_signal_1367, n2164}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2345 ( .a ({new_AGEMA_signal_3240, new_AGEMA_signal_3238}), .b ({new_AGEMA_signal_1370, n2177}), .clk ( clk ), .r ( Fresh[496] ), .c ({new_AGEMA_signal_1513, n2179}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2359 ( .a ({new_AGEMA_signal_3248, new_AGEMA_signal_3244}), .b ({new_AGEMA_signal_1373, n2191}), .clk ( clk ), .r ( Fresh[497] ), .c ({new_AGEMA_signal_1514, n2192}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2370 ( .a ({new_AGEMA_signal_1374, n2201}), .b ({new_AGEMA_signal_1515, n2200}), .clk ( clk ), .r ( Fresh[498] ), .c ({new_AGEMA_signal_1613, n2203}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2382 ( .a ({new_AGEMA_signal_1376, n2217}), .b ({new_AGEMA_signal_1210, n2216}), .clk ( clk ), .r ( Fresh[499] ), .c ({new_AGEMA_signal_1517, n2224}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2388 ( .a ({new_AGEMA_signal_1377, n2222}), .b ({new_AGEMA_signal_1378, n2221}), .clk ( clk ), .r ( Fresh[500] ), .c ({new_AGEMA_signal_1518, n2223}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2392 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1213, n2226}), .clk ( clk ), .r ( Fresh[501] ), .c ({new_AGEMA_signal_1379, n2229}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2399 ( .a ({new_AGEMA_signal_3096, new_AGEMA_signal_3094}), .b ({new_AGEMA_signal_1520, n2233}), .clk ( clk ), .r ( Fresh[502] ), .c ({new_AGEMA_signal_1616, n2234}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2410 ( .a ({new_AGEMA_signal_3100, new_AGEMA_signal_3098}), .b ({new_AGEMA_signal_1381, n2244}), .clk ( clk ), .r ( Fresh[503] ), .c ({new_AGEMA_signal_1521, n2246}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2418 ( .a ({new_AGEMA_signal_3252, new_AGEMA_signal_3250}), .b ({new_AGEMA_signal_1383, n2253}), .clk ( clk ), .r ( Fresh[504] ), .c ({new_AGEMA_signal_1522, n2254}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2425 ( .a ({new_AGEMA_signal_3256, new_AGEMA_signal_3254}), .b ({new_AGEMA_signal_1384, n2260}), .clk ( clk ), .r ( Fresh[505] ), .c ({new_AGEMA_signal_1523, n2263}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2434 ( .a ({new_AGEMA_signal_3260, new_AGEMA_signal_3258}), .b ({new_AGEMA_signal_1223, n2265}), .clk ( clk ), .r ( Fresh[506] ), .c ({new_AGEMA_signal_1385, n2267}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2438 ( .a ({new_AGEMA_signal_3096, new_AGEMA_signal_3094}), .b ({new_AGEMA_signal_1224, n2269}), .clk ( clk ), .r ( Fresh[507] ), .c ({new_AGEMA_signal_1386, n2270}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2445 ( .a ({new_AGEMA_signal_3264, new_AGEMA_signal_3262}), .b ({new_AGEMA_signal_1226, n2277}), .clk ( clk ), .r ( Fresh[508] ), .c ({new_AGEMA_signal_1387, n2279}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2450 ( .a ({new_AGEMA_signal_3144, new_AGEMA_signal_3140}), .b ({new_AGEMA_signal_1227, n2282}), .clk ( clk ), .r ( Fresh[509] ), .c ({new_AGEMA_signal_1388, n2283}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2453 ( .a ({new_AGEMA_signal_3184, new_AGEMA_signal_3182}), .b ({new_AGEMA_signal_1389, n2284}), .clk ( clk ), .r ( Fresh[510] ), .c ({new_AGEMA_signal_1528, n2285}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2457 ( .a ({new_AGEMA_signal_3092, new_AGEMA_signal_3088}), .b ({new_AGEMA_signal_1390, n2459}), .clk ( clk ), .r ( Fresh[511] ), .c ({new_AGEMA_signal_1529, n2686}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2460 ( .a ({new_AGEMA_signal_3100, new_AGEMA_signal_3098}), .b ({new_AGEMA_signal_1391, n2288}), .clk ( clk ), .r ( Fresh[512] ), .c ({new_AGEMA_signal_1530, n2289}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2463 ( .a ({new_AGEMA_signal_1392, n2458}), .b ({new_AGEMA_signal_3268, new_AGEMA_signal_3266}), .clk ( clk ), .r ( Fresh[513] ), .c ({new_AGEMA_signal_1531, n2297}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2465 ( .a ({new_AGEMA_signal_3272, new_AGEMA_signal_3270}), .b ({new_AGEMA_signal_1358, n2291}), .clk ( clk ), .r ( Fresh[514] ), .c ({new_AGEMA_signal_1532, n2292}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2473 ( .a ({new_AGEMA_signal_3276, new_AGEMA_signal_3274}), .b ({new_AGEMA_signal_1394, n2300}), .clk ( clk ), .r ( Fresh[515] ), .c ({new_AGEMA_signal_1533, n2301}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2483 ( .a ({new_AGEMA_signal_3280, new_AGEMA_signal_3278}), .b ({new_AGEMA_signal_1396, n2314}), .clk ( clk ), .r ( Fresh[516] ), .c ({new_AGEMA_signal_1534, n2321}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2487 ( .a ({new_AGEMA_signal_1097, n2319}), .b ({new_AGEMA_signal_3284, new_AGEMA_signal_3282}), .clk ( clk ), .r ( Fresh[517] ), .c ({new_AGEMA_signal_1233, n2320}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2493 ( .a ({new_AGEMA_signal_1234, n2326}), .b ({new_AGEMA_signal_3288, new_AGEMA_signal_3286}), .clk ( clk ), .r ( Fresh[518] ), .c ({new_AGEMA_signal_1397, n2334}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2497 ( .a ({new_AGEMA_signal_1398, n2329}), .b ({new_AGEMA_signal_3144, new_AGEMA_signal_3140}), .clk ( clk ), .r ( Fresh[519] ), .c ({new_AGEMA_signal_1535, n2332}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2498 ( .a ({new_AGEMA_signal_3292, new_AGEMA_signal_3290}), .b ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .r ( Fresh[520] ), .c ({new_AGEMA_signal_1536, n2331}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2502 ( .a ({new_AGEMA_signal_3296, new_AGEMA_signal_3294}), .b ({new_AGEMA_signal_1537, n2335}), .clk ( clk ), .r ( Fresh[521] ), .c ({new_AGEMA_signal_1626, n2336}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2508 ( .a ({new_AGEMA_signal_1399, n2341}), .b ({new_AGEMA_signal_1238, n2340}), .clk ( clk ), .r ( Fresh[522] ), .c ({new_AGEMA_signal_1538, n2342}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2519 ( .a ({new_AGEMA_signal_1242, n2352}), .b ({new_AGEMA_signal_3300, new_AGEMA_signal_3298}), .clk ( clk ), .r ( Fresh[523] ), .c ({new_AGEMA_signal_1400, n2367}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2523 ( .a ({new_AGEMA_signal_1401, n2354}), .b ({new_AGEMA_signal_3304, new_AGEMA_signal_3302}), .clk ( clk ), .r ( Fresh[524] ), .c ({new_AGEMA_signal_1539, n2358}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2547 ( .a ({new_AGEMA_signal_1247, n2385}), .b ({new_AGEMA_signal_1248, n2384}), .clk ( clk ), .r ( Fresh[525] ), .c ({new_AGEMA_signal_1406, n2387}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2555 ( .a ({new_AGEMA_signal_1250, n2391}), .b ({new_AGEMA_signal_1408, n2390}), .clk ( clk ), .r ( Fresh[526] ), .c ({new_AGEMA_signal_1542, n2392}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2566 ( .a ({new_AGEMA_signal_1252, n2403}), .b ({new_AGEMA_signal_3308, new_AGEMA_signal_3306}), .clk ( clk ), .r ( Fresh[527] ), .c ({new_AGEMA_signal_1410, n2404}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2570 ( .a ({new_AGEMA_signal_3168, new_AGEMA_signal_3166}), .b ({new_AGEMA_signal_1411, n2408}), .clk ( clk ), .r ( Fresh[528] ), .c ({new_AGEMA_signal_1544, n2409}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2575 ( .a ({new_AGEMA_signal_1412, n2574}), .b ({new_AGEMA_signal_1253, n2413}), .clk ( clk ), .r ( Fresh[529] ), .c ({new_AGEMA_signal_1545, n2414}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2578 ( .a ({new_AGEMA_signal_3312, new_AGEMA_signal_3310}), .b ({new_AGEMA_signal_1254, n2416}), .clk ( clk ), .r ( Fresh[530] ), .c ({new_AGEMA_signal_1413, n2418}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2589 ( .a ({new_AGEMA_signal_1415, n2689}), .b ({new_AGEMA_signal_3316, new_AGEMA_signal_3314}), .clk ( clk ), .r ( Fresh[531] ), .c ({new_AGEMA_signal_1547, n2432}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2592 ( .a ({new_AGEMA_signal_3328, new_AGEMA_signal_3322}), .b ({new_AGEMA_signal_1257, n2434}), .clk ( clk ), .r ( Fresh[532] ), .c ({new_AGEMA_signal_1416, n2435}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2601 ( .a ({new_AGEMA_signal_1418, n2445}), .b ({new_AGEMA_signal_1419, n2444}), .clk ( clk ), .r ( Fresh[533] ), .c ({new_AGEMA_signal_1548, n2449}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2603 ( .a ({new_AGEMA_signal_3280, new_AGEMA_signal_3278}), .b ({new_AGEMA_signal_1420, n2447}), .clk ( clk ), .r ( Fresh[534] ), .c ({new_AGEMA_signal_1549, n2448}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2609 ( .a ({new_AGEMA_signal_1421, n2454}), .b ({new_AGEMA_signal_3332, new_AGEMA_signal_3330}), .clk ( clk ), .r ( Fresh[535] ), .c ({new_AGEMA_signal_1550, n2455}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2612 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_1392, n2458}), .clk ( clk ), .r ( Fresh[536] ), .c ({new_AGEMA_signal_1551, n2460}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2618 ( .a ({new_AGEMA_signal_3272, new_AGEMA_signal_3270}), .b ({new_AGEMA_signal_1260, n2465}), .clk ( clk ), .r ( Fresh[537] ), .c ({new_AGEMA_signal_1422, n2466}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2629 ( .a ({new_AGEMA_signal_1262, n2476}), .b ({new_AGEMA_signal_3336, new_AGEMA_signal_3334}), .clk ( clk ), .r ( Fresh[538] ), .c ({new_AGEMA_signal_1423, n2477}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2634 ( .a ({new_AGEMA_signal_3164, new_AGEMA_signal_3162}), .b ({new_AGEMA_signal_1424, n2481}), .clk ( clk ), .r ( Fresh[539] ), .c ({new_AGEMA_signal_1554, n2482}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2640 ( .a ({new_AGEMA_signal_3340, new_AGEMA_signal_3338}), .b ({new_AGEMA_signal_1265, n2486}), .clk ( clk ), .r ( Fresh[540] ), .c ({new_AGEMA_signal_1425, n2490}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2648 ( .a ({new_AGEMA_signal_1268, n2495}), .b ({new_AGEMA_signal_1426, n2494}), .clk ( clk ), .r ( Fresh[541] ), .c ({new_AGEMA_signal_1556, n2496}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2654 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1557, n2503}), .clk ( clk ), .r ( Fresh[542] ), .c ({new_AGEMA_signal_1643, n2507}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2664 ( .a ({new_AGEMA_signal_1428, n2518}), .b ({new_AGEMA_signal_1558, n2517}), .clk ( clk ), .r ( Fresh[543] ), .c ({new_AGEMA_signal_1644, n2525}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2669 ( .a ({new_AGEMA_signal_1429, n2523}), .b ({new_AGEMA_signal_1430, n2522}), .clk ( clk ), .r ( Fresh[544] ), .c ({new_AGEMA_signal_1559, n2524}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2676 ( .a ({new_AGEMA_signal_1431, n2532}), .b ({new_AGEMA_signal_3348, new_AGEMA_signal_3344}), .clk ( clk ), .r ( Fresh[545] ), .c ({new_AGEMA_signal_1560, n2537}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2678 ( .a ({new_AGEMA_signal_3168, new_AGEMA_signal_3166}), .b ({new_AGEMA_signal_1432, n2534}), .clk ( clk ), .r ( Fresh[546] ), .c ({new_AGEMA_signal_1561, n2536}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2684 ( .a ({new_AGEMA_signal_3352, new_AGEMA_signal_3350}), .b ({new_AGEMA_signal_1272, n2546}), .clk ( clk ), .r ( Fresh[547] ), .c ({new_AGEMA_signal_1434, n2547}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2693 ( .a ({new_AGEMA_signal_3356, new_AGEMA_signal_3354}), .b ({new_AGEMA_signal_1437, n2556}), .clk ( clk ), .r ( Fresh[548] ), .c ({new_AGEMA_signal_1562, n2557}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2699 ( .a ({new_AGEMA_signal_1439, n2715}), .b ({new_AGEMA_signal_3360, new_AGEMA_signal_3358}), .clk ( clk ), .r ( Fresh[549] ), .c ({new_AGEMA_signal_1563, n2565}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2704 ( .a ({new_AGEMA_signal_1412, n2574}), .b ({new_AGEMA_signal_1440, n2573}), .clk ( clk ), .r ( Fresh[550] ), .c ({new_AGEMA_signal_1564, n2591}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2709 ( .a ({new_AGEMA_signal_1442, n2579}), .b ({new_AGEMA_signal_1277, n2578}), .clk ( clk ), .r ( Fresh[551] ), .c ({new_AGEMA_signal_1565, n2580}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2727 ( .a ({new_AGEMA_signal_1118, n2601}), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3364}), .clk ( clk ), .r ( Fresh[552] ), .c ({new_AGEMA_signal_1282, n2602}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2738 ( .a ({new_AGEMA_signal_1448, n2618}), .b ({new_AGEMA_signal_3372, new_AGEMA_signal_3370}), .clk ( clk ), .r ( Fresh[553] ), .c ({new_AGEMA_signal_1567, n2619}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2744 ( .a ({new_AGEMA_signal_3188, new_AGEMA_signal_3186}), .b ({new_AGEMA_signal_1449, n2626}), .clk ( clk ), .r ( Fresh[554] ), .c ({new_AGEMA_signal_1568, n2628}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2753 ( .a ({new_AGEMA_signal_1450, n2644}), .b ({new_AGEMA_signal_3216, new_AGEMA_signal_3214}), .clk ( clk ), .r ( Fresh[555] ), .c ({new_AGEMA_signal_1569, n2649}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2755 ( .a ({new_AGEMA_signal_3376, new_AGEMA_signal_3374}), .b ({new_AGEMA_signal_1288, n2646}), .clk ( clk ), .r ( Fresh[556] ), .c ({new_AGEMA_signal_1451, n2648}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2765 ( .a ({new_AGEMA_signal_3100, new_AGEMA_signal_3098}), .b ({new_AGEMA_signal_1453, n2663}), .clk ( clk ), .r ( Fresh[557] ), .c ({new_AGEMA_signal_1570, n2664}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2771 ( .a ({new_AGEMA_signal_1290, n2675}), .b ({new_AGEMA_signal_3380, new_AGEMA_signal_3378}), .clk ( clk ), .r ( Fresh[558] ), .c ({new_AGEMA_signal_1571, n2681}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2773 ( .a ({new_AGEMA_signal_3232, new_AGEMA_signal_3230}), .b ({new_AGEMA_signal_1291, n2678}), .clk ( clk ), .r ( Fresh[559] ), .c ({new_AGEMA_signal_1454, n2680}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2776 ( .a ({new_AGEMA_signal_1325, n2684}), .b ({new_AGEMA_signal_3384, new_AGEMA_signal_3382}), .clk ( clk ), .r ( Fresh[560] ), .c ({new_AGEMA_signal_1572, n2685}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2778 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_3352, new_AGEMA_signal_3350}), .clk ( clk ), .r ( Fresh[561] ), .c ({new_AGEMA_signal_1573, n2698}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2779 ( .a ({new_AGEMA_signal_1415, n2689}), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3354}), .clk ( clk ), .r ( Fresh[562] ), .c ({new_AGEMA_signal_1574, n2692}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2793 ( .a ({new_AGEMA_signal_1439, n2715}), .b ({new_AGEMA_signal_3388, new_AGEMA_signal_3386}), .clk ( clk ), .r ( Fresh[563] ), .c ({new_AGEMA_signal_1575, n2716}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2800 ( .a ({new_AGEMA_signal_1296, n2727}), .b ({new_AGEMA_signal_3392, new_AGEMA_signal_3390}), .clk ( clk ), .r ( Fresh[564] ), .c ({new_AGEMA_signal_1457, n2728}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2804 ( .a ({new_AGEMA_signal_3396, new_AGEMA_signal_3394}), .b ({new_AGEMA_signal_1458, n2733}), .clk ( clk ), .r ( Fresh[565] ), .c ({new_AGEMA_signal_1577, n2735}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2808 ( .a ({new_AGEMA_signal_3124, new_AGEMA_signal_3122}), .b ({new_AGEMA_signal_1459, n2740}), .clk ( clk ), .r ( Fresh[566] ), .c ({new_AGEMA_signal_1578, n2743}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2813 ( .a ({new_AGEMA_signal_3404, new_AGEMA_signal_3400}), .b ({new_AGEMA_signal_1299, n2749}), .clk ( clk ), .r ( Fresh[567] ), .c ({new_AGEMA_signal_1460, n2751}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2817 ( .a ({new_AGEMA_signal_1461, n2757}), .b ({new_AGEMA_signal_1300, n2756}), .clk ( clk ), .r ( Fresh[568] ), .c ({new_AGEMA_signal_1579, n2758}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2820 ( .a ({new_AGEMA_signal_3408, new_AGEMA_signal_3406}), .b ({new_AGEMA_signal_1462, n2762}), .clk ( clk ), .r ( Fresh[569] ), .c ({new_AGEMA_signal_1580, n2764}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2827 ( .a ({new_AGEMA_signal_1464, n2776}), .b ({new_AGEMA_signal_1465, n2775}), .clk ( clk ), .r ( Fresh[570] ), .c ({new_AGEMA_signal_1581, n2800}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2831 ( .a ({new_AGEMA_signal_3412, new_AGEMA_signal_3410}), .b ({new_AGEMA_signal_1302, n2783}), .clk ( clk ), .r ( Fresh[571] ), .c ({new_AGEMA_signal_1466, n2788}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2837 ( .a ({new_AGEMA_signal_3420, new_AGEMA_signal_3416}), .b ({new_AGEMA_signal_1467, n2795}), .clk ( clk ), .r ( Fresh[572] ), .c ({new_AGEMA_signal_1583, n2797}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2846 ( .a ({new_AGEMA_signal_1468, n2814}), .b ({new_AGEMA_signal_3136, new_AGEMA_signal_3134}), .clk ( clk ), .r ( Fresh[573] ), .c ({new_AGEMA_signal_1584, n2822}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2849 ( .a ({new_AGEMA_signal_3424, new_AGEMA_signal_3422}), .b ({new_AGEMA_signal_1307, n2819}), .clk ( clk ), .r ( Fresh[574] ), .c ({new_AGEMA_signal_1469, n2821}) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C ( clk ), .D ( new_AGEMA_signal_3427 ), .Q ( new_AGEMA_signal_3428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C ( clk ), .D ( new_AGEMA_signal_3431 ), .Q ( new_AGEMA_signal_3432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C ( clk ), .D ( new_AGEMA_signal_3435 ), .Q ( new_AGEMA_signal_3436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C ( clk ), .D ( new_AGEMA_signal_3439 ), .Q ( new_AGEMA_signal_3440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C ( clk ), .D ( new_AGEMA_signal_3441 ), .Q ( new_AGEMA_signal_3442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C ( clk ), .D ( new_AGEMA_signal_3443 ), .Q ( new_AGEMA_signal_3444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C ( clk ), .D ( new_AGEMA_signal_3445 ), .Q ( new_AGEMA_signal_3446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C ( clk ), .D ( new_AGEMA_signal_3447 ), .Q ( new_AGEMA_signal_3448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C ( clk ), .D ( new_AGEMA_signal_3451 ), .Q ( new_AGEMA_signal_3452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C ( clk ), .D ( new_AGEMA_signal_3455 ), .Q ( new_AGEMA_signal_3456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C ( clk ), .D ( new_AGEMA_signal_3457 ), .Q ( new_AGEMA_signal_3458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C ( clk ), .D ( new_AGEMA_signal_3459 ), .Q ( new_AGEMA_signal_3460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C ( clk ), .D ( new_AGEMA_signal_3463 ), .Q ( new_AGEMA_signal_3464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C ( clk ), .D ( new_AGEMA_signal_3467 ), .Q ( new_AGEMA_signal_3468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C ( clk ), .D ( new_AGEMA_signal_3469 ), .Q ( new_AGEMA_signal_3470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C ( clk ), .D ( new_AGEMA_signal_3471 ), .Q ( new_AGEMA_signal_3472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C ( clk ), .D ( new_AGEMA_signal_3475 ), .Q ( new_AGEMA_signal_3476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C ( clk ), .D ( new_AGEMA_signal_3479 ), .Q ( new_AGEMA_signal_3480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C ( clk ), .D ( new_AGEMA_signal_3483 ), .Q ( new_AGEMA_signal_3484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C ( clk ), .D ( new_AGEMA_signal_3487 ), .Q ( new_AGEMA_signal_3488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C ( clk ), .D ( new_AGEMA_signal_3489 ), .Q ( new_AGEMA_signal_3490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C ( clk ), .D ( new_AGEMA_signal_3491 ), .Q ( new_AGEMA_signal_3492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C ( clk ), .D ( new_AGEMA_signal_3493 ), .Q ( new_AGEMA_signal_3494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C ( clk ), .D ( new_AGEMA_signal_3495 ), .Q ( new_AGEMA_signal_3496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C ( clk ), .D ( new_AGEMA_signal_3497 ), .Q ( new_AGEMA_signal_3498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C ( clk ), .D ( new_AGEMA_signal_3499 ), .Q ( new_AGEMA_signal_3500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C ( clk ), .D ( new_AGEMA_signal_3501 ), .Q ( new_AGEMA_signal_3502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C ( clk ), .D ( new_AGEMA_signal_3503 ), .Q ( new_AGEMA_signal_3504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C ( clk ), .D ( new_AGEMA_signal_3507 ), .Q ( new_AGEMA_signal_3508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C ( clk ), .D ( new_AGEMA_signal_3511 ), .Q ( new_AGEMA_signal_3512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C ( clk ), .D ( new_AGEMA_signal_3515 ), .Q ( new_AGEMA_signal_3516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C ( clk ), .D ( new_AGEMA_signal_3519 ), .Q ( new_AGEMA_signal_3520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C ( clk ), .D ( new_AGEMA_signal_3523 ), .Q ( new_AGEMA_signal_3524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C ( clk ), .D ( new_AGEMA_signal_3527 ), .Q ( new_AGEMA_signal_3528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C ( clk ), .D ( new_AGEMA_signal_3529 ), .Q ( new_AGEMA_signal_3530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C ( clk ), .D ( new_AGEMA_signal_3531 ), .Q ( new_AGEMA_signal_3532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C ( clk ), .D ( new_AGEMA_signal_3533 ), .Q ( new_AGEMA_signal_3534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C ( clk ), .D ( new_AGEMA_signal_3535 ), .Q ( new_AGEMA_signal_3536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C ( clk ), .D ( new_AGEMA_signal_3537 ), .Q ( new_AGEMA_signal_3538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C ( clk ), .D ( new_AGEMA_signal_3539 ), .Q ( new_AGEMA_signal_3540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C ( clk ), .D ( new_AGEMA_signal_3543 ), .Q ( new_AGEMA_signal_3544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C ( clk ), .D ( new_AGEMA_signal_3547 ), .Q ( new_AGEMA_signal_3548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C ( clk ), .D ( new_AGEMA_signal_3549 ), .Q ( new_AGEMA_signal_3550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C ( clk ), .D ( new_AGEMA_signal_3551 ), .Q ( new_AGEMA_signal_3552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C ( clk ), .D ( new_AGEMA_signal_3555 ), .Q ( new_AGEMA_signal_3556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C ( clk ), .D ( new_AGEMA_signal_3559 ), .Q ( new_AGEMA_signal_3560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C ( clk ), .D ( new_AGEMA_signal_3565 ), .Q ( new_AGEMA_signal_3566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C ( clk ), .D ( new_AGEMA_signal_3571 ), .Q ( new_AGEMA_signal_3572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C ( clk ), .D ( new_AGEMA_signal_3575 ), .Q ( new_AGEMA_signal_3576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C ( clk ), .D ( new_AGEMA_signal_3579 ), .Q ( new_AGEMA_signal_3580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C ( clk ), .D ( new_AGEMA_signal_3583 ), .Q ( new_AGEMA_signal_3584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C ( clk ), .D ( new_AGEMA_signal_3587 ), .Q ( new_AGEMA_signal_3588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C ( clk ), .D ( new_AGEMA_signal_3589 ), .Q ( new_AGEMA_signal_3590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C ( clk ), .D ( new_AGEMA_signal_3591 ), .Q ( new_AGEMA_signal_3592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C ( clk ), .D ( new_AGEMA_signal_3593 ), .Q ( new_AGEMA_signal_3594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C ( clk ), .D ( new_AGEMA_signal_3595 ), .Q ( new_AGEMA_signal_3596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C ( clk ), .D ( new_AGEMA_signal_3597 ), .Q ( new_AGEMA_signal_3598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C ( clk ), .D ( new_AGEMA_signal_3599 ), .Q ( new_AGEMA_signal_3600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C ( clk ), .D ( new_AGEMA_signal_3601 ), .Q ( new_AGEMA_signal_3602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C ( clk ), .D ( new_AGEMA_signal_3603 ), .Q ( new_AGEMA_signal_3604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C ( clk ), .D ( new_AGEMA_signal_3607 ), .Q ( new_AGEMA_signal_3608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C ( clk ), .D ( new_AGEMA_signal_3611 ), .Q ( new_AGEMA_signal_3612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C ( clk ), .D ( new_AGEMA_signal_3617 ), .Q ( new_AGEMA_signal_3618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C ( clk ), .D ( new_AGEMA_signal_3623 ), .Q ( new_AGEMA_signal_3624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C ( clk ), .D ( new_AGEMA_signal_3627 ), .Q ( new_AGEMA_signal_3628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C ( clk ), .D ( new_AGEMA_signal_3631 ), .Q ( new_AGEMA_signal_3632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C ( clk ), .D ( new_AGEMA_signal_3633 ), .Q ( new_AGEMA_signal_3634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C ( clk ), .D ( new_AGEMA_signal_3635 ), .Q ( new_AGEMA_signal_3636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C ( clk ), .D ( new_AGEMA_signal_3637 ), .Q ( new_AGEMA_signal_3638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C ( clk ), .D ( new_AGEMA_signal_3639 ), .Q ( new_AGEMA_signal_3640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C ( clk ), .D ( new_AGEMA_signal_3641 ), .Q ( new_AGEMA_signal_3642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C ( clk ), .D ( new_AGEMA_signal_3643 ), .Q ( new_AGEMA_signal_3644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C ( clk ), .D ( new_AGEMA_signal_3647 ), .Q ( new_AGEMA_signal_3648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C ( clk ), .D ( new_AGEMA_signal_3651 ), .Q ( new_AGEMA_signal_3652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C ( clk ), .D ( new_AGEMA_signal_3653 ), .Q ( new_AGEMA_signal_3654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C ( clk ), .D ( new_AGEMA_signal_3655 ), .Q ( new_AGEMA_signal_3656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C ( clk ), .D ( new_AGEMA_signal_3657 ), .Q ( new_AGEMA_signal_3658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C ( clk ), .D ( new_AGEMA_signal_3659 ), .Q ( new_AGEMA_signal_3660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C ( clk ), .D ( new_AGEMA_signal_3663 ), .Q ( new_AGEMA_signal_3664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C ( clk ), .D ( new_AGEMA_signal_3667 ), .Q ( new_AGEMA_signal_3668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C ( clk ), .D ( new_AGEMA_signal_3671 ), .Q ( new_AGEMA_signal_3672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C ( clk ), .D ( new_AGEMA_signal_3675 ), .Q ( new_AGEMA_signal_3676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C ( clk ), .D ( new_AGEMA_signal_3679 ), .Q ( new_AGEMA_signal_3680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C ( clk ), .D ( new_AGEMA_signal_3683 ), .Q ( new_AGEMA_signal_3684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C ( clk ), .D ( new_AGEMA_signal_3687 ), .Q ( new_AGEMA_signal_3688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C ( clk ), .D ( new_AGEMA_signal_3691 ), .Q ( new_AGEMA_signal_3692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C ( clk ), .D ( new_AGEMA_signal_3695 ), .Q ( new_AGEMA_signal_3696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C ( clk ), .D ( new_AGEMA_signal_3699 ), .Q ( new_AGEMA_signal_3700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C ( clk ), .D ( new_AGEMA_signal_3701 ), .Q ( new_AGEMA_signal_3702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C ( clk ), .D ( new_AGEMA_signal_3703 ), .Q ( new_AGEMA_signal_3704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C ( clk ), .D ( new_AGEMA_signal_3705 ), .Q ( new_AGEMA_signal_3706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C ( clk ), .D ( new_AGEMA_signal_3707 ), .Q ( new_AGEMA_signal_3708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C ( clk ), .D ( new_AGEMA_signal_3709 ), .Q ( new_AGEMA_signal_3710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C ( clk ), .D ( new_AGEMA_signal_3711 ), .Q ( new_AGEMA_signal_3712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C ( clk ), .D ( new_AGEMA_signal_3713 ), .Q ( new_AGEMA_signal_3714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C ( clk ), .D ( new_AGEMA_signal_3715 ), .Q ( new_AGEMA_signal_3716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C ( clk ), .D ( new_AGEMA_signal_3719 ), .Q ( new_AGEMA_signal_3720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C ( clk ), .D ( new_AGEMA_signal_3723 ), .Q ( new_AGEMA_signal_3724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C ( clk ), .D ( new_AGEMA_signal_3727 ), .Q ( new_AGEMA_signal_3728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C ( clk ), .D ( new_AGEMA_signal_3731 ), .Q ( new_AGEMA_signal_3732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C ( clk ), .D ( new_AGEMA_signal_3733 ), .Q ( new_AGEMA_signal_3734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C ( clk ), .D ( new_AGEMA_signal_3735 ), .Q ( new_AGEMA_signal_3736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C ( clk ), .D ( new_AGEMA_signal_3737 ), .Q ( new_AGEMA_signal_3738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C ( clk ), .D ( new_AGEMA_signal_3739 ), .Q ( new_AGEMA_signal_3740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C ( clk ), .D ( new_AGEMA_signal_3741 ), .Q ( new_AGEMA_signal_3742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C ( clk ), .D ( new_AGEMA_signal_3743 ), .Q ( new_AGEMA_signal_3744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C ( clk ), .D ( new_AGEMA_signal_3745 ), .Q ( new_AGEMA_signal_3746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C ( clk ), .D ( new_AGEMA_signal_3747 ), .Q ( new_AGEMA_signal_3748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C ( clk ), .D ( new_AGEMA_signal_3749 ), .Q ( new_AGEMA_signal_3750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C ( clk ), .D ( new_AGEMA_signal_3751 ), .Q ( new_AGEMA_signal_3752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C ( clk ), .D ( new_AGEMA_signal_3753 ), .Q ( new_AGEMA_signal_3754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C ( clk ), .D ( new_AGEMA_signal_3755 ), .Q ( new_AGEMA_signal_3756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C ( clk ), .D ( new_AGEMA_signal_3757 ), .Q ( new_AGEMA_signal_3758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C ( clk ), .D ( new_AGEMA_signal_3759 ), .Q ( new_AGEMA_signal_3760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C ( clk ), .D ( new_AGEMA_signal_3761 ), .Q ( new_AGEMA_signal_3762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C ( clk ), .D ( new_AGEMA_signal_3763 ), .Q ( new_AGEMA_signal_3764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C ( clk ), .D ( new_AGEMA_signal_3765 ), .Q ( new_AGEMA_signal_3766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C ( clk ), .D ( new_AGEMA_signal_3767 ), .Q ( new_AGEMA_signal_3768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C ( clk ), .D ( new_AGEMA_signal_3771 ), .Q ( new_AGEMA_signal_3772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C ( clk ), .D ( new_AGEMA_signal_3775 ), .Q ( new_AGEMA_signal_3776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C ( clk ), .D ( new_AGEMA_signal_3777 ), .Q ( new_AGEMA_signal_3778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C ( clk ), .D ( new_AGEMA_signal_3779 ), .Q ( new_AGEMA_signal_3780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C ( clk ), .D ( new_AGEMA_signal_3781 ), .Q ( new_AGEMA_signal_3782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C ( clk ), .D ( new_AGEMA_signal_3783 ), .Q ( new_AGEMA_signal_3784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C ( clk ), .D ( new_AGEMA_signal_3785 ), .Q ( new_AGEMA_signal_3786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C ( clk ), .D ( new_AGEMA_signal_3787 ), .Q ( new_AGEMA_signal_3788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C ( clk ), .D ( new_AGEMA_signal_3789 ), .Q ( new_AGEMA_signal_3790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C ( clk ), .D ( new_AGEMA_signal_3791 ), .Q ( new_AGEMA_signal_3792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C ( clk ), .D ( new_AGEMA_signal_3793 ), .Q ( new_AGEMA_signal_3794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C ( clk ), .D ( new_AGEMA_signal_3795 ), .Q ( new_AGEMA_signal_3796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C ( clk ), .D ( new_AGEMA_signal_3799 ), .Q ( new_AGEMA_signal_3800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C ( clk ), .D ( new_AGEMA_signal_3803 ), .Q ( new_AGEMA_signal_3804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C ( clk ), .D ( new_AGEMA_signal_3807 ), .Q ( new_AGEMA_signal_3808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C ( clk ), .D ( new_AGEMA_signal_3811 ), .Q ( new_AGEMA_signal_3812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C ( clk ), .D ( new_AGEMA_signal_3815 ), .Q ( new_AGEMA_signal_3816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C ( clk ), .D ( new_AGEMA_signal_3819 ), .Q ( new_AGEMA_signal_3820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C ( clk ), .D ( new_AGEMA_signal_3823 ), .Q ( new_AGEMA_signal_3824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C ( clk ), .D ( new_AGEMA_signal_3827 ), .Q ( new_AGEMA_signal_3828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C ( clk ), .D ( new_AGEMA_signal_3829 ), .Q ( new_AGEMA_signal_3830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C ( clk ), .D ( new_AGEMA_signal_3833 ), .Q ( new_AGEMA_signal_3834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C ( clk ), .D ( new_AGEMA_signal_3837 ), .Q ( new_AGEMA_signal_3838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C ( clk ), .D ( new_AGEMA_signal_3841 ), .Q ( new_AGEMA_signal_3842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C ( clk ), .D ( new_AGEMA_signal_3849 ), .Q ( new_AGEMA_signal_3850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C ( clk ), .D ( new_AGEMA_signal_3857 ), .Q ( new_AGEMA_signal_3858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C ( clk ), .D ( new_AGEMA_signal_3869 ), .Q ( new_AGEMA_signal_3870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C ( clk ), .D ( new_AGEMA_signal_3877 ), .Q ( new_AGEMA_signal_3878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C ( clk ), .D ( new_AGEMA_signal_3883 ), .Q ( new_AGEMA_signal_3884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C ( clk ), .D ( new_AGEMA_signal_3889 ), .Q ( new_AGEMA_signal_3890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C ( clk ), .D ( new_AGEMA_signal_3893 ), .Q ( new_AGEMA_signal_3894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C ( clk ), .D ( new_AGEMA_signal_3897 ), .Q ( new_AGEMA_signal_3898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C ( clk ), .D ( new_AGEMA_signal_3903 ), .Q ( new_AGEMA_signal_3904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C ( clk ), .D ( new_AGEMA_signal_3909 ), .Q ( new_AGEMA_signal_3910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C ( clk ), .D ( new_AGEMA_signal_3919 ), .Q ( new_AGEMA_signal_3920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C ( clk ), .D ( new_AGEMA_signal_3925 ), .Q ( new_AGEMA_signal_3926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C ( clk ), .D ( new_AGEMA_signal_3931 ), .Q ( new_AGEMA_signal_3932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C ( clk ), .D ( new_AGEMA_signal_3937 ), .Q ( new_AGEMA_signal_3938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C ( clk ), .D ( new_AGEMA_signal_3945 ), .Q ( new_AGEMA_signal_3946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C ( clk ), .D ( new_AGEMA_signal_3949 ), .Q ( new_AGEMA_signal_3950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C ( clk ), .D ( new_AGEMA_signal_3955 ), .Q ( new_AGEMA_signal_3956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C ( clk ), .D ( new_AGEMA_signal_3961 ), .Q ( new_AGEMA_signal_3962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C ( clk ), .D ( new_AGEMA_signal_3967 ), .Q ( new_AGEMA_signal_3968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C ( clk ), .D ( new_AGEMA_signal_3973 ), .Q ( new_AGEMA_signal_3974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C ( clk ), .D ( new_AGEMA_signal_3983 ), .Q ( new_AGEMA_signal_3984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C ( clk ), .D ( new_AGEMA_signal_3989 ), .Q ( new_AGEMA_signal_3990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C ( clk ), .D ( new_AGEMA_signal_3997 ), .Q ( new_AGEMA_signal_3998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C ( clk ), .D ( new_AGEMA_signal_4001 ), .Q ( new_AGEMA_signal_4002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C ( clk ), .D ( new_AGEMA_signal_4005 ), .Q ( new_AGEMA_signal_4006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C ( clk ), .D ( new_AGEMA_signal_4009 ), .Q ( new_AGEMA_signal_4010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C ( clk ), .D ( new_AGEMA_signal_4021 ), .Q ( new_AGEMA_signal_4022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C ( clk ), .D ( new_AGEMA_signal_4029 ), .Q ( new_AGEMA_signal_4030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C ( clk ), .D ( new_AGEMA_signal_4035 ), .Q ( new_AGEMA_signal_4036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C ( clk ), .D ( new_AGEMA_signal_4041 ), .Q ( new_AGEMA_signal_4042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C ( clk ), .D ( new_AGEMA_signal_4045 ), .Q ( new_AGEMA_signal_4046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C ( clk ), .D ( new_AGEMA_signal_4049 ), .Q ( new_AGEMA_signal_4050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C ( clk ), .D ( new_AGEMA_signal_4053 ), .Q ( new_AGEMA_signal_4054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C ( clk ), .D ( new_AGEMA_signal_4057 ), .Q ( new_AGEMA_signal_4058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C ( clk ), .D ( new_AGEMA_signal_4069 ), .Q ( new_AGEMA_signal_4070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C ( clk ), .D ( new_AGEMA_signal_4073 ), .Q ( new_AGEMA_signal_4074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C ( clk ), .D ( new_AGEMA_signal_4077 ), .Q ( new_AGEMA_signal_4078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C ( clk ), .D ( new_AGEMA_signal_4081 ), .Q ( new_AGEMA_signal_4082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C ( clk ), .D ( new_AGEMA_signal_4091 ), .Q ( new_AGEMA_signal_4092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C ( clk ), .D ( new_AGEMA_signal_4097 ), .Q ( new_AGEMA_signal_4098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C ( clk ), .D ( new_AGEMA_signal_4101 ), .Q ( new_AGEMA_signal_4102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C ( clk ), .D ( new_AGEMA_signal_4105 ), .Q ( new_AGEMA_signal_4106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C ( clk ), .D ( new_AGEMA_signal_4113 ), .Q ( new_AGEMA_signal_4114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C ( clk ), .D ( new_AGEMA_signal_4117 ), .Q ( new_AGEMA_signal_4118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C ( clk ), .D ( new_AGEMA_signal_4121 ), .Q ( new_AGEMA_signal_4122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C ( clk ), .D ( new_AGEMA_signal_4125 ), .Q ( new_AGEMA_signal_4126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C ( clk ), .D ( new_AGEMA_signal_4129 ), .Q ( new_AGEMA_signal_4130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C ( clk ), .D ( new_AGEMA_signal_4133 ), .Q ( new_AGEMA_signal_4134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C ( clk ), .D ( new_AGEMA_signal_4141 ), .Q ( new_AGEMA_signal_4142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C ( clk ), .D ( new_AGEMA_signal_4145 ), .Q ( new_AGEMA_signal_4146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C ( clk ), .D ( new_AGEMA_signal_4155 ), .Q ( new_AGEMA_signal_4156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C ( clk ), .D ( new_AGEMA_signal_4161 ), .Q ( new_AGEMA_signal_4162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C ( clk ), .D ( new_AGEMA_signal_4167 ), .Q ( new_AGEMA_signal_4168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C ( clk ), .D ( new_AGEMA_signal_4173 ), .Q ( new_AGEMA_signal_4174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C ( clk ), .D ( new_AGEMA_signal_4177 ), .Q ( new_AGEMA_signal_4178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C ( clk ), .D ( new_AGEMA_signal_4181 ), .Q ( new_AGEMA_signal_4182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C ( clk ), .D ( new_AGEMA_signal_4193 ), .Q ( new_AGEMA_signal_4194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C ( clk ), .D ( new_AGEMA_signal_4201 ), .Q ( new_AGEMA_signal_4202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C ( clk ), .D ( new_AGEMA_signal_4209 ), .Q ( new_AGEMA_signal_4210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C ( clk ), .D ( new_AGEMA_signal_4213 ), .Q ( new_AGEMA_signal_4214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C ( clk ), .D ( new_AGEMA_signal_4217 ), .Q ( new_AGEMA_signal_4218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C ( clk ), .D ( new_AGEMA_signal_4221 ), .Q ( new_AGEMA_signal_4222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C ( clk ), .D ( new_AGEMA_signal_4225 ), .Q ( new_AGEMA_signal_4226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C ( clk ), .D ( new_AGEMA_signal_4229 ), .Q ( new_AGEMA_signal_4230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C ( clk ), .D ( new_AGEMA_signal_4233 ), .Q ( new_AGEMA_signal_4234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C ( clk ), .D ( new_AGEMA_signal_4237 ), .Q ( new_AGEMA_signal_4238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C ( clk ), .D ( new_AGEMA_signal_4241 ), .Q ( new_AGEMA_signal_4242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C ( clk ), .D ( new_AGEMA_signal_4245 ), .Q ( new_AGEMA_signal_4246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C ( clk ), .D ( new_AGEMA_signal_4253 ), .Q ( new_AGEMA_signal_4254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C ( clk ), .D ( new_AGEMA_signal_4261 ), .Q ( new_AGEMA_signal_4262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C ( clk ), .D ( new_AGEMA_signal_4269 ), .Q ( new_AGEMA_signal_4270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C ( clk ), .D ( new_AGEMA_signal_4273 ), .Q ( new_AGEMA_signal_4274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C ( clk ), .D ( new_AGEMA_signal_4283 ), .Q ( new_AGEMA_signal_4284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C ( clk ), .D ( new_AGEMA_signal_4289 ), .Q ( new_AGEMA_signal_4290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C ( clk ), .D ( new_AGEMA_signal_4299 ), .Q ( new_AGEMA_signal_4300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C ( clk ), .D ( new_AGEMA_signal_4307 ), .Q ( new_AGEMA_signal_4308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C ( clk ), .D ( new_AGEMA_signal_4327 ), .Q ( new_AGEMA_signal_4328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C ( clk ), .D ( new_AGEMA_signal_4335 ), .Q ( new_AGEMA_signal_4336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C ( clk ), .D ( new_AGEMA_signal_4345 ), .Q ( new_AGEMA_signal_4346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C ( clk ), .D ( new_AGEMA_signal_4351 ), .Q ( new_AGEMA_signal_4352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C ( clk ), .D ( new_AGEMA_signal_4367 ), .Q ( new_AGEMA_signal_4368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C ( clk ), .D ( new_AGEMA_signal_4375 ), .Q ( new_AGEMA_signal_4376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C ( clk ), .D ( new_AGEMA_signal_4389 ), .Q ( new_AGEMA_signal_4390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C ( clk ), .D ( new_AGEMA_signal_4395 ), .Q ( new_AGEMA_signal_4396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C ( clk ), .D ( new_AGEMA_signal_4401 ), .Q ( new_AGEMA_signal_4402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C ( clk ), .D ( new_AGEMA_signal_4407 ), .Q ( new_AGEMA_signal_4408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C ( clk ), .D ( new_AGEMA_signal_4413 ), .Q ( new_AGEMA_signal_4414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C ( clk ), .D ( new_AGEMA_signal_4419 ), .Q ( new_AGEMA_signal_4420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C ( clk ), .D ( new_AGEMA_signal_4425 ), .Q ( new_AGEMA_signal_4426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C ( clk ), .D ( new_AGEMA_signal_4431 ), .Q ( new_AGEMA_signal_4432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C ( clk ), .D ( new_AGEMA_signal_4437 ), .Q ( new_AGEMA_signal_4438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C ( clk ), .D ( new_AGEMA_signal_4443 ), .Q ( new_AGEMA_signal_4444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C ( clk ), .D ( new_AGEMA_signal_4459 ), .Q ( new_AGEMA_signal_4460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C ( clk ), .D ( new_AGEMA_signal_4467 ), .Q ( new_AGEMA_signal_4468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C ( clk ), .D ( new_AGEMA_signal_4481 ), .Q ( new_AGEMA_signal_4482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C ( clk ), .D ( new_AGEMA_signal_4487 ), .Q ( new_AGEMA_signal_4488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C ( clk ), .D ( new_AGEMA_signal_4495 ), .Q ( new_AGEMA_signal_4496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C ( clk ), .D ( new_AGEMA_signal_4503 ), .Q ( new_AGEMA_signal_4504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C ( clk ), .D ( new_AGEMA_signal_4513 ), .Q ( new_AGEMA_signal_4514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C ( clk ), .D ( new_AGEMA_signal_4519 ), .Q ( new_AGEMA_signal_4520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C ( clk ), .D ( new_AGEMA_signal_4533 ), .Q ( new_AGEMA_signal_4534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C ( clk ), .D ( new_AGEMA_signal_4539 ), .Q ( new_AGEMA_signal_4540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C ( clk ), .D ( new_AGEMA_signal_4545 ), .Q ( new_AGEMA_signal_4546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C ( clk ), .D ( new_AGEMA_signal_4551 ), .Q ( new_AGEMA_signal_4552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C ( clk ), .D ( new_AGEMA_signal_4559 ), .Q ( new_AGEMA_signal_4560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C ( clk ), .D ( new_AGEMA_signal_4567 ), .Q ( new_AGEMA_signal_4568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C ( clk ), .D ( new_AGEMA_signal_4575 ), .Q ( new_AGEMA_signal_4576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C ( clk ), .D ( new_AGEMA_signal_4583 ), .Q ( new_AGEMA_signal_4584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C ( clk ), .D ( new_AGEMA_signal_4589 ), .Q ( new_AGEMA_signal_4590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C ( clk ), .D ( new_AGEMA_signal_4595 ), .Q ( new_AGEMA_signal_4596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C ( clk ), .D ( new_AGEMA_signal_4601 ), .Q ( new_AGEMA_signal_4602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C ( clk ), .D ( new_AGEMA_signal_4607 ), .Q ( new_AGEMA_signal_4608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C ( clk ), .D ( new_AGEMA_signal_4669 ), .Q ( new_AGEMA_signal_4670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C ( clk ), .D ( new_AGEMA_signal_4677 ), .Q ( new_AGEMA_signal_4678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C ( clk ), .D ( new_AGEMA_signal_4685 ), .Q ( new_AGEMA_signal_4686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C ( clk ), .D ( new_AGEMA_signal_4693 ), .Q ( new_AGEMA_signal_4694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C ( clk ), .D ( new_AGEMA_signal_4701 ), .Q ( new_AGEMA_signal_4702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C ( clk ), .D ( new_AGEMA_signal_4709 ), .Q ( new_AGEMA_signal_4710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C ( clk ), .D ( new_AGEMA_signal_4717 ), .Q ( new_AGEMA_signal_4718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C ( clk ), .D ( new_AGEMA_signal_4725 ), .Q ( new_AGEMA_signal_4726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C ( clk ), .D ( new_AGEMA_signal_4747 ), .Q ( new_AGEMA_signal_4748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C ( clk ), .D ( new_AGEMA_signal_4757 ), .Q ( new_AGEMA_signal_4758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C ( clk ), .D ( new_AGEMA_signal_4765 ), .Q ( new_AGEMA_signal_4766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C ( clk ), .D ( new_AGEMA_signal_4773 ), .Q ( new_AGEMA_signal_4774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C ( clk ), .D ( new_AGEMA_signal_4781 ), .Q ( new_AGEMA_signal_4782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C ( clk ), .D ( new_AGEMA_signal_4789 ), .Q ( new_AGEMA_signal_4790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C ( clk ), .D ( new_AGEMA_signal_4797 ), .Q ( new_AGEMA_signal_4798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C ( clk ), .D ( new_AGEMA_signal_4805 ), .Q ( new_AGEMA_signal_4806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C ( clk ), .D ( new_AGEMA_signal_4847 ), .Q ( new_AGEMA_signal_4848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C ( clk ), .D ( new_AGEMA_signal_4857 ), .Q ( new_AGEMA_signal_4858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C ( clk ), .D ( new_AGEMA_signal_4865 ), .Q ( new_AGEMA_signal_4866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C ( clk ), .D ( new_AGEMA_signal_4873 ), .Q ( new_AGEMA_signal_4874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C ( clk ), .D ( new_AGEMA_signal_4893 ), .Q ( new_AGEMA_signal_4894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C ( clk ), .D ( new_AGEMA_signal_4901 ), .Q ( new_AGEMA_signal_4902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C ( clk ), .D ( new_AGEMA_signal_4909 ), .Q ( new_AGEMA_signal_4910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C ( clk ), .D ( new_AGEMA_signal_4917 ), .Q ( new_AGEMA_signal_4918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C ( clk ), .D ( new_AGEMA_signal_4945 ), .Q ( new_AGEMA_signal_4946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C ( clk ), .D ( new_AGEMA_signal_4953 ), .Q ( new_AGEMA_signal_4954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C ( clk ), .D ( new_AGEMA_signal_5077 ), .Q ( new_AGEMA_signal_5078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C ( clk ), .D ( new_AGEMA_signal_5087 ), .Q ( new_AGEMA_signal_5088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C ( clk ), .D ( new_AGEMA_signal_5469 ), .Q ( new_AGEMA_signal_5470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C ( clk ), .D ( new_AGEMA_signal_5483 ), .Q ( new_AGEMA_signal_5484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C ( clk ), .D ( new_AGEMA_signal_5513 ), .Q ( new_AGEMA_signal_5514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C ( clk ), .D ( new_AGEMA_signal_5527 ), .Q ( new_AGEMA_signal_5528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C ( clk ), .D ( new_AGEMA_signal_5585 ), .Q ( new_AGEMA_signal_5586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C ( clk ), .D ( new_AGEMA_signal_5601 ), .Q ( new_AGEMA_signal_5602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C ( clk ), .D ( new_AGEMA_signal_5629 ), .Q ( new_AGEMA_signal_5630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C ( clk ), .D ( new_AGEMA_signal_5645 ), .Q ( new_AGEMA_signal_5646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C ( clk ), .D ( new_AGEMA_signal_5781 ), .Q ( new_AGEMA_signal_5782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C ( clk ), .D ( new_AGEMA_signal_5799 ), .Q ( new_AGEMA_signal_5800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C ( clk ), .D ( new_AGEMA_signal_5881 ), .Q ( new_AGEMA_signal_5882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C ( clk ), .D ( new_AGEMA_signal_5901 ), .Q ( new_AGEMA_signal_5902 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_2013 ( .C ( clk ), .D ( new_AGEMA_signal_3830 ), .Q ( new_AGEMA_signal_3831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C ( clk ), .D ( new_AGEMA_signal_3834 ), .Q ( new_AGEMA_signal_3835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C ( clk ), .D ( new_AGEMA_signal_3838 ), .Q ( new_AGEMA_signal_3839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C ( clk ), .D ( new_AGEMA_signal_3842 ), .Q ( new_AGEMA_signal_3843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C ( clk ), .D ( new_AGEMA_signal_3850 ), .Q ( new_AGEMA_signal_3851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C ( clk ), .D ( new_AGEMA_signal_3858 ), .Q ( new_AGEMA_signal_3859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C ( clk ), .D ( n1978 ), .Q ( new_AGEMA_signal_3861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C ( clk ), .D ( new_AGEMA_signal_1482 ), .Q ( new_AGEMA_signal_3863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C ( clk ), .D ( new_AGEMA_signal_3870 ), .Q ( new_AGEMA_signal_3871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C ( clk ), .D ( new_AGEMA_signal_3878 ), .Q ( new_AGEMA_signal_3879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C ( clk ), .D ( new_AGEMA_signal_3884 ), .Q ( new_AGEMA_signal_3885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C ( clk ), .D ( new_AGEMA_signal_3890 ), .Q ( new_AGEMA_signal_3891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C ( clk ), .D ( new_AGEMA_signal_3894 ), .Q ( new_AGEMA_signal_3895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C ( clk ), .D ( new_AGEMA_signal_3898 ), .Q ( new_AGEMA_signal_3899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C ( clk ), .D ( new_AGEMA_signal_3904 ), .Q ( new_AGEMA_signal_3905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C ( clk ), .D ( new_AGEMA_signal_3910 ), .Q ( new_AGEMA_signal_3911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C ( clk ), .D ( new_AGEMA_signal_3720 ), .Q ( new_AGEMA_signal_3913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C ( clk ), .D ( new_AGEMA_signal_3724 ), .Q ( new_AGEMA_signal_3915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C ( clk ), .D ( new_AGEMA_signal_3920 ), .Q ( new_AGEMA_signal_3921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C ( clk ), .D ( new_AGEMA_signal_3926 ), .Q ( new_AGEMA_signal_3927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C ( clk ), .D ( new_AGEMA_signal_3932 ), .Q ( new_AGEMA_signal_3933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C ( clk ), .D ( new_AGEMA_signal_3938 ), .Q ( new_AGEMA_signal_3939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C ( clk ), .D ( n2091 ), .Q ( new_AGEMA_signal_3941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C ( clk ), .D ( new_AGEMA_signal_1500 ), .Q ( new_AGEMA_signal_3943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C ( clk ), .D ( new_AGEMA_signal_3946 ), .Q ( new_AGEMA_signal_3947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C ( clk ), .D ( new_AGEMA_signal_3950 ), .Q ( new_AGEMA_signal_3951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C ( clk ), .D ( new_AGEMA_signal_3956 ), .Q ( new_AGEMA_signal_3957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C ( clk ), .D ( new_AGEMA_signal_3962 ), .Q ( new_AGEMA_signal_3963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C ( clk ), .D ( new_AGEMA_signal_3968 ), .Q ( new_AGEMA_signal_3969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C ( clk ), .D ( new_AGEMA_signal_3974 ), .Q ( new_AGEMA_signal_3975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C ( clk ), .D ( n2543 ), .Q ( new_AGEMA_signal_3977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C ( clk ), .D ( new_AGEMA_signal_1506 ), .Q ( new_AGEMA_signal_3979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C ( clk ), .D ( new_AGEMA_signal_3984 ), .Q ( new_AGEMA_signal_3985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C ( clk ), .D ( new_AGEMA_signal_3990 ), .Q ( new_AGEMA_signal_3991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C ( clk ), .D ( n2159 ), .Q ( new_AGEMA_signal_3993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C ( clk ), .D ( new_AGEMA_signal_1510 ), .Q ( new_AGEMA_signal_3995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C ( clk ), .D ( new_AGEMA_signal_3998 ), .Q ( new_AGEMA_signal_3999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C ( clk ), .D ( new_AGEMA_signal_4002 ), .Q ( new_AGEMA_signal_4003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C ( clk ), .D ( new_AGEMA_signal_4006 ), .Q ( new_AGEMA_signal_4007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C ( clk ), .D ( new_AGEMA_signal_4010 ), .Q ( new_AGEMA_signal_4011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C ( clk ), .D ( new_AGEMA_signal_3706 ), .Q ( new_AGEMA_signal_4013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C ( clk ), .D ( new_AGEMA_signal_3708 ), .Q ( new_AGEMA_signal_4015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C ( clk ), .D ( new_AGEMA_signal_4022 ), .Q ( new_AGEMA_signal_4023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C ( clk ), .D ( new_AGEMA_signal_4030 ), .Q ( new_AGEMA_signal_4031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C ( clk ), .D ( new_AGEMA_signal_4036 ), .Q ( new_AGEMA_signal_4037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C ( clk ), .D ( new_AGEMA_signal_4042 ), .Q ( new_AGEMA_signal_4043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C ( clk ), .D ( new_AGEMA_signal_4046 ), .Q ( new_AGEMA_signal_4047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C ( clk ), .D ( new_AGEMA_signal_4050 ), .Q ( new_AGEMA_signal_4051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C ( clk ), .D ( new_AGEMA_signal_4054 ), .Q ( new_AGEMA_signal_4055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C ( clk ), .D ( new_AGEMA_signal_4058 ), .Q ( new_AGEMA_signal_4059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C ( clk ), .D ( n2270 ), .Q ( new_AGEMA_signal_4061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C ( clk ), .D ( new_AGEMA_signal_1386 ), .Q ( new_AGEMA_signal_4063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C ( clk ), .D ( n2285 ), .Q ( new_AGEMA_signal_4065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C ( clk ), .D ( new_AGEMA_signal_1528 ), .Q ( new_AGEMA_signal_4067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C ( clk ), .D ( new_AGEMA_signal_4070 ), .Q ( new_AGEMA_signal_4071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C ( clk ), .D ( new_AGEMA_signal_4074 ), .Q ( new_AGEMA_signal_4075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C ( clk ), .D ( new_AGEMA_signal_4078 ), .Q ( new_AGEMA_signal_4079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C ( clk ), .D ( new_AGEMA_signal_4082 ), .Q ( new_AGEMA_signal_4083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C ( clk ), .D ( n2334 ), .Q ( new_AGEMA_signal_4085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C ( clk ), .D ( new_AGEMA_signal_1397 ), .Q ( new_AGEMA_signal_4087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C ( clk ), .D ( new_AGEMA_signal_4092 ), .Q ( new_AGEMA_signal_4093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C ( clk ), .D ( new_AGEMA_signal_4098 ), .Q ( new_AGEMA_signal_4099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C ( clk ), .D ( new_AGEMA_signal_4102 ), .Q ( new_AGEMA_signal_4103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C ( clk ), .D ( new_AGEMA_signal_4106 ), .Q ( new_AGEMA_signal_4107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C ( clk ), .D ( new_AGEMA_signal_3714 ), .Q ( new_AGEMA_signal_4109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C ( clk ), .D ( new_AGEMA_signal_3716 ), .Q ( new_AGEMA_signal_4111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C ( clk ), .D ( new_AGEMA_signal_4114 ), .Q ( new_AGEMA_signal_4115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C ( clk ), .D ( new_AGEMA_signal_4118 ), .Q ( new_AGEMA_signal_4119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C ( clk ), .D ( new_AGEMA_signal_4122 ), .Q ( new_AGEMA_signal_4123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C ( clk ), .D ( new_AGEMA_signal_4126 ), .Q ( new_AGEMA_signal_4127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C ( clk ), .D ( new_AGEMA_signal_4130 ), .Q ( new_AGEMA_signal_4131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C ( clk ), .D ( new_AGEMA_signal_4134 ), .Q ( new_AGEMA_signal_4135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C ( clk ), .D ( n2435 ), .Q ( new_AGEMA_signal_4137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C ( clk ), .D ( new_AGEMA_signal_1416 ), .Q ( new_AGEMA_signal_4139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C ( clk ), .D ( new_AGEMA_signal_4142 ), .Q ( new_AGEMA_signal_4143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C ( clk ), .D ( new_AGEMA_signal_4146 ), .Q ( new_AGEMA_signal_4147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C ( clk ), .D ( new_AGEMA_signal_3638 ), .Q ( new_AGEMA_signal_4149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C ( clk ), .D ( new_AGEMA_signal_3640 ), .Q ( new_AGEMA_signal_4151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C ( clk ), .D ( new_AGEMA_signal_4156 ), .Q ( new_AGEMA_signal_4157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C ( clk ), .D ( new_AGEMA_signal_4162 ), .Q ( new_AGEMA_signal_4163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C ( clk ), .D ( new_AGEMA_signal_4168 ), .Q ( new_AGEMA_signal_4169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C ( clk ), .D ( new_AGEMA_signal_4174 ), .Q ( new_AGEMA_signal_4175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C ( clk ), .D ( new_AGEMA_signal_4178 ), .Q ( new_AGEMA_signal_4179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C ( clk ), .D ( new_AGEMA_signal_4182 ), .Q ( new_AGEMA_signal_4183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C ( clk ), .D ( new_AGEMA_signal_3618 ), .Q ( new_AGEMA_signal_4185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C ( clk ), .D ( new_AGEMA_signal_3624 ), .Q ( new_AGEMA_signal_4187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C ( clk ), .D ( new_AGEMA_signal_4194 ), .Q ( new_AGEMA_signal_4195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C ( clk ), .D ( new_AGEMA_signal_4202 ), .Q ( new_AGEMA_signal_4203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C ( clk ), .D ( n2547 ), .Q ( new_AGEMA_signal_4205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C ( clk ), .D ( new_AGEMA_signal_1434 ), .Q ( new_AGEMA_signal_4207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C ( clk ), .D ( new_AGEMA_signal_4210 ), .Q ( new_AGEMA_signal_4211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C ( clk ), .D ( new_AGEMA_signal_4214 ), .Q ( new_AGEMA_signal_4215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C ( clk ), .D ( new_AGEMA_signal_4218 ), .Q ( new_AGEMA_signal_4219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C ( clk ), .D ( new_AGEMA_signal_4222 ), .Q ( new_AGEMA_signal_4223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C ( clk ), .D ( new_AGEMA_signal_4226 ), .Q ( new_AGEMA_signal_4227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C ( clk ), .D ( new_AGEMA_signal_4230 ), .Q ( new_AGEMA_signal_4231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C ( clk ), .D ( new_AGEMA_signal_4234 ), .Q ( new_AGEMA_signal_4235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C ( clk ), .D ( new_AGEMA_signal_4238 ), .Q ( new_AGEMA_signal_4239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C ( clk ), .D ( new_AGEMA_signal_4242 ), .Q ( new_AGEMA_signal_4243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C ( clk ), .D ( new_AGEMA_signal_4246 ), .Q ( new_AGEMA_signal_4247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C ( clk ), .D ( new_AGEMA_signal_4254 ), .Q ( new_AGEMA_signal_4255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C ( clk ), .D ( new_AGEMA_signal_4262 ), .Q ( new_AGEMA_signal_4263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C ( clk ), .D ( n2758 ), .Q ( new_AGEMA_signal_4265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C ( clk ), .D ( new_AGEMA_signal_1579 ), .Q ( new_AGEMA_signal_4267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C ( clk ), .D ( new_AGEMA_signal_4270 ), .Q ( new_AGEMA_signal_4271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C ( clk ), .D ( new_AGEMA_signal_4274 ), .Q ( new_AGEMA_signal_4275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C ( clk ), .D ( n2797 ), .Q ( new_AGEMA_signal_4277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C ( clk ), .D ( new_AGEMA_signal_1583 ), .Q ( new_AGEMA_signal_4279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C ( clk ), .D ( new_AGEMA_signal_4284 ), .Q ( new_AGEMA_signal_4285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C ( clk ), .D ( new_AGEMA_signal_4290 ), .Q ( new_AGEMA_signal_4291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C ( clk ), .D ( new_AGEMA_signal_4300 ), .Q ( new_AGEMA_signal_4301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C ( clk ), .D ( new_AGEMA_signal_4308 ), .Q ( new_AGEMA_signal_4309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C ( clk ), .D ( n2012 ), .Q ( new_AGEMA_signal_4317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C ( clk ), .D ( new_AGEMA_signal_1487 ), .Q ( new_AGEMA_signal_4321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C ( clk ), .D ( new_AGEMA_signal_4328 ), .Q ( new_AGEMA_signal_4329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C ( clk ), .D ( new_AGEMA_signal_4336 ), .Q ( new_AGEMA_signal_4337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C ( clk ), .D ( new_AGEMA_signal_4346 ), .Q ( new_AGEMA_signal_4347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C ( clk ), .D ( new_AGEMA_signal_4352 ), .Q ( new_AGEMA_signal_4353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C ( clk ), .D ( n2652 ), .Q ( new_AGEMA_signal_4357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C ( clk ), .D ( new_AGEMA_signal_1496 ), .Q ( new_AGEMA_signal_4361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C ( clk ), .D ( new_AGEMA_signal_4368 ), .Q ( new_AGEMA_signal_4369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C ( clk ), .D ( new_AGEMA_signal_4376 ), .Q ( new_AGEMA_signal_4377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C ( clk ), .D ( n2143 ), .Q ( new_AGEMA_signal_4381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C ( clk ), .D ( new_AGEMA_signal_1508 ), .Q ( new_AGEMA_signal_4385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C ( clk ), .D ( new_AGEMA_signal_4390 ), .Q ( new_AGEMA_signal_4391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C ( clk ), .D ( new_AGEMA_signal_4396 ), .Q ( new_AGEMA_signal_4397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C ( clk ), .D ( new_AGEMA_signal_4402 ), .Q ( new_AGEMA_signal_4403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C ( clk ), .D ( new_AGEMA_signal_4408 ), .Q ( new_AGEMA_signal_4409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C ( clk ), .D ( new_AGEMA_signal_4414 ), .Q ( new_AGEMA_signal_4415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C ( clk ), .D ( new_AGEMA_signal_4420 ), .Q ( new_AGEMA_signal_4421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C ( clk ), .D ( new_AGEMA_signal_4426 ), .Q ( new_AGEMA_signal_4427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C ( clk ), .D ( new_AGEMA_signal_4432 ), .Q ( new_AGEMA_signal_4433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C ( clk ), .D ( new_AGEMA_signal_4438 ), .Q ( new_AGEMA_signal_4439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C ( clk ), .D ( new_AGEMA_signal_4444 ), .Q ( new_AGEMA_signal_4445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C ( clk ), .D ( n2297 ), .Q ( new_AGEMA_signal_4449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C ( clk ), .D ( new_AGEMA_signal_1531 ), .Q ( new_AGEMA_signal_4453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C ( clk ), .D ( new_AGEMA_signal_4460 ), .Q ( new_AGEMA_signal_4461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C ( clk ), .D ( new_AGEMA_signal_4468 ), .Q ( new_AGEMA_signal_4469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C ( clk ), .D ( n2336 ), .Q ( new_AGEMA_signal_4473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C ( clk ), .D ( new_AGEMA_signal_1626 ), .Q ( new_AGEMA_signal_4477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C ( clk ), .D ( new_AGEMA_signal_4482 ), .Q ( new_AGEMA_signal_4483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C ( clk ), .D ( new_AGEMA_signal_4488 ), .Q ( new_AGEMA_signal_4489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C ( clk ), .D ( new_AGEMA_signal_4496 ), .Q ( new_AGEMA_signal_4497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C ( clk ), .D ( new_AGEMA_signal_4504 ), .Q ( new_AGEMA_signal_4505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C ( clk ), .D ( new_AGEMA_signal_4514 ), .Q ( new_AGEMA_signal_4515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C ( clk ), .D ( new_AGEMA_signal_4520 ), .Q ( new_AGEMA_signal_4521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C ( clk ), .D ( new_AGEMA_signal_4534 ), .Q ( new_AGEMA_signal_4535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C ( clk ), .D ( new_AGEMA_signal_4540 ), .Q ( new_AGEMA_signal_4541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C ( clk ), .D ( new_AGEMA_signal_4546 ), .Q ( new_AGEMA_signal_4547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C ( clk ), .D ( new_AGEMA_signal_4552 ), .Q ( new_AGEMA_signal_4553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C ( clk ), .D ( new_AGEMA_signal_4560 ), .Q ( new_AGEMA_signal_4561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C ( clk ), .D ( new_AGEMA_signal_4568 ), .Q ( new_AGEMA_signal_4569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C ( clk ), .D ( new_AGEMA_signal_4576 ), .Q ( new_AGEMA_signal_4577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C ( clk ), .D ( new_AGEMA_signal_4584 ), .Q ( new_AGEMA_signal_4585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C ( clk ), .D ( new_AGEMA_signal_4590 ), .Q ( new_AGEMA_signal_4591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C ( clk ), .D ( new_AGEMA_signal_4596 ), .Q ( new_AGEMA_signal_4597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C ( clk ), .D ( new_AGEMA_signal_4602 ), .Q ( new_AGEMA_signal_4603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C ( clk ), .D ( new_AGEMA_signal_4608 ), .Q ( new_AGEMA_signal_4609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C ( clk ), .D ( n2658 ), .Q ( new_AGEMA_signal_4617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C ( clk ), .D ( new_AGEMA_signal_1478 ), .Q ( new_AGEMA_signal_4621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C ( clk ), .D ( n2698 ), .Q ( new_AGEMA_signal_4625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C ( clk ), .D ( new_AGEMA_signal_1573 ), .Q ( new_AGEMA_signal_4629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C ( clk ), .D ( n2800 ), .Q ( new_AGEMA_signal_4633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C ( clk ), .D ( new_AGEMA_signal_1581 ), .Q ( new_AGEMA_signal_4637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C ( clk ), .D ( n1936 ), .Q ( new_AGEMA_signal_4645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C ( clk ), .D ( new_AGEMA_signal_1470 ), .Q ( new_AGEMA_signal_4651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C ( clk ), .D ( new_AGEMA_signal_4670 ), .Q ( new_AGEMA_signal_4671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C ( clk ), .D ( new_AGEMA_signal_4678 ), .Q ( new_AGEMA_signal_4679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C ( clk ), .D ( new_AGEMA_signal_4686 ), .Q ( new_AGEMA_signal_4687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C ( clk ), .D ( new_AGEMA_signal_4694 ), .Q ( new_AGEMA_signal_4695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C ( clk ), .D ( new_AGEMA_signal_4702 ), .Q ( new_AGEMA_signal_4703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C ( clk ), .D ( new_AGEMA_signal_4710 ), .Q ( new_AGEMA_signal_4711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C ( clk ), .D ( new_AGEMA_signal_4718 ), .Q ( new_AGEMA_signal_4719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C ( clk ), .D ( new_AGEMA_signal_4726 ), .Q ( new_AGEMA_signal_4727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C ( clk ), .D ( n2099 ), .Q ( new_AGEMA_signal_4733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C ( clk ), .D ( new_AGEMA_signal_1499 ), .Q ( new_AGEMA_signal_4739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C ( clk ), .D ( new_AGEMA_signal_4748 ), .Q ( new_AGEMA_signal_4749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C ( clk ), .D ( new_AGEMA_signal_4758 ), .Q ( new_AGEMA_signal_4759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C ( clk ), .D ( new_AGEMA_signal_4766 ), .Q ( new_AGEMA_signal_4767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C ( clk ), .D ( new_AGEMA_signal_4774 ), .Q ( new_AGEMA_signal_4775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C ( clk ), .D ( new_AGEMA_signal_4782 ), .Q ( new_AGEMA_signal_4783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C ( clk ), .D ( new_AGEMA_signal_4790 ), .Q ( new_AGEMA_signal_4791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C ( clk ), .D ( new_AGEMA_signal_4798 ), .Q ( new_AGEMA_signal_4799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C ( clk ), .D ( new_AGEMA_signal_4806 ), .Q ( new_AGEMA_signal_4807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C ( clk ), .D ( n2301 ), .Q ( new_AGEMA_signal_4825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C ( clk ), .D ( new_AGEMA_signal_1533 ), .Q ( new_AGEMA_signal_4831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C ( clk ), .D ( new_AGEMA_signal_4848 ), .Q ( new_AGEMA_signal_4849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C ( clk ), .D ( new_AGEMA_signal_4858 ), .Q ( new_AGEMA_signal_4859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C ( clk ), .D ( new_AGEMA_signal_4866 ), .Q ( new_AGEMA_signal_4867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C ( clk ), .D ( new_AGEMA_signal_4874 ), .Q ( new_AGEMA_signal_4875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C ( clk ), .D ( new_AGEMA_signal_4894 ), .Q ( new_AGEMA_signal_4895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C ( clk ), .D ( new_AGEMA_signal_4902 ), .Q ( new_AGEMA_signal_4903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C ( clk ), .D ( new_AGEMA_signal_4910 ), .Q ( new_AGEMA_signal_4911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C ( clk ), .D ( new_AGEMA_signal_4918 ), .Q ( new_AGEMA_signal_4919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C ( clk ), .D ( new_AGEMA_signal_3584 ), .Q ( new_AGEMA_signal_4925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C ( clk ), .D ( new_AGEMA_signal_3588 ), .Q ( new_AGEMA_signal_4931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C ( clk ), .D ( new_AGEMA_signal_4946 ), .Q ( new_AGEMA_signal_4947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C ( clk ), .D ( new_AGEMA_signal_4954 ), .Q ( new_AGEMA_signal_4955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C ( clk ), .D ( new_AGEMA_signal_3808 ), .Q ( new_AGEMA_signal_5009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C ( clk ), .D ( new_AGEMA_signal_3812 ), .Q ( new_AGEMA_signal_5017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C ( clk ), .D ( n2102 ), .Q ( new_AGEMA_signal_5045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C ( clk ), .D ( new_AGEMA_signal_1503 ), .Q ( new_AGEMA_signal_5053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C ( clk ), .D ( new_AGEMA_signal_3502 ), .Q ( new_AGEMA_signal_5061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C ( clk ), .D ( new_AGEMA_signal_3504 ), .Q ( new_AGEMA_signal_5069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C ( clk ), .D ( new_AGEMA_signal_5078 ), .Q ( new_AGEMA_signal_5079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C ( clk ), .D ( new_AGEMA_signal_5088 ), .Q ( new_AGEMA_signal_5089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C ( clk ), .D ( new_AGEMA_signal_3688 ), .Q ( new_AGEMA_signal_5097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C ( clk ), .D ( new_AGEMA_signal_3692 ), .Q ( new_AGEMA_signal_5105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C ( clk ), .D ( n2367 ), .Q ( new_AGEMA_signal_5145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C ( clk ), .D ( new_AGEMA_signal_1400 ), .Q ( new_AGEMA_signal_5153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C ( clk ), .D ( n2591 ), .Q ( new_AGEMA_signal_5177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C ( clk ), .D ( new_AGEMA_signal_1564 ), .Q ( new_AGEMA_signal_5185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C ( clk ), .D ( n2105 ), .Q ( new_AGEMA_signal_5265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C ( clk ), .D ( new_AGEMA_signal_1498 ), .Q ( new_AGEMA_signal_5275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C ( clk ), .D ( n2106 ), .Q ( new_AGEMA_signal_5445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C ( clk ), .D ( new_AGEMA_signal_1357 ), .Q ( new_AGEMA_signal_5457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C ( clk ), .D ( new_AGEMA_signal_5470 ), .Q ( new_AGEMA_signal_5471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C ( clk ), .D ( new_AGEMA_signal_5484 ), .Q ( new_AGEMA_signal_5485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C ( clk ), .D ( new_AGEMA_signal_5514 ), .Q ( new_AGEMA_signal_5515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C ( clk ), .D ( new_AGEMA_signal_5528 ), .Q ( new_AGEMA_signal_5529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C ( clk ), .D ( new_AGEMA_signal_5586 ), .Q ( new_AGEMA_signal_5587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C ( clk ), .D ( new_AGEMA_signal_5602 ), .Q ( new_AGEMA_signal_5603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C ( clk ), .D ( new_AGEMA_signal_5630 ), .Q ( new_AGEMA_signal_5631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C ( clk ), .D ( new_AGEMA_signal_5646 ), .Q ( new_AGEMA_signal_5647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C ( clk ), .D ( n2155 ), .Q ( new_AGEMA_signal_5729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C ( clk ), .D ( new_AGEMA_signal_1359 ), .Q ( new_AGEMA_signal_5745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C ( clk ), .D ( new_AGEMA_signal_5782 ), .Q ( new_AGEMA_signal_5783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C ( clk ), .D ( new_AGEMA_signal_5800 ), .Q ( new_AGEMA_signal_5801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C ( clk ), .D ( new_AGEMA_signal_5882 ), .Q ( new_AGEMA_signal_5883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C ( clk ), .D ( new_AGEMA_signal_5902 ), .Q ( new_AGEMA_signal_5903 ) ) ;

    /* cells in depth 10 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1983 ( .a ({new_AGEMA_signal_3432, new_AGEMA_signal_3428}), .b ({new_AGEMA_signal_1471, n1928}), .clk ( clk ), .r ( Fresh[575] ), .c ({new_AGEMA_signal_1585, n1934}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U1998 ( .a ({new_AGEMA_signal_1472, n1931}), .b ({new_AGEMA_signal_3440, new_AGEMA_signal_3436}), .clk ( clk ), .r ( Fresh[576] ), .c ({new_AGEMA_signal_1586, n1932}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2015 ( .a ({new_AGEMA_signal_1473, n1939}), .b ({new_AGEMA_signal_3444, new_AGEMA_signal_3442}), .clk ( clk ), .r ( Fresh[577] ), .c ({new_AGEMA_signal_1587, n1940}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2033 ( .a ({new_AGEMA_signal_1474, n1948}), .b ({new_AGEMA_signal_1475, n1947}), .clk ( clk ), .r ( Fresh[578] ), .c ({new_AGEMA_signal_1588, n1961}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2050 ( .a ({new_AGEMA_signal_1476, n1954}), .b ({new_AGEMA_signal_1477, n1953}), .clk ( clk ), .r ( Fresh[579] ), .c ({new_AGEMA_signal_1589, n1955}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2066 ( .a ({new_AGEMA_signal_3448, new_AGEMA_signal_3446}), .b ({new_AGEMA_signal_1322, n1965}), .clk ( clk ), .r ( Fresh[580] ), .c ({new_AGEMA_signal_1479, n1967}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2085 ( .a ({new_AGEMA_signal_1591, n1970}), .b ({new_AGEMA_signal_1481, n1969}), .clk ( clk ), .r ( Fresh[581] ), .c ({new_AGEMA_signal_1669, n1984}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2103 ( .a ({new_AGEMA_signal_3456, new_AGEMA_signal_3452}), .b ({new_AGEMA_signal_1483, n1975}), .clk ( clk ), .r ( Fresh[582] ), .c ({new_AGEMA_signal_1592, n1977}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2108 ( .a ({new_AGEMA_signal_3460, new_AGEMA_signal_3458}), .b ({new_AGEMA_signal_1484, n1980}), .clk ( clk ), .r ( Fresh[583] ), .c ({new_AGEMA_signal_1593, n1981}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2115 ( .a ({new_AGEMA_signal_3468, new_AGEMA_signal_3464}), .b ({new_AGEMA_signal_1329, n1986}), .clk ( clk ), .r ( Fresh[584] ), .c ({new_AGEMA_signal_1485, n1987}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2127 ( .a ({new_AGEMA_signal_1486, n1997}), .b ({new_AGEMA_signal_3472, new_AGEMA_signal_3470}), .clk ( clk ), .r ( Fresh[585] ), .c ({new_AGEMA_signal_1594, n1998}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2146 ( .a ({new_AGEMA_signal_3480, new_AGEMA_signal_3476}), .b ({new_AGEMA_signal_1488, n2007}), .clk ( clk ), .r ( Fresh[586] ), .c ({new_AGEMA_signal_1595, n2010}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2162 ( .a ({new_AGEMA_signal_3488, new_AGEMA_signal_3484}), .b ({new_AGEMA_signal_1336, n2021}), .clk ( clk ), .r ( Fresh[587] ), .c ({new_AGEMA_signal_1489, n2024}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2177 ( .a ({new_AGEMA_signal_3492, new_AGEMA_signal_3490}), .b ({new_AGEMA_signal_1490, n2032}), .clk ( clk ), .r ( Fresh[588] ), .c ({new_AGEMA_signal_1597, n2035}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2186 ( .a ({new_AGEMA_signal_1491, n2041}), .b ({new_AGEMA_signal_3496, new_AGEMA_signal_3494}), .clk ( clk ), .r ( Fresh[589] ), .c ({new_AGEMA_signal_1598, n2054}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2190 ( .a ({new_AGEMA_signal_3500, new_AGEMA_signal_3498}), .b ({new_AGEMA_signal_1492, n2043}), .clk ( clk ), .r ( Fresh[590] ), .c ({new_AGEMA_signal_1599, n2048}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2195 ( .a ({new_AGEMA_signal_1493, n2046}), .b ({new_AGEMA_signal_3504, new_AGEMA_signal_3502}), .clk ( clk ), .r ( Fresh[591] ), .c ({new_AGEMA_signal_1600, n2047}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2206 ( .a ({new_AGEMA_signal_1494, n2058}), .b ({new_AGEMA_signal_3512, new_AGEMA_signal_3508}), .clk ( clk ), .r ( Fresh[592] ), .c ({new_AGEMA_signal_1601, n2059}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2213 ( .a ({new_AGEMA_signal_1495, n2063}), .b ({new_AGEMA_signal_3520, new_AGEMA_signal_3516}), .clk ( clk ), .r ( Fresh[593] ), .c ({new_AGEMA_signal_1602, n2064}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2229 ( .a ({new_AGEMA_signal_1497, n2076}), .b ({new_AGEMA_signal_3528, new_AGEMA_signal_3524}), .clk ( clk ), .r ( Fresh[594] ), .c ({new_AGEMA_signal_1603, n2077}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2249 ( .a ({new_AGEMA_signal_1501, n2090}), .b ({new_AGEMA_signal_3532, new_AGEMA_signal_3530}), .clk ( clk ), .r ( Fresh[595] ), .c ({new_AGEMA_signal_1604, n2158}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2255 ( .a ({new_AGEMA_signal_1502, n2093}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3534}), .clk ( clk ), .r ( Fresh[596] ), .c ({new_AGEMA_signal_1605, n2095}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2274 ( .a ({new_AGEMA_signal_1606, n2116}), .b ({new_AGEMA_signal_3540, new_AGEMA_signal_3538}), .clk ( clk ), .r ( Fresh[597] ), .c ({new_AGEMA_signal_1681, n2117}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2283 ( .a ({new_AGEMA_signal_3548, new_AGEMA_signal_3544}), .b ({new_AGEMA_signal_1505, n2120}), .clk ( clk ), .r ( Fresh[598] ), .c ({new_AGEMA_signal_1607, n2123}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2300 ( .a ({new_AGEMA_signal_3552, new_AGEMA_signal_3550}), .b ({new_AGEMA_signal_1360, n2134}), .clk ( clk ), .r ( Fresh[599] ), .c ({new_AGEMA_signal_1507, n2135}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2309 ( .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3556}), .b ({new_AGEMA_signal_1509, n2140}), .clk ( clk ), .r ( Fresh[600] ), .c ({new_AGEMA_signal_1609, n2141}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2327 ( .a ({new_AGEMA_signal_3572, new_AGEMA_signal_3566}), .b ({new_AGEMA_signal_1511, n2161}), .clk ( clk ), .r ( Fresh[601] ), .c ({new_AGEMA_signal_1610, n2166}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2331 ( .a ({new_AGEMA_signal_3580, new_AGEMA_signal_3576}), .b ({new_AGEMA_signal_1367, n2164}), .clk ( clk ), .r ( Fresh[602] ), .c ({new_AGEMA_signal_1512, n2165}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2346 ( .a ({new_AGEMA_signal_1513, n2179}), .b ({new_AGEMA_signal_3588, new_AGEMA_signal_3584}), .clk ( clk ), .r ( Fresh[603] ), .c ({new_AGEMA_signal_1611, n2180}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2360 ( .a ({new_AGEMA_signal_3592, new_AGEMA_signal_3590}), .b ({new_AGEMA_signal_1514, n2192}), .clk ( clk ), .r ( Fresh[604] ), .c ({new_AGEMA_signal_1612, n2194}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2372 ( .a ({new_AGEMA_signal_1613, n2203}), .b ({new_AGEMA_signal_3596, new_AGEMA_signal_3594}), .clk ( clk ), .r ( Fresh[605] ), .c ({new_AGEMA_signal_1688, n2204}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2389 ( .a ({new_AGEMA_signal_1517, n2224}), .b ({new_AGEMA_signal_1518, n2223}), .clk ( clk ), .r ( Fresh[606] ), .c ({new_AGEMA_signal_1614, n2225}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2394 ( .a ({new_AGEMA_signal_1379, n2229}), .b ({new_AGEMA_signal_3600, new_AGEMA_signal_3598}), .clk ( clk ), .r ( Fresh[607] ), .c ({new_AGEMA_signal_1519, n2230}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2400 ( .a ({new_AGEMA_signal_3604, new_AGEMA_signal_3602}), .b ({new_AGEMA_signal_1616, n2234}), .clk ( clk ), .r ( Fresh[608] ), .c ({new_AGEMA_signal_1690, n2236}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2412 ( .a ({new_AGEMA_signal_1521, n2246}), .b ({new_AGEMA_signal_3612, new_AGEMA_signal_3608}), .clk ( clk ), .r ( Fresh[609] ), .c ({new_AGEMA_signal_1617, n2247}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2419 ( .a ({new_AGEMA_signal_1522, n2254}), .b ({new_AGEMA_signal_3624, new_AGEMA_signal_3618}), .clk ( clk ), .r ( Fresh[610] ), .c ({new_AGEMA_signal_1618, n2255}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2427 ( .a ({new_AGEMA_signal_1523, n2263}), .b ({new_AGEMA_signal_3632, new_AGEMA_signal_3628}), .clk ( clk ), .r ( Fresh[611] ), .c ({new_AGEMA_signal_1619, n2264}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2435 ( .a ({new_AGEMA_signal_3636, new_AGEMA_signal_3634}), .b ({new_AGEMA_signal_1385, n2267}), .clk ( clk ), .r ( Fresh[612] ), .c ({new_AGEMA_signal_1620, n2271}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2446 ( .a ({new_AGEMA_signal_3468, new_AGEMA_signal_3464}), .b ({new_AGEMA_signal_1387, n2279}), .clk ( clk ), .r ( Fresh[613] ), .c ({new_AGEMA_signal_1526, n2280}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2451 ( .a ({new_AGEMA_signal_3640, new_AGEMA_signal_3638}), .b ({new_AGEMA_signal_1388, n2283}), .clk ( clk ), .r ( Fresh[614] ), .c ({new_AGEMA_signal_1527, n2286}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2461 ( .a ({new_AGEMA_signal_1529, n2686}), .b ({new_AGEMA_signal_1530, n2289}), .clk ( clk ), .r ( Fresh[615] ), .c ({new_AGEMA_signal_1622, n2304}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2466 ( .a ({new_AGEMA_signal_3644, new_AGEMA_signal_3642}), .b ({new_AGEMA_signal_1532, n2292}), .clk ( clk ), .r ( Fresh[616] ), .c ({new_AGEMA_signal_1623, n2295}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2488 ( .a ({new_AGEMA_signal_1534, n2321}), .b ({new_AGEMA_signal_1233, n2320}), .clk ( clk ), .r ( Fresh[617] ), .c ({new_AGEMA_signal_1624, n2322}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2499 ( .a ({new_AGEMA_signal_1535, n2332}), .b ({new_AGEMA_signal_1536, n2331}), .clk ( clk ), .r ( Fresh[618] ), .c ({new_AGEMA_signal_1625, n2333}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2509 ( .a ({new_AGEMA_signal_3652, new_AGEMA_signal_3648}), .b ({new_AGEMA_signal_1538, n2342}), .clk ( clk ), .r ( Fresh[619] ), .c ({new_AGEMA_signal_1627, n2345}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2526 ( .a ({new_AGEMA_signal_1539, n2358}), .b ({new_AGEMA_signal_3656, new_AGEMA_signal_3654}), .clk ( clk ), .r ( Fresh[620] ), .c ({new_AGEMA_signal_1628, n2361}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2549 ( .a ({new_AGEMA_signal_1406, n2387}), .b ({new_AGEMA_signal_3660, new_AGEMA_signal_3658}), .clk ( clk ), .r ( Fresh[621] ), .c ({new_AGEMA_signal_1541, n2388}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2556 ( .a ({new_AGEMA_signal_3668, new_AGEMA_signal_3664}), .b ({new_AGEMA_signal_1542, n2392}), .clk ( clk ), .r ( Fresh[622] ), .c ({new_AGEMA_signal_1630, n2393}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2567 ( .a ({new_AGEMA_signal_3676, new_AGEMA_signal_3672}), .b ({new_AGEMA_signal_1410, n2404}), .clk ( clk ), .r ( Fresh[623] ), .c ({new_AGEMA_signal_1543, n2405}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2571 ( .a ({new_AGEMA_signal_1544, n2409}), .b ({new_AGEMA_signal_3684, new_AGEMA_signal_3680}), .clk ( clk ), .r ( Fresh[624] ), .c ({new_AGEMA_signal_1632, n2410}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2576 ( .a ({new_AGEMA_signal_3692, new_AGEMA_signal_3688}), .b ({new_AGEMA_signal_1545, n2414}), .clk ( clk ), .r ( Fresh[625] ), .c ({new_AGEMA_signal_1633, n2421}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2579 ( .a ({new_AGEMA_signal_1413, n2418}), .b ({new_AGEMA_signal_3700, new_AGEMA_signal_3696}), .clk ( clk ), .r ( Fresh[626] ), .c ({new_AGEMA_signal_1546, n2419}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2590 ( .a ({new_AGEMA_signal_3704, new_AGEMA_signal_3702}), .b ({new_AGEMA_signal_1547, n2432}), .clk ( clk ), .r ( Fresh[627] ), .c ({new_AGEMA_signal_1635, n2436}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2604 ( .a ({new_AGEMA_signal_1548, n2449}), .b ({new_AGEMA_signal_1549, n2448}), .clk ( clk ), .r ( Fresh[628] ), .c ({new_AGEMA_signal_1636, n2450}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2610 ( .a ({new_AGEMA_signal_3708, new_AGEMA_signal_3706}), .b ({new_AGEMA_signal_1550, n2455}), .clk ( clk ), .r ( Fresh[629] ), .c ({new_AGEMA_signal_1637, n2456}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2613 ( .a ({new_AGEMA_signal_1551, n2460}), .b ({new_AGEMA_signal_3712, new_AGEMA_signal_3710}), .clk ( clk ), .r ( Fresh[630] ), .c ({new_AGEMA_signal_1638, n2461}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2619 ( .a ({new_AGEMA_signal_3716, new_AGEMA_signal_3714}), .b ({new_AGEMA_signal_1422, n2466}), .clk ( clk ), .r ( Fresh[631] ), .c ({new_AGEMA_signal_1552, n2469}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2630 ( .a ({new_AGEMA_signal_3724, new_AGEMA_signal_3720}), .b ({new_AGEMA_signal_1423, n2477}), .clk ( clk ), .r ( Fresh[632] ), .c ({new_AGEMA_signal_1553, n2478}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2635 ( .a ({new_AGEMA_signal_3732, new_AGEMA_signal_3728}), .b ({new_AGEMA_signal_1554, n2482}), .clk ( clk ), .r ( Fresh[633] ), .c ({new_AGEMA_signal_1640, n2484}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2643 ( .a ({new_AGEMA_signal_1425, n2490}), .b ({new_AGEMA_signal_3736, new_AGEMA_signal_3734}), .clk ( clk ), .r ( Fresh[634] ), .c ({new_AGEMA_signal_1555, n2491}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2649 ( .a ({new_AGEMA_signal_3740, new_AGEMA_signal_3738}), .b ({new_AGEMA_signal_1556, n2496}), .clk ( clk ), .r ( Fresh[635] ), .c ({new_AGEMA_signal_1642, n2500}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2656 ( .a ({new_AGEMA_signal_1643, n2507}), .b ({new_AGEMA_signal_3744, new_AGEMA_signal_3742}), .clk ( clk ), .r ( Fresh[636] ), .c ({new_AGEMA_signal_1708, n2508}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2670 ( .a ({new_AGEMA_signal_1644, n2525}), .b ({new_AGEMA_signal_1559, n2524}), .clk ( clk ), .r ( Fresh[637] ), .c ({new_AGEMA_signal_1709, n2526}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2679 ( .a ({new_AGEMA_signal_1560, n2537}), .b ({new_AGEMA_signal_1561, n2536}), .clk ( clk ), .r ( Fresh[638] ), .c ({new_AGEMA_signal_1645, n2539}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2682 ( .a ({new_AGEMA_signal_1506, n2543}), .b ({new_AGEMA_signal_3748, new_AGEMA_signal_3746}), .clk ( clk ), .r ( Fresh[639] ), .c ({new_AGEMA_signal_1646, n2548}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2694 ( .a ({new_AGEMA_signal_3752, new_AGEMA_signal_3750}), .b ({new_AGEMA_signal_1562, n2557}), .clk ( clk ), .r ( Fresh[640] ), .c ({new_AGEMA_signal_1647, n2568}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2700 ( .a ({new_AGEMA_signal_3756, new_AGEMA_signal_3754}), .b ({new_AGEMA_signal_1563, n2565}), .clk ( clk ), .r ( Fresh[641] ), .c ({new_AGEMA_signal_1648, n2567}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2710 ( .a ({new_AGEMA_signal_3760, new_AGEMA_signal_3758}), .b ({new_AGEMA_signal_1565, n2580}), .clk ( clk ), .r ( Fresh[642] ), .c ({new_AGEMA_signal_1649, n2583}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2728 ( .a ({new_AGEMA_signal_3764, new_AGEMA_signal_3762}), .b ({new_AGEMA_signal_1282, n2602}), .clk ( clk ), .r ( Fresh[643] ), .c ({new_AGEMA_signal_1566, n2604}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2739 ( .a ({new_AGEMA_signal_3768, new_AGEMA_signal_3766}), .b ({new_AGEMA_signal_1567, n2619}), .clk ( clk ), .r ( Fresh[644] ), .c ({new_AGEMA_signal_1651, n2621}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2745 ( .a ({new_AGEMA_signal_3776, new_AGEMA_signal_3772}), .b ({new_AGEMA_signal_1568, n2628}), .clk ( clk ), .r ( Fresh[645] ), .c ({new_AGEMA_signal_1652, n2633}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2756 ( .a ({new_AGEMA_signal_1569, n2649}), .b ({new_AGEMA_signal_1451, n2648}), .clk ( clk ), .r ( Fresh[646] ), .c ({new_AGEMA_signal_1653, n2660}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2759 ( .a ({new_AGEMA_signal_3780, new_AGEMA_signal_3778}), .b ({new_AGEMA_signal_1496, n2652}), .clk ( clk ), .r ( Fresh[647] ), .c ({new_AGEMA_signal_1654, n2656}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2766 ( .a ({new_AGEMA_signal_3784, new_AGEMA_signal_3782}), .b ({new_AGEMA_signal_1570, n2664}), .clk ( clk ), .r ( Fresh[648] ), .c ({new_AGEMA_signal_1655, n2666}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2774 ( .a ({new_AGEMA_signal_1571, n2681}), .b ({new_AGEMA_signal_1454, n2680}), .clk ( clk ), .r ( Fresh[649] ), .c ({new_AGEMA_signal_1656, n2706}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2777 ( .a ({new_AGEMA_signal_1529, n2686}), .b ({new_AGEMA_signal_1572, n2685}), .clk ( clk ), .r ( Fresh[650] ), .c ({new_AGEMA_signal_1657, n2704}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2781 ( .a ({new_AGEMA_signal_1574, n2692}), .b ({new_AGEMA_signal_3788, new_AGEMA_signal_3786}), .clk ( clk ), .r ( Fresh[651] ), .c ({new_AGEMA_signal_1658, n2696}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2794 ( .a ({new_AGEMA_signal_3792, new_AGEMA_signal_3790}), .b ({new_AGEMA_signal_1575, n2716}), .clk ( clk ), .r ( Fresh[652] ), .c ({new_AGEMA_signal_1659, n2718}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2801 ( .a ({new_AGEMA_signal_3796, new_AGEMA_signal_3794}), .b ({new_AGEMA_signal_1457, n2728}), .clk ( clk ), .r ( Fresh[653] ), .c ({new_AGEMA_signal_1660, n2730}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2805 ( .a ({new_AGEMA_signal_3804, new_AGEMA_signal_3800}), .b ({new_AGEMA_signal_1577, n2735}), .clk ( clk ), .r ( Fresh[654] ), .c ({new_AGEMA_signal_1661, n2745}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2809 ( .a ({new_AGEMA_signal_1578, n2743}), .b ({new_AGEMA_signal_3812, new_AGEMA_signal_3808}), .clk ( clk ), .r ( Fresh[655] ), .c ({new_AGEMA_signal_1662, n2744}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2814 ( .a ({new_AGEMA_signal_3636, new_AGEMA_signal_3634}), .b ({new_AGEMA_signal_1460, n2751}), .clk ( clk ), .r ( Fresh[656] ), .c ({new_AGEMA_signal_1663, n2759}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2821 ( .a ({new_AGEMA_signal_3820, new_AGEMA_signal_3816}), .b ({new_AGEMA_signal_1580, n2764}), .clk ( clk ), .r ( Fresh[657] ), .c ({new_AGEMA_signal_1664, n2771}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2833 ( .a ({new_AGEMA_signal_1466, n2788}), .b ({new_AGEMA_signal_3828, new_AGEMA_signal_3824}), .clk ( clk ), .r ( Fresh[658] ), .c ({new_AGEMA_signal_1582, n2798}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2850 ( .a ({new_AGEMA_signal_1584, n2822}), .b ({new_AGEMA_signal_1469, n2821}), .clk ( clk ), .r ( Fresh[659] ), .c ({new_AGEMA_signal_1666, n2826}) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C ( clk ), .D ( new_AGEMA_signal_3831 ), .Q ( new_AGEMA_signal_3832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C ( clk ), .D ( new_AGEMA_signal_3835 ), .Q ( new_AGEMA_signal_3836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C ( clk ), .D ( new_AGEMA_signal_3839 ), .Q ( new_AGEMA_signal_3840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C ( clk ), .D ( new_AGEMA_signal_3843 ), .Q ( new_AGEMA_signal_3844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C ( clk ), .D ( new_AGEMA_signal_3851 ), .Q ( new_AGEMA_signal_3852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C ( clk ), .D ( new_AGEMA_signal_3859 ), .Q ( new_AGEMA_signal_3860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C ( clk ), .D ( new_AGEMA_signal_3861 ), .Q ( new_AGEMA_signal_3862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C ( clk ), .D ( new_AGEMA_signal_3863 ), .Q ( new_AGEMA_signal_3864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C ( clk ), .D ( new_AGEMA_signal_3871 ), .Q ( new_AGEMA_signal_3872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C ( clk ), .D ( new_AGEMA_signal_3879 ), .Q ( new_AGEMA_signal_3880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C ( clk ), .D ( new_AGEMA_signal_3885 ), .Q ( new_AGEMA_signal_3886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C ( clk ), .D ( new_AGEMA_signal_3891 ), .Q ( new_AGEMA_signal_3892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C ( clk ), .D ( new_AGEMA_signal_3895 ), .Q ( new_AGEMA_signal_3896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C ( clk ), .D ( new_AGEMA_signal_3899 ), .Q ( new_AGEMA_signal_3900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C ( clk ), .D ( new_AGEMA_signal_3905 ), .Q ( new_AGEMA_signal_3906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C ( clk ), .D ( new_AGEMA_signal_3911 ), .Q ( new_AGEMA_signal_3912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C ( clk ), .D ( new_AGEMA_signal_3913 ), .Q ( new_AGEMA_signal_3914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C ( clk ), .D ( new_AGEMA_signal_3915 ), .Q ( new_AGEMA_signal_3916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C ( clk ), .D ( new_AGEMA_signal_3921 ), .Q ( new_AGEMA_signal_3922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C ( clk ), .D ( new_AGEMA_signal_3927 ), .Q ( new_AGEMA_signal_3928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C ( clk ), .D ( new_AGEMA_signal_3933 ), .Q ( new_AGEMA_signal_3934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C ( clk ), .D ( new_AGEMA_signal_3939 ), .Q ( new_AGEMA_signal_3940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C ( clk ), .D ( new_AGEMA_signal_3941 ), .Q ( new_AGEMA_signal_3942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C ( clk ), .D ( new_AGEMA_signal_3943 ), .Q ( new_AGEMA_signal_3944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C ( clk ), .D ( new_AGEMA_signal_3947 ), .Q ( new_AGEMA_signal_3948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C ( clk ), .D ( new_AGEMA_signal_3951 ), .Q ( new_AGEMA_signal_3952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C ( clk ), .D ( new_AGEMA_signal_3957 ), .Q ( new_AGEMA_signal_3958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C ( clk ), .D ( new_AGEMA_signal_3963 ), .Q ( new_AGEMA_signal_3964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C ( clk ), .D ( new_AGEMA_signal_3969 ), .Q ( new_AGEMA_signal_3970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C ( clk ), .D ( new_AGEMA_signal_3975 ), .Q ( new_AGEMA_signal_3976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C ( clk ), .D ( new_AGEMA_signal_3977 ), .Q ( new_AGEMA_signal_3978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C ( clk ), .D ( new_AGEMA_signal_3979 ), .Q ( new_AGEMA_signal_3980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C ( clk ), .D ( new_AGEMA_signal_3985 ), .Q ( new_AGEMA_signal_3986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C ( clk ), .D ( new_AGEMA_signal_3991 ), .Q ( new_AGEMA_signal_3992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C ( clk ), .D ( new_AGEMA_signal_3993 ), .Q ( new_AGEMA_signal_3994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C ( clk ), .D ( new_AGEMA_signal_3995 ), .Q ( new_AGEMA_signal_3996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C ( clk ), .D ( new_AGEMA_signal_3999 ), .Q ( new_AGEMA_signal_4000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C ( clk ), .D ( new_AGEMA_signal_4003 ), .Q ( new_AGEMA_signal_4004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C ( clk ), .D ( new_AGEMA_signal_4007 ), .Q ( new_AGEMA_signal_4008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C ( clk ), .D ( new_AGEMA_signal_4011 ), .Q ( new_AGEMA_signal_4012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C ( clk ), .D ( new_AGEMA_signal_4013 ), .Q ( new_AGEMA_signal_4014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C ( clk ), .D ( new_AGEMA_signal_4015 ), .Q ( new_AGEMA_signal_4016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C ( clk ), .D ( new_AGEMA_signal_4023 ), .Q ( new_AGEMA_signal_4024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C ( clk ), .D ( new_AGEMA_signal_4031 ), .Q ( new_AGEMA_signal_4032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C ( clk ), .D ( new_AGEMA_signal_4037 ), .Q ( new_AGEMA_signal_4038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C ( clk ), .D ( new_AGEMA_signal_4043 ), .Q ( new_AGEMA_signal_4044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C ( clk ), .D ( new_AGEMA_signal_4047 ), .Q ( new_AGEMA_signal_4048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C ( clk ), .D ( new_AGEMA_signal_4051 ), .Q ( new_AGEMA_signal_4052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C ( clk ), .D ( new_AGEMA_signal_4055 ), .Q ( new_AGEMA_signal_4056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C ( clk ), .D ( new_AGEMA_signal_4059 ), .Q ( new_AGEMA_signal_4060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C ( clk ), .D ( new_AGEMA_signal_4061 ), .Q ( new_AGEMA_signal_4062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C ( clk ), .D ( new_AGEMA_signal_4063 ), .Q ( new_AGEMA_signal_4064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C ( clk ), .D ( new_AGEMA_signal_4065 ), .Q ( new_AGEMA_signal_4066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C ( clk ), .D ( new_AGEMA_signal_4067 ), .Q ( new_AGEMA_signal_4068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C ( clk ), .D ( new_AGEMA_signal_4071 ), .Q ( new_AGEMA_signal_4072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C ( clk ), .D ( new_AGEMA_signal_4075 ), .Q ( new_AGEMA_signal_4076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C ( clk ), .D ( new_AGEMA_signal_4079 ), .Q ( new_AGEMA_signal_4080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C ( clk ), .D ( new_AGEMA_signal_4083 ), .Q ( new_AGEMA_signal_4084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C ( clk ), .D ( new_AGEMA_signal_4085 ), .Q ( new_AGEMA_signal_4086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C ( clk ), .D ( new_AGEMA_signal_4087 ), .Q ( new_AGEMA_signal_4088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C ( clk ), .D ( new_AGEMA_signal_4093 ), .Q ( new_AGEMA_signal_4094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C ( clk ), .D ( new_AGEMA_signal_4099 ), .Q ( new_AGEMA_signal_4100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C ( clk ), .D ( new_AGEMA_signal_4103 ), .Q ( new_AGEMA_signal_4104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C ( clk ), .D ( new_AGEMA_signal_4107 ), .Q ( new_AGEMA_signal_4108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C ( clk ), .D ( new_AGEMA_signal_4109 ), .Q ( new_AGEMA_signal_4110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C ( clk ), .D ( new_AGEMA_signal_4111 ), .Q ( new_AGEMA_signal_4112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C ( clk ), .D ( new_AGEMA_signal_4115 ), .Q ( new_AGEMA_signal_4116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C ( clk ), .D ( new_AGEMA_signal_4119 ), .Q ( new_AGEMA_signal_4120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C ( clk ), .D ( new_AGEMA_signal_4123 ), .Q ( new_AGEMA_signal_4124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C ( clk ), .D ( new_AGEMA_signal_4127 ), .Q ( new_AGEMA_signal_4128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C ( clk ), .D ( new_AGEMA_signal_4131 ), .Q ( new_AGEMA_signal_4132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C ( clk ), .D ( new_AGEMA_signal_4135 ), .Q ( new_AGEMA_signal_4136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C ( clk ), .D ( new_AGEMA_signal_4137 ), .Q ( new_AGEMA_signal_4138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C ( clk ), .D ( new_AGEMA_signal_4139 ), .Q ( new_AGEMA_signal_4140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C ( clk ), .D ( new_AGEMA_signal_4143 ), .Q ( new_AGEMA_signal_4144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C ( clk ), .D ( new_AGEMA_signal_4147 ), .Q ( new_AGEMA_signal_4148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C ( clk ), .D ( new_AGEMA_signal_4149 ), .Q ( new_AGEMA_signal_4150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C ( clk ), .D ( new_AGEMA_signal_4151 ), .Q ( new_AGEMA_signal_4152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C ( clk ), .D ( new_AGEMA_signal_4157 ), .Q ( new_AGEMA_signal_4158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C ( clk ), .D ( new_AGEMA_signal_4163 ), .Q ( new_AGEMA_signal_4164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C ( clk ), .D ( new_AGEMA_signal_4169 ), .Q ( new_AGEMA_signal_4170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C ( clk ), .D ( new_AGEMA_signal_4175 ), .Q ( new_AGEMA_signal_4176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C ( clk ), .D ( new_AGEMA_signal_4179 ), .Q ( new_AGEMA_signal_4180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C ( clk ), .D ( new_AGEMA_signal_4183 ), .Q ( new_AGEMA_signal_4184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C ( clk ), .D ( new_AGEMA_signal_4185 ), .Q ( new_AGEMA_signal_4186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C ( clk ), .D ( new_AGEMA_signal_4187 ), .Q ( new_AGEMA_signal_4188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C ( clk ), .D ( new_AGEMA_signal_4195 ), .Q ( new_AGEMA_signal_4196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C ( clk ), .D ( new_AGEMA_signal_4203 ), .Q ( new_AGEMA_signal_4204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C ( clk ), .D ( new_AGEMA_signal_4205 ), .Q ( new_AGEMA_signal_4206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C ( clk ), .D ( new_AGEMA_signal_4207 ), .Q ( new_AGEMA_signal_4208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C ( clk ), .D ( new_AGEMA_signal_4211 ), .Q ( new_AGEMA_signal_4212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C ( clk ), .D ( new_AGEMA_signal_4215 ), .Q ( new_AGEMA_signal_4216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C ( clk ), .D ( new_AGEMA_signal_4219 ), .Q ( new_AGEMA_signal_4220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C ( clk ), .D ( new_AGEMA_signal_4223 ), .Q ( new_AGEMA_signal_4224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C ( clk ), .D ( new_AGEMA_signal_4227 ), .Q ( new_AGEMA_signal_4228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C ( clk ), .D ( new_AGEMA_signal_4231 ), .Q ( new_AGEMA_signal_4232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C ( clk ), .D ( new_AGEMA_signal_4235 ), .Q ( new_AGEMA_signal_4236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C ( clk ), .D ( new_AGEMA_signal_4239 ), .Q ( new_AGEMA_signal_4240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C ( clk ), .D ( new_AGEMA_signal_4243 ), .Q ( new_AGEMA_signal_4244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C ( clk ), .D ( new_AGEMA_signal_4247 ), .Q ( new_AGEMA_signal_4248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C ( clk ), .D ( new_AGEMA_signal_4255 ), .Q ( new_AGEMA_signal_4256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C ( clk ), .D ( new_AGEMA_signal_4263 ), .Q ( new_AGEMA_signal_4264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C ( clk ), .D ( new_AGEMA_signal_4265 ), .Q ( new_AGEMA_signal_4266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C ( clk ), .D ( new_AGEMA_signal_4267 ), .Q ( new_AGEMA_signal_4268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C ( clk ), .D ( new_AGEMA_signal_4271 ), .Q ( new_AGEMA_signal_4272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C ( clk ), .D ( new_AGEMA_signal_4275 ), .Q ( new_AGEMA_signal_4276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C ( clk ), .D ( new_AGEMA_signal_4277 ), .Q ( new_AGEMA_signal_4278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C ( clk ), .D ( new_AGEMA_signal_4279 ), .Q ( new_AGEMA_signal_4280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C ( clk ), .D ( new_AGEMA_signal_4285 ), .Q ( new_AGEMA_signal_4286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C ( clk ), .D ( new_AGEMA_signal_4291 ), .Q ( new_AGEMA_signal_4292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C ( clk ), .D ( new_AGEMA_signal_4301 ), .Q ( new_AGEMA_signal_4302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C ( clk ), .D ( new_AGEMA_signal_4309 ), .Q ( new_AGEMA_signal_4310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C ( clk ), .D ( new_AGEMA_signal_4317 ), .Q ( new_AGEMA_signal_4318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C ( clk ), .D ( new_AGEMA_signal_4321 ), .Q ( new_AGEMA_signal_4322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C ( clk ), .D ( new_AGEMA_signal_4329 ), .Q ( new_AGEMA_signal_4330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C ( clk ), .D ( new_AGEMA_signal_4337 ), .Q ( new_AGEMA_signal_4338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C ( clk ), .D ( new_AGEMA_signal_4347 ), .Q ( new_AGEMA_signal_4348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C ( clk ), .D ( new_AGEMA_signal_4353 ), .Q ( new_AGEMA_signal_4354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C ( clk ), .D ( new_AGEMA_signal_4357 ), .Q ( new_AGEMA_signal_4358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C ( clk ), .D ( new_AGEMA_signal_4361 ), .Q ( new_AGEMA_signal_4362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C ( clk ), .D ( new_AGEMA_signal_4369 ), .Q ( new_AGEMA_signal_4370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C ( clk ), .D ( new_AGEMA_signal_4377 ), .Q ( new_AGEMA_signal_4378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C ( clk ), .D ( new_AGEMA_signal_4381 ), .Q ( new_AGEMA_signal_4382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C ( clk ), .D ( new_AGEMA_signal_4385 ), .Q ( new_AGEMA_signal_4386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C ( clk ), .D ( new_AGEMA_signal_4391 ), .Q ( new_AGEMA_signal_4392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C ( clk ), .D ( new_AGEMA_signal_4397 ), .Q ( new_AGEMA_signal_4398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C ( clk ), .D ( new_AGEMA_signal_4403 ), .Q ( new_AGEMA_signal_4404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C ( clk ), .D ( new_AGEMA_signal_4409 ), .Q ( new_AGEMA_signal_4410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C ( clk ), .D ( new_AGEMA_signal_4415 ), .Q ( new_AGEMA_signal_4416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C ( clk ), .D ( new_AGEMA_signal_4421 ), .Q ( new_AGEMA_signal_4422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C ( clk ), .D ( new_AGEMA_signal_4427 ), .Q ( new_AGEMA_signal_4428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C ( clk ), .D ( new_AGEMA_signal_4433 ), .Q ( new_AGEMA_signal_4434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C ( clk ), .D ( new_AGEMA_signal_4439 ), .Q ( new_AGEMA_signal_4440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C ( clk ), .D ( new_AGEMA_signal_4445 ), .Q ( new_AGEMA_signal_4446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C ( clk ), .D ( new_AGEMA_signal_4449 ), .Q ( new_AGEMA_signal_4450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C ( clk ), .D ( new_AGEMA_signal_4453 ), .Q ( new_AGEMA_signal_4454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C ( clk ), .D ( new_AGEMA_signal_4461 ), .Q ( new_AGEMA_signal_4462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C ( clk ), .D ( new_AGEMA_signal_4469 ), .Q ( new_AGEMA_signal_4470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C ( clk ), .D ( new_AGEMA_signal_4473 ), .Q ( new_AGEMA_signal_4474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C ( clk ), .D ( new_AGEMA_signal_4477 ), .Q ( new_AGEMA_signal_4478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C ( clk ), .D ( new_AGEMA_signal_4483 ), .Q ( new_AGEMA_signal_4484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C ( clk ), .D ( new_AGEMA_signal_4489 ), .Q ( new_AGEMA_signal_4490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C ( clk ), .D ( new_AGEMA_signal_4497 ), .Q ( new_AGEMA_signal_4498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C ( clk ), .D ( new_AGEMA_signal_4505 ), .Q ( new_AGEMA_signal_4506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C ( clk ), .D ( new_AGEMA_signal_4515 ), .Q ( new_AGEMA_signal_4516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C ( clk ), .D ( new_AGEMA_signal_4521 ), .Q ( new_AGEMA_signal_4522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C ( clk ), .D ( new_AGEMA_signal_4535 ), .Q ( new_AGEMA_signal_4536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C ( clk ), .D ( new_AGEMA_signal_4541 ), .Q ( new_AGEMA_signal_4542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C ( clk ), .D ( new_AGEMA_signal_4547 ), .Q ( new_AGEMA_signal_4548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C ( clk ), .D ( new_AGEMA_signal_4553 ), .Q ( new_AGEMA_signal_4554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C ( clk ), .D ( new_AGEMA_signal_4561 ), .Q ( new_AGEMA_signal_4562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C ( clk ), .D ( new_AGEMA_signal_4569 ), .Q ( new_AGEMA_signal_4570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C ( clk ), .D ( new_AGEMA_signal_4577 ), .Q ( new_AGEMA_signal_4578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C ( clk ), .D ( new_AGEMA_signal_4585 ), .Q ( new_AGEMA_signal_4586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C ( clk ), .D ( new_AGEMA_signal_4591 ), .Q ( new_AGEMA_signal_4592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C ( clk ), .D ( new_AGEMA_signal_4597 ), .Q ( new_AGEMA_signal_4598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C ( clk ), .D ( new_AGEMA_signal_4603 ), .Q ( new_AGEMA_signal_4604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C ( clk ), .D ( new_AGEMA_signal_4609 ), .Q ( new_AGEMA_signal_4610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C ( clk ), .D ( new_AGEMA_signal_4617 ), .Q ( new_AGEMA_signal_4618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C ( clk ), .D ( new_AGEMA_signal_4621 ), .Q ( new_AGEMA_signal_4622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C ( clk ), .D ( new_AGEMA_signal_4625 ), .Q ( new_AGEMA_signal_4626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C ( clk ), .D ( new_AGEMA_signal_4629 ), .Q ( new_AGEMA_signal_4630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C ( clk ), .D ( new_AGEMA_signal_4633 ), .Q ( new_AGEMA_signal_4634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C ( clk ), .D ( new_AGEMA_signal_4637 ), .Q ( new_AGEMA_signal_4638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C ( clk ), .D ( new_AGEMA_signal_4645 ), .Q ( new_AGEMA_signal_4646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C ( clk ), .D ( new_AGEMA_signal_4651 ), .Q ( new_AGEMA_signal_4652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C ( clk ), .D ( new_AGEMA_signal_4671 ), .Q ( new_AGEMA_signal_4672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C ( clk ), .D ( new_AGEMA_signal_4679 ), .Q ( new_AGEMA_signal_4680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C ( clk ), .D ( new_AGEMA_signal_4687 ), .Q ( new_AGEMA_signal_4688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C ( clk ), .D ( new_AGEMA_signal_4695 ), .Q ( new_AGEMA_signal_4696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C ( clk ), .D ( new_AGEMA_signal_4703 ), .Q ( new_AGEMA_signal_4704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C ( clk ), .D ( new_AGEMA_signal_4711 ), .Q ( new_AGEMA_signal_4712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C ( clk ), .D ( new_AGEMA_signal_4719 ), .Q ( new_AGEMA_signal_4720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C ( clk ), .D ( new_AGEMA_signal_4727 ), .Q ( new_AGEMA_signal_4728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C ( clk ), .D ( new_AGEMA_signal_4733 ), .Q ( new_AGEMA_signal_4734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C ( clk ), .D ( new_AGEMA_signal_4739 ), .Q ( new_AGEMA_signal_4740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C ( clk ), .D ( new_AGEMA_signal_4749 ), .Q ( new_AGEMA_signal_4750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C ( clk ), .D ( new_AGEMA_signal_4759 ), .Q ( new_AGEMA_signal_4760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C ( clk ), .D ( new_AGEMA_signal_4767 ), .Q ( new_AGEMA_signal_4768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C ( clk ), .D ( new_AGEMA_signal_4775 ), .Q ( new_AGEMA_signal_4776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C ( clk ), .D ( new_AGEMA_signal_4783 ), .Q ( new_AGEMA_signal_4784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C ( clk ), .D ( new_AGEMA_signal_4791 ), .Q ( new_AGEMA_signal_4792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C ( clk ), .D ( new_AGEMA_signal_4799 ), .Q ( new_AGEMA_signal_4800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C ( clk ), .D ( new_AGEMA_signal_4807 ), .Q ( new_AGEMA_signal_4808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C ( clk ), .D ( new_AGEMA_signal_4825 ), .Q ( new_AGEMA_signal_4826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C ( clk ), .D ( new_AGEMA_signal_4831 ), .Q ( new_AGEMA_signal_4832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C ( clk ), .D ( new_AGEMA_signal_4849 ), .Q ( new_AGEMA_signal_4850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C ( clk ), .D ( new_AGEMA_signal_4859 ), .Q ( new_AGEMA_signal_4860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C ( clk ), .D ( new_AGEMA_signal_4867 ), .Q ( new_AGEMA_signal_4868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C ( clk ), .D ( new_AGEMA_signal_4875 ), .Q ( new_AGEMA_signal_4876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C ( clk ), .D ( new_AGEMA_signal_4895 ), .Q ( new_AGEMA_signal_4896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C ( clk ), .D ( new_AGEMA_signal_4903 ), .Q ( new_AGEMA_signal_4904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C ( clk ), .D ( new_AGEMA_signal_4911 ), .Q ( new_AGEMA_signal_4912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C ( clk ), .D ( new_AGEMA_signal_4919 ), .Q ( new_AGEMA_signal_4920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C ( clk ), .D ( new_AGEMA_signal_4925 ), .Q ( new_AGEMA_signal_4926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C ( clk ), .D ( new_AGEMA_signal_4931 ), .Q ( new_AGEMA_signal_4932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C ( clk ), .D ( new_AGEMA_signal_4947 ), .Q ( new_AGEMA_signal_4948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C ( clk ), .D ( new_AGEMA_signal_4955 ), .Q ( new_AGEMA_signal_4956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C ( clk ), .D ( new_AGEMA_signal_5009 ), .Q ( new_AGEMA_signal_5010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C ( clk ), .D ( new_AGEMA_signal_5017 ), .Q ( new_AGEMA_signal_5018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C ( clk ), .D ( new_AGEMA_signal_5045 ), .Q ( new_AGEMA_signal_5046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C ( clk ), .D ( new_AGEMA_signal_5053 ), .Q ( new_AGEMA_signal_5054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C ( clk ), .D ( new_AGEMA_signal_5061 ), .Q ( new_AGEMA_signal_5062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C ( clk ), .D ( new_AGEMA_signal_5069 ), .Q ( new_AGEMA_signal_5070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C ( clk ), .D ( new_AGEMA_signal_5079 ), .Q ( new_AGEMA_signal_5080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C ( clk ), .D ( new_AGEMA_signal_5089 ), .Q ( new_AGEMA_signal_5090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C ( clk ), .D ( new_AGEMA_signal_5097 ), .Q ( new_AGEMA_signal_5098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C ( clk ), .D ( new_AGEMA_signal_5105 ), .Q ( new_AGEMA_signal_5106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C ( clk ), .D ( new_AGEMA_signal_5145 ), .Q ( new_AGEMA_signal_5146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C ( clk ), .D ( new_AGEMA_signal_5153 ), .Q ( new_AGEMA_signal_5154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C ( clk ), .D ( new_AGEMA_signal_5177 ), .Q ( new_AGEMA_signal_5178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C ( clk ), .D ( new_AGEMA_signal_5185 ), .Q ( new_AGEMA_signal_5186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C ( clk ), .D ( new_AGEMA_signal_5265 ), .Q ( new_AGEMA_signal_5266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C ( clk ), .D ( new_AGEMA_signal_5275 ), .Q ( new_AGEMA_signal_5276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C ( clk ), .D ( new_AGEMA_signal_5445 ), .Q ( new_AGEMA_signal_5446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C ( clk ), .D ( new_AGEMA_signal_5457 ), .Q ( new_AGEMA_signal_5458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C ( clk ), .D ( new_AGEMA_signal_5471 ), .Q ( new_AGEMA_signal_5472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C ( clk ), .D ( new_AGEMA_signal_5485 ), .Q ( new_AGEMA_signal_5486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C ( clk ), .D ( new_AGEMA_signal_5515 ), .Q ( new_AGEMA_signal_5516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C ( clk ), .D ( new_AGEMA_signal_5529 ), .Q ( new_AGEMA_signal_5530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C ( clk ), .D ( new_AGEMA_signal_5587 ), .Q ( new_AGEMA_signal_5588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C ( clk ), .D ( new_AGEMA_signal_5603 ), .Q ( new_AGEMA_signal_5604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C ( clk ), .D ( new_AGEMA_signal_5631 ), .Q ( new_AGEMA_signal_5632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C ( clk ), .D ( new_AGEMA_signal_5647 ), .Q ( new_AGEMA_signal_5648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C ( clk ), .D ( new_AGEMA_signal_5729 ), .Q ( new_AGEMA_signal_5730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C ( clk ), .D ( new_AGEMA_signal_5745 ), .Q ( new_AGEMA_signal_5746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C ( clk ), .D ( new_AGEMA_signal_5783 ), .Q ( new_AGEMA_signal_5784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C ( clk ), .D ( new_AGEMA_signal_5801 ), .Q ( new_AGEMA_signal_5802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C ( clk ), .D ( new_AGEMA_signal_5883 ), .Q ( new_AGEMA_signal_5884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C ( clk ), .D ( new_AGEMA_signal_5903 ), .Q ( new_AGEMA_signal_5904 ) ) ;

    /* cells in depth 11 */
    buf_clk new_AGEMA_reg_buffer_2475 ( .C ( clk ), .D ( n1934 ), .Q ( new_AGEMA_signal_4293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C ( clk ), .D ( new_AGEMA_signal_1585 ), .Q ( new_AGEMA_signal_4295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C ( clk ), .D ( new_AGEMA_signal_4302 ), .Q ( new_AGEMA_signal_4303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C ( clk ), .D ( new_AGEMA_signal_4310 ), .Q ( new_AGEMA_signal_4311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C ( clk ), .D ( n1981 ), .Q ( new_AGEMA_signal_4313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C ( clk ), .D ( new_AGEMA_signal_1593 ), .Q ( new_AGEMA_signal_4315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C ( clk ), .D ( new_AGEMA_signal_4318 ), .Q ( new_AGEMA_signal_4319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C ( clk ), .D ( new_AGEMA_signal_4322 ), .Q ( new_AGEMA_signal_4323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C ( clk ), .D ( new_AGEMA_signal_4330 ), .Q ( new_AGEMA_signal_4331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C ( clk ), .D ( new_AGEMA_signal_4338 ), .Q ( new_AGEMA_signal_4339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C ( clk ), .D ( new_AGEMA_signal_3872 ), .Q ( new_AGEMA_signal_4341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C ( clk ), .D ( new_AGEMA_signal_3880 ), .Q ( new_AGEMA_signal_4343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C ( clk ), .D ( new_AGEMA_signal_4348 ), .Q ( new_AGEMA_signal_4349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C ( clk ), .D ( new_AGEMA_signal_4354 ), .Q ( new_AGEMA_signal_4355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C ( clk ), .D ( new_AGEMA_signal_4358 ), .Q ( new_AGEMA_signal_4359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C ( clk ), .D ( new_AGEMA_signal_4362 ), .Q ( new_AGEMA_signal_4363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C ( clk ), .D ( new_AGEMA_signal_4370 ), .Q ( new_AGEMA_signal_4371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C ( clk ), .D ( new_AGEMA_signal_4378 ), .Q ( new_AGEMA_signal_4379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C ( clk ), .D ( new_AGEMA_signal_4382 ), .Q ( new_AGEMA_signal_4383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C ( clk ), .D ( new_AGEMA_signal_4386 ), .Q ( new_AGEMA_signal_4387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C ( clk ), .D ( new_AGEMA_signal_4392 ), .Q ( new_AGEMA_signal_4393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C ( clk ), .D ( new_AGEMA_signal_4398 ), .Q ( new_AGEMA_signal_4399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C ( clk ), .D ( new_AGEMA_signal_4404 ), .Q ( new_AGEMA_signal_4405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C ( clk ), .D ( new_AGEMA_signal_4410 ), .Q ( new_AGEMA_signal_4411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C ( clk ), .D ( new_AGEMA_signal_4416 ), .Q ( new_AGEMA_signal_4417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C ( clk ), .D ( new_AGEMA_signal_4422 ), .Q ( new_AGEMA_signal_4423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C ( clk ), .D ( new_AGEMA_signal_4428 ), .Q ( new_AGEMA_signal_4429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C ( clk ), .D ( new_AGEMA_signal_4434 ), .Q ( new_AGEMA_signal_4435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C ( clk ), .D ( new_AGEMA_signal_4440 ), .Q ( new_AGEMA_signal_4441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C ( clk ), .D ( new_AGEMA_signal_4446 ), .Q ( new_AGEMA_signal_4447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C ( clk ), .D ( new_AGEMA_signal_4450 ), .Q ( new_AGEMA_signal_4451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C ( clk ), .D ( new_AGEMA_signal_4454 ), .Q ( new_AGEMA_signal_4455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C ( clk ), .D ( new_AGEMA_signal_4462 ), .Q ( new_AGEMA_signal_4463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C ( clk ), .D ( new_AGEMA_signal_4470 ), .Q ( new_AGEMA_signal_4471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C ( clk ), .D ( new_AGEMA_signal_4474 ), .Q ( new_AGEMA_signal_4475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C ( clk ), .D ( new_AGEMA_signal_4478 ), .Q ( new_AGEMA_signal_4479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C ( clk ), .D ( new_AGEMA_signal_4484 ), .Q ( new_AGEMA_signal_4485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C ( clk ), .D ( new_AGEMA_signal_4490 ), .Q ( new_AGEMA_signal_4491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C ( clk ), .D ( new_AGEMA_signal_4498 ), .Q ( new_AGEMA_signal_4499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C ( clk ), .D ( new_AGEMA_signal_4506 ), .Q ( new_AGEMA_signal_4507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C ( clk ), .D ( new_AGEMA_signal_4150 ), .Q ( new_AGEMA_signal_4509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C ( clk ), .D ( new_AGEMA_signal_4152 ), .Q ( new_AGEMA_signal_4511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C ( clk ), .D ( new_AGEMA_signal_4516 ), .Q ( new_AGEMA_signal_4517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C ( clk ), .D ( new_AGEMA_signal_4522 ), .Q ( new_AGEMA_signal_4523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C ( clk ), .D ( n2410 ), .Q ( new_AGEMA_signal_4525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C ( clk ), .D ( new_AGEMA_signal_1632 ), .Q ( new_AGEMA_signal_4527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C ( clk ), .D ( n2421 ), .Q ( new_AGEMA_signal_4529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C ( clk ), .D ( new_AGEMA_signal_1633 ), .Q ( new_AGEMA_signal_4531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C ( clk ), .D ( new_AGEMA_signal_4536 ), .Q ( new_AGEMA_signal_4537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C ( clk ), .D ( new_AGEMA_signal_4542 ), .Q ( new_AGEMA_signal_4543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C ( clk ), .D ( new_AGEMA_signal_4548 ), .Q ( new_AGEMA_signal_4549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C ( clk ), .D ( new_AGEMA_signal_4554 ), .Q ( new_AGEMA_signal_4555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C ( clk ), .D ( new_AGEMA_signal_4562 ), .Q ( new_AGEMA_signal_4563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C ( clk ), .D ( new_AGEMA_signal_4570 ), .Q ( new_AGEMA_signal_4571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C ( clk ), .D ( new_AGEMA_signal_4578 ), .Q ( new_AGEMA_signal_4579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C ( clk ), .D ( new_AGEMA_signal_4586 ), .Q ( new_AGEMA_signal_4587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C ( clk ), .D ( new_AGEMA_signal_4592 ), .Q ( new_AGEMA_signal_4593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C ( clk ), .D ( new_AGEMA_signal_4598 ), .Q ( new_AGEMA_signal_4599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C ( clk ), .D ( new_AGEMA_signal_4604 ), .Q ( new_AGEMA_signal_4605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C ( clk ), .D ( new_AGEMA_signal_4610 ), .Q ( new_AGEMA_signal_4611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C ( clk ), .D ( new_AGEMA_signal_4132 ), .Q ( new_AGEMA_signal_4613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C ( clk ), .D ( new_AGEMA_signal_4136 ), .Q ( new_AGEMA_signal_4615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C ( clk ), .D ( new_AGEMA_signal_4618 ), .Q ( new_AGEMA_signal_4619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C ( clk ), .D ( new_AGEMA_signal_4622 ), .Q ( new_AGEMA_signal_4623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C ( clk ), .D ( new_AGEMA_signal_4626 ), .Q ( new_AGEMA_signal_4627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C ( clk ), .D ( new_AGEMA_signal_4630 ), .Q ( new_AGEMA_signal_4631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C ( clk ), .D ( new_AGEMA_signal_4634 ), .Q ( new_AGEMA_signal_4635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C ( clk ), .D ( new_AGEMA_signal_4638 ), .Q ( new_AGEMA_signal_4639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C ( clk ), .D ( new_AGEMA_signal_4024 ), .Q ( new_AGEMA_signal_4641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C ( clk ), .D ( new_AGEMA_signal_4032 ), .Q ( new_AGEMA_signal_4643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C ( clk ), .D ( new_AGEMA_signal_4646 ), .Q ( new_AGEMA_signal_4647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C ( clk ), .D ( new_AGEMA_signal_4652 ), .Q ( new_AGEMA_signal_4653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C ( clk ), .D ( n1984 ), .Q ( new_AGEMA_signal_4661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C ( clk ), .D ( new_AGEMA_signal_1669 ), .Q ( new_AGEMA_signal_4665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C ( clk ), .D ( new_AGEMA_signal_4672 ), .Q ( new_AGEMA_signal_4673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C ( clk ), .D ( new_AGEMA_signal_4680 ), .Q ( new_AGEMA_signal_4681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C ( clk ), .D ( new_AGEMA_signal_4688 ), .Q ( new_AGEMA_signal_4689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C ( clk ), .D ( new_AGEMA_signal_4696 ), .Q ( new_AGEMA_signal_4697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C ( clk ), .D ( new_AGEMA_signal_4704 ), .Q ( new_AGEMA_signal_4705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C ( clk ), .D ( new_AGEMA_signal_4712 ), .Q ( new_AGEMA_signal_4713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C ( clk ), .D ( new_AGEMA_signal_4720 ), .Q ( new_AGEMA_signal_4721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C ( clk ), .D ( new_AGEMA_signal_4728 ), .Q ( new_AGEMA_signal_4729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C ( clk ), .D ( new_AGEMA_signal_4734 ), .Q ( new_AGEMA_signal_4735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C ( clk ), .D ( new_AGEMA_signal_4740 ), .Q ( new_AGEMA_signal_4741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C ( clk ), .D ( new_AGEMA_signal_4750 ), .Q ( new_AGEMA_signal_4751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C ( clk ), .D ( new_AGEMA_signal_4760 ), .Q ( new_AGEMA_signal_4761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C ( clk ), .D ( new_AGEMA_signal_4768 ), .Q ( new_AGEMA_signal_4769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C ( clk ), .D ( new_AGEMA_signal_4776 ), .Q ( new_AGEMA_signal_4777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C ( clk ), .D ( new_AGEMA_signal_4784 ), .Q ( new_AGEMA_signal_4785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C ( clk ), .D ( new_AGEMA_signal_4792 ), .Q ( new_AGEMA_signal_4793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C ( clk ), .D ( new_AGEMA_signal_4800 ), .Q ( new_AGEMA_signal_4801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C ( clk ), .D ( new_AGEMA_signal_4808 ), .Q ( new_AGEMA_signal_4809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C ( clk ), .D ( new_AGEMA_signal_4144 ), .Q ( new_AGEMA_signal_4817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C ( clk ), .D ( new_AGEMA_signal_4148 ), .Q ( new_AGEMA_signal_4821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C ( clk ), .D ( new_AGEMA_signal_4826 ), .Q ( new_AGEMA_signal_4827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C ( clk ), .D ( new_AGEMA_signal_4832 ), .Q ( new_AGEMA_signal_4833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C ( clk ), .D ( new_AGEMA_signal_3922 ), .Q ( new_AGEMA_signal_4837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C ( clk ), .D ( new_AGEMA_signal_3928 ), .Q ( new_AGEMA_signal_4841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C ( clk ), .D ( new_AGEMA_signal_4850 ), .Q ( new_AGEMA_signal_4851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C ( clk ), .D ( new_AGEMA_signal_4860 ), .Q ( new_AGEMA_signal_4861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C ( clk ), .D ( new_AGEMA_signal_4868 ), .Q ( new_AGEMA_signal_4869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C ( clk ), .D ( new_AGEMA_signal_4876 ), .Q ( new_AGEMA_signal_4877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C ( clk ), .D ( n2478 ), .Q ( new_AGEMA_signal_4881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C ( clk ), .D ( new_AGEMA_signal_1553 ), .Q ( new_AGEMA_signal_4885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C ( clk ), .D ( new_AGEMA_signal_4896 ), .Q ( new_AGEMA_signal_4897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C ( clk ), .D ( new_AGEMA_signal_4904 ), .Q ( new_AGEMA_signal_4905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C ( clk ), .D ( new_AGEMA_signal_4912 ), .Q ( new_AGEMA_signal_4913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C ( clk ), .D ( new_AGEMA_signal_4920 ), .Q ( new_AGEMA_signal_4921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C ( clk ), .D ( new_AGEMA_signal_4926 ), .Q ( new_AGEMA_signal_4927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C ( clk ), .D ( new_AGEMA_signal_4932 ), .Q ( new_AGEMA_signal_4933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C ( clk ), .D ( n2660 ), .Q ( new_AGEMA_signal_4937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_4941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C ( clk ), .D ( new_AGEMA_signal_4948 ), .Q ( new_AGEMA_signal_4949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C ( clk ), .D ( new_AGEMA_signal_4956 ), .Q ( new_AGEMA_signal_4957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C ( clk ), .D ( n1940 ), .Q ( new_AGEMA_signal_4965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C ( clk ), .D ( new_AGEMA_signal_1587 ), .Q ( new_AGEMA_signal_4971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C ( clk ), .D ( n1961 ), .Q ( new_AGEMA_signal_4977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C ( clk ), .D ( new_AGEMA_signal_1588 ), .Q ( new_AGEMA_signal_4983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C ( clk ), .D ( n1987 ), .Q ( new_AGEMA_signal_4989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C ( clk ), .D ( new_AGEMA_signal_1485 ), .Q ( new_AGEMA_signal_4995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C ( clk ), .D ( new_AGEMA_signal_5010 ), .Q ( new_AGEMA_signal_5011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C ( clk ), .D ( new_AGEMA_signal_5018 ), .Q ( new_AGEMA_signal_5019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C ( clk ), .D ( n2054 ), .Q ( new_AGEMA_signal_5025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C ( clk ), .D ( new_AGEMA_signal_1598 ), .Q ( new_AGEMA_signal_5031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C ( clk ), .D ( new_AGEMA_signal_5046 ), .Q ( new_AGEMA_signal_5047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C ( clk ), .D ( new_AGEMA_signal_5054 ), .Q ( new_AGEMA_signal_5055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C ( clk ), .D ( new_AGEMA_signal_5062 ), .Q ( new_AGEMA_signal_5063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C ( clk ), .D ( new_AGEMA_signal_5070 ), .Q ( new_AGEMA_signal_5071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C ( clk ), .D ( new_AGEMA_signal_5080 ), .Q ( new_AGEMA_signal_5081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C ( clk ), .D ( new_AGEMA_signal_5090 ), .Q ( new_AGEMA_signal_5091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C ( clk ), .D ( new_AGEMA_signal_5098 ), .Q ( new_AGEMA_signal_5099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C ( clk ), .D ( new_AGEMA_signal_5106 ), .Q ( new_AGEMA_signal_5107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C ( clk ), .D ( n2255 ), .Q ( new_AGEMA_signal_5113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C ( clk ), .D ( new_AGEMA_signal_1618 ), .Q ( new_AGEMA_signal_5119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C ( clk ), .D ( n2304 ), .Q ( new_AGEMA_signal_5133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C ( clk ), .D ( new_AGEMA_signal_1622 ), .Q ( new_AGEMA_signal_5139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C ( clk ), .D ( new_AGEMA_signal_5146 ), .Q ( new_AGEMA_signal_5147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C ( clk ), .D ( new_AGEMA_signal_5154 ), .Q ( new_AGEMA_signal_5155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C ( clk ), .D ( n2450 ), .Q ( new_AGEMA_signal_5161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C ( clk ), .D ( new_AGEMA_signal_1636 ), .Q ( new_AGEMA_signal_5167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C ( clk ), .D ( new_AGEMA_signal_5178 ), .Q ( new_AGEMA_signal_5179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C ( clk ), .D ( new_AGEMA_signal_5186 ), .Q ( new_AGEMA_signal_5187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C ( clk ), .D ( n2666 ), .Q ( new_AGEMA_signal_5201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C ( clk ), .D ( new_AGEMA_signal_1655 ), .Q ( new_AGEMA_signal_5207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C ( clk ), .D ( n2704 ), .Q ( new_AGEMA_signal_5213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C ( clk ), .D ( new_AGEMA_signal_1657 ), .Q ( new_AGEMA_signal_5219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C ( clk ), .D ( new_AGEMA_signal_5266 ), .Q ( new_AGEMA_signal_5267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C ( clk ), .D ( new_AGEMA_signal_5276 ), .Q ( new_AGEMA_signal_5277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C ( clk ), .D ( n2280 ), .Q ( new_AGEMA_signal_5325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C ( clk ), .D ( new_AGEMA_signal_1526 ), .Q ( new_AGEMA_signal_5333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C ( clk ), .D ( new_AGEMA_signal_3914 ), .Q ( new_AGEMA_signal_5353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C ( clk ), .D ( new_AGEMA_signal_3916 ), .Q ( new_AGEMA_signal_5361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C ( clk ), .D ( n2456 ), .Q ( new_AGEMA_signal_5369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C ( clk ), .D ( new_AGEMA_signal_1637 ), .Q ( new_AGEMA_signal_5377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C ( clk ), .D ( n2706 ), .Q ( new_AGEMA_signal_5405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C ( clk ), .D ( new_AGEMA_signal_1656 ), .Q ( new_AGEMA_signal_5413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C ( clk ), .D ( new_AGEMA_signal_5446 ), .Q ( new_AGEMA_signal_5447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C ( clk ), .D ( new_AGEMA_signal_5458 ), .Q ( new_AGEMA_signal_5459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C ( clk ), .D ( new_AGEMA_signal_5472 ), .Q ( new_AGEMA_signal_5473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C ( clk ), .D ( new_AGEMA_signal_5486 ), .Q ( new_AGEMA_signal_5487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C ( clk ), .D ( new_AGEMA_signal_5516 ), .Q ( new_AGEMA_signal_5517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C ( clk ), .D ( new_AGEMA_signal_5530 ), .Q ( new_AGEMA_signal_5531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C ( clk ), .D ( new_AGEMA_signal_5588 ), .Q ( new_AGEMA_signal_5589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C ( clk ), .D ( new_AGEMA_signal_5604 ), .Q ( new_AGEMA_signal_5605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C ( clk ), .D ( new_AGEMA_signal_5632 ), .Q ( new_AGEMA_signal_5633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C ( clk ), .D ( new_AGEMA_signal_5648 ), .Q ( new_AGEMA_signal_5649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C ( clk ), .D ( new_AGEMA_signal_5730 ), .Q ( new_AGEMA_signal_5731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C ( clk ), .D ( new_AGEMA_signal_5746 ), .Q ( new_AGEMA_signal_5747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C ( clk ), .D ( new_AGEMA_signal_5784 ), .Q ( new_AGEMA_signal_5785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C ( clk ), .D ( new_AGEMA_signal_5802 ), .Q ( new_AGEMA_signal_5803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C ( clk ), .D ( new_AGEMA_signal_5884 ), .Q ( new_AGEMA_signal_5885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C ( clk ), .D ( new_AGEMA_signal_5904 ), .Q ( new_AGEMA_signal_5905 ) ) ;

    /* cells in depth 12 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2001 ( .a ({new_AGEMA_signal_1586, n1932}), .b ({new_AGEMA_signal_3836, new_AGEMA_signal_3832}), .clk ( clk ), .r ( Fresh[660] ), .c ({new_AGEMA_signal_1667, n1933}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2051 ( .a ({new_AGEMA_signal_3844, new_AGEMA_signal_3840}), .b ({new_AGEMA_signal_1589, n1955}), .clk ( clk ), .r ( Fresh[661] ), .c ({new_AGEMA_signal_1668, n1958}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2067 ( .a ({new_AGEMA_signal_1479, n1967}), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3852}), .clk ( clk ), .r ( Fresh[662] ), .c ({new_AGEMA_signal_1590, n1990}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2104 ( .a ({new_AGEMA_signal_3864, new_AGEMA_signal_3862}), .b ({new_AGEMA_signal_1592, n1977}), .clk ( clk ), .r ( Fresh[663] ), .c ({new_AGEMA_signal_1670, n1982}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2128 ( .a ({new_AGEMA_signal_3880, new_AGEMA_signal_3872}), .b ({new_AGEMA_signal_1594, n1998}), .clk ( clk ), .r ( Fresh[664] ), .c ({new_AGEMA_signal_1671, n1999}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2148 ( .a ({new_AGEMA_signal_1595, n2010}), .b ({new_AGEMA_signal_3892, new_AGEMA_signal_3886}), .clk ( clk ), .r ( Fresh[665] ), .c ({new_AGEMA_signal_1672, n2011}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2165 ( .a ({new_AGEMA_signal_1489, n2024}), .b ({new_AGEMA_signal_3900, new_AGEMA_signal_3896}), .clk ( clk ), .r ( Fresh[666] ), .c ({new_AGEMA_signal_1596, n2025}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2179 ( .a ({new_AGEMA_signal_1597, n2035}), .b ({new_AGEMA_signal_3912, new_AGEMA_signal_3906}), .clk ( clk ), .r ( Fresh[667] ), .c ({new_AGEMA_signal_1674, n2036}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2196 ( .a ({new_AGEMA_signal_1599, n2048}), .b ({new_AGEMA_signal_1600, n2047}), .clk ( clk ), .r ( Fresh[668] ), .c ({new_AGEMA_signal_1675, n2049}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2207 ( .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3914}), .b ({new_AGEMA_signal_1601, n2059}), .clk ( clk ), .r ( Fresh[669] ), .c ({new_AGEMA_signal_1676, n2072}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2214 ( .a ({new_AGEMA_signal_3928, new_AGEMA_signal_3922}), .b ({new_AGEMA_signal_1602, n2064}), .clk ( clk ), .r ( Fresh[670] ), .c ({new_AGEMA_signal_1677, n2067}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2230 ( .a ({new_AGEMA_signal_3940, new_AGEMA_signal_3934}), .b ({new_AGEMA_signal_1603, n2077}), .clk ( clk ), .r ( Fresh[671] ), .c ({new_AGEMA_signal_1678, n2078}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2250 ( .a ({new_AGEMA_signal_3944, new_AGEMA_signal_3942}), .b ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .r ( Fresh[672] ), .c ({new_AGEMA_signal_1679, n2097}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2257 ( .a ({new_AGEMA_signal_1605, n2095}), .b ({new_AGEMA_signal_3952, new_AGEMA_signal_3948}), .clk ( clk ), .r ( Fresh[673] ), .c ({new_AGEMA_signal_1680, n2096}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2275 ( .a ({new_AGEMA_signal_3964, new_AGEMA_signal_3958}), .b ({new_AGEMA_signal_1681, n2117}), .clk ( clk ), .r ( Fresh[674] ), .c ({new_AGEMA_signal_1735, n2128}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2285 ( .a ({new_AGEMA_signal_1607, n2123}), .b ({new_AGEMA_signal_3976, new_AGEMA_signal_3970}), .clk ( clk ), .r ( Fresh[675] ), .c ({new_AGEMA_signal_1682, n2124}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2301 ( .a ({new_AGEMA_signal_3980, new_AGEMA_signal_3978}), .b ({new_AGEMA_signal_1507, n2135}), .clk ( clk ), .r ( Fresh[676] ), .c ({new_AGEMA_signal_1608, n2148}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2310 ( .a ({new_AGEMA_signal_3992, new_AGEMA_signal_3986}), .b ({new_AGEMA_signal_1609, n2141}), .clk ( clk ), .r ( Fresh[677] ), .c ({new_AGEMA_signal_1683, n2142}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2325 ( .a ({new_AGEMA_signal_3996, new_AGEMA_signal_3994}), .b ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .r ( Fresh[678] ), .c ({new_AGEMA_signal_1684, n2168}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2332 ( .a ({new_AGEMA_signal_1610, n2166}), .b ({new_AGEMA_signal_1512, n2165}), .clk ( clk ), .r ( Fresh[679] ), .c ({new_AGEMA_signal_1685, n2167}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2347 ( .a ({new_AGEMA_signal_4004, new_AGEMA_signal_4000}), .b ({new_AGEMA_signal_1611, n2180}), .clk ( clk ), .r ( Fresh[680] ), .c ({new_AGEMA_signal_1686, n2184}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2361 ( .a ({new_AGEMA_signal_4012, new_AGEMA_signal_4008}), .b ({new_AGEMA_signal_1612, n2194}), .clk ( clk ), .r ( Fresh[681] ), .c ({new_AGEMA_signal_1687, n2197}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2373 ( .a ({new_AGEMA_signal_4016, new_AGEMA_signal_4014}), .b ({new_AGEMA_signal_1688, n2204}), .clk ( clk ), .r ( Fresh[682] ), .c ({new_AGEMA_signal_1741, n2205}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2390 ( .a ({new_AGEMA_signal_4032, new_AGEMA_signal_4024}), .b ({new_AGEMA_signal_1614, n2225}), .clk ( clk ), .r ( Fresh[683] ), .c ({new_AGEMA_signal_1689, n2232}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2395 ( .a ({new_AGEMA_signal_1519, n2230}), .b ({new_AGEMA_signal_4044, new_AGEMA_signal_4038}), .clk ( clk ), .r ( Fresh[684] ), .c ({new_AGEMA_signal_1615, n2231}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2401 ( .a ({new_AGEMA_signal_4052, new_AGEMA_signal_4048}), .b ({new_AGEMA_signal_1690, n2236}), .clk ( clk ), .r ( Fresh[685] ), .c ({new_AGEMA_signal_1743, n2239}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2413 ( .a ({new_AGEMA_signal_4060, new_AGEMA_signal_4056}), .b ({new_AGEMA_signal_1617, n2247}), .clk ( clk ), .r ( Fresh[686] ), .c ({new_AGEMA_signal_1691, n2250}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2428 ( .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3914}), .b ({new_AGEMA_signal_1619, n2264}), .clk ( clk ), .r ( Fresh[687] ), .c ({new_AGEMA_signal_1692, n2276}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2439 ( .a ({new_AGEMA_signal_1620, n2271}), .b ({new_AGEMA_signal_4064, new_AGEMA_signal_4062}), .clk ( clk ), .r ( Fresh[688] ), .c ({new_AGEMA_signal_1693, n2272}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2454 ( .a ({new_AGEMA_signal_1527, n2286}), .b ({new_AGEMA_signal_4068, new_AGEMA_signal_4066}), .clk ( clk ), .r ( Fresh[689] ), .c ({new_AGEMA_signal_1621, n2306}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2468 ( .a ({new_AGEMA_signal_1623, n2295}), .b ({new_AGEMA_signal_4076, new_AGEMA_signal_4072}), .clk ( clk ), .r ( Fresh[690] ), .c ({new_AGEMA_signal_1694, n2296}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2489 ( .a ({new_AGEMA_signal_4084, new_AGEMA_signal_4080}), .b ({new_AGEMA_signal_1624, n2322}), .clk ( clk ), .r ( Fresh[691] ), .c ({new_AGEMA_signal_1695, n2324}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2500 ( .a ({new_AGEMA_signal_4088, new_AGEMA_signal_4086}), .b ({new_AGEMA_signal_1625, n2333}), .clk ( clk ), .r ( Fresh[692] ), .c ({new_AGEMA_signal_1696, n2337}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2511 ( .a ({new_AGEMA_signal_1627, n2345}), .b ({new_AGEMA_signal_4100, new_AGEMA_signal_4094}), .clk ( clk ), .r ( Fresh[693] ), .c ({new_AGEMA_signal_1697, n2350}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2528 ( .a ({new_AGEMA_signal_1628, n2361}), .b ({new_AGEMA_signal_4108, new_AGEMA_signal_4104}), .clk ( clk ), .r ( Fresh[694] ), .c ({new_AGEMA_signal_1698, n2362}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2550 ( .a ({new_AGEMA_signal_4112, new_AGEMA_signal_4110}), .b ({new_AGEMA_signal_1541, n2388}), .clk ( clk ), .r ( Fresh[695] ), .c ({new_AGEMA_signal_1629, n2389}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2557 ( .a ({new_AGEMA_signal_4120, new_AGEMA_signal_4116}), .b ({new_AGEMA_signal_1630, n2393}), .clk ( clk ), .r ( Fresh[696] ), .c ({new_AGEMA_signal_1700, n2397}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2568 ( .a ({new_AGEMA_signal_4128, new_AGEMA_signal_4124}), .b ({new_AGEMA_signal_1543, n2405}), .clk ( clk ), .r ( Fresh[697] ), .c ({new_AGEMA_signal_1631, n2411}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2580 ( .a ({new_AGEMA_signal_4136, new_AGEMA_signal_4132}), .b ({new_AGEMA_signal_1546, n2419}), .clk ( clk ), .r ( Fresh[698] ), .c ({new_AGEMA_signal_1634, n2420}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2593 ( .a ({new_AGEMA_signal_1635, n2436}), .b ({new_AGEMA_signal_4140, new_AGEMA_signal_4138}), .clk ( clk ), .r ( Fresh[699] ), .c ({new_AGEMA_signal_1703, n2440}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2614 ( .a ({new_AGEMA_signal_4148, new_AGEMA_signal_4144}), .b ({new_AGEMA_signal_1638, n2461}), .clk ( clk ), .r ( Fresh[700] ), .c ({new_AGEMA_signal_1704, n2516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2621 ( .s ({new_AGEMA_signal_4152, new_AGEMA_signal_4150}), .b ({new_AGEMA_signal_1552, n2469}), .a ({new_AGEMA_signal_4164, new_AGEMA_signal_4158}), .clk ( clk ), .r ( Fresh[701] ), .c ({new_AGEMA_signal_1639, n2471}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2636 ( .a ({new_AGEMA_signal_4176, new_AGEMA_signal_4170}), .b ({new_AGEMA_signal_1640, n2484}), .clk ( clk ), .r ( Fresh[702] ), .c ({new_AGEMA_signal_1706, n2485}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2644 ( .a ({new_AGEMA_signal_3928, new_AGEMA_signal_3922}), .b ({new_AGEMA_signal_1555, n2491}), .clk ( clk ), .r ( Fresh[703] ), .c ({new_AGEMA_signal_1641, n2502}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2651 ( .a ({new_AGEMA_signal_1642, n2500}), .b ({new_AGEMA_signal_4184, new_AGEMA_signal_4180}), .clk ( clk ), .r ( Fresh[704] ), .c ({new_AGEMA_signal_1707, n2501}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2657 ( .a ({new_AGEMA_signal_4136, new_AGEMA_signal_4132}), .b ({new_AGEMA_signal_1708, n2508}), .clk ( clk ), .r ( Fresh[705] ), .c ({new_AGEMA_signal_1757, n2509}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2671 ( .a ({new_AGEMA_signal_4188, new_AGEMA_signal_4186}), .b ({new_AGEMA_signal_1709, n2526}), .clk ( clk ), .r ( Fresh[706] ), .c ({new_AGEMA_signal_1758, n2527}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2680 ( .a ({new_AGEMA_signal_1645, n2539}), .b ({new_AGEMA_signal_4204, new_AGEMA_signal_4196}), .clk ( clk ), .r ( Fresh[707] ), .c ({new_AGEMA_signal_1710, n2550}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2685 ( .a ({new_AGEMA_signal_1646, n2548}), .b ({new_AGEMA_signal_4208, new_AGEMA_signal_4206}), .clk ( clk ), .r ( Fresh[708] ), .c ({new_AGEMA_signal_1711, n2549}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2701 ( .a ({new_AGEMA_signal_1647, n2568}), .b ({new_AGEMA_signal_1648, n2567}), .clk ( clk ), .r ( Fresh[709] ), .c ({new_AGEMA_signal_1712, n2569}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2712 ( .a ({new_AGEMA_signal_1649, n2583}), .b ({new_AGEMA_signal_4216, new_AGEMA_signal_4212}), .clk ( clk ), .r ( Fresh[710] ), .c ({new_AGEMA_signal_1713, n2584}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2729 ( .a ({new_AGEMA_signal_4224, new_AGEMA_signal_4220}), .b ({new_AGEMA_signal_1566, n2604}), .clk ( clk ), .r ( Fresh[711] ), .c ({new_AGEMA_signal_1650, n2606}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2740 ( .a ({new_AGEMA_signal_3928, new_AGEMA_signal_3922}), .b ({new_AGEMA_signal_1651, n2621}), .clk ( clk ), .r ( Fresh[712] ), .c ({new_AGEMA_signal_1715, n2622}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2747 ( .a ({new_AGEMA_signal_1652, n2633}), .b ({new_AGEMA_signal_4232, new_AGEMA_signal_4228}), .clk ( clk ), .r ( Fresh[713] ), .c ({new_AGEMA_signal_1716, n2634}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2761 ( .a ({new_AGEMA_signal_1654, n2656}), .b ({new_AGEMA_signal_4240, new_AGEMA_signal_4236}), .clk ( clk ), .r ( Fresh[714] ), .c ({new_AGEMA_signal_1717, n2657}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2783 ( .a ({new_AGEMA_signal_1658, n2696}), .b ({new_AGEMA_signal_4248, new_AGEMA_signal_4244}), .clk ( clk ), .r ( Fresh[715] ), .c ({new_AGEMA_signal_1718, n2697}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2795 ( .a ({new_AGEMA_signal_3916, new_AGEMA_signal_3914}), .b ({new_AGEMA_signal_1659, n2718}), .clk ( clk ), .r ( Fresh[716] ), .c ({new_AGEMA_signal_1719, n2808}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2802 ( .a ({new_AGEMA_signal_1660, n2730}), .b ({new_AGEMA_signal_4264, new_AGEMA_signal_4256}), .clk ( clk ), .r ( Fresh[717] ), .c ({new_AGEMA_signal_1720, n2747}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2810 ( .a ({new_AGEMA_signal_1661, n2745}), .b ({new_AGEMA_signal_1662, n2744}), .clk ( clk ), .r ( Fresh[718] ), .c ({new_AGEMA_signal_1721, n2746}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2818 ( .a ({new_AGEMA_signal_1663, n2759}), .b ({new_AGEMA_signal_4268, new_AGEMA_signal_4266}), .clk ( clk ), .r ( Fresh[719] ), .c ({new_AGEMA_signal_1722, n2804}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2824 ( .a ({new_AGEMA_signal_1664, n2771}), .b ({new_AGEMA_signal_4276, new_AGEMA_signal_4272}), .clk ( clk ), .r ( Fresh[720] ), .c ({new_AGEMA_signal_1723, n2802}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2838 ( .a ({new_AGEMA_signal_1582, n2798}), .b ({new_AGEMA_signal_4280, new_AGEMA_signal_4278}), .clk ( clk ), .r ( Fresh[721] ), .c ({new_AGEMA_signal_1665, n2799}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2852 ( .a ({new_AGEMA_signal_1666, n2826}), .b ({new_AGEMA_signal_4292, new_AGEMA_signal_4286}), .clk ( clk ), .r ( Fresh[722] ), .c ({new_AGEMA_signal_1725, n2827}) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C ( clk ), .D ( new_AGEMA_signal_4293 ), .Q ( new_AGEMA_signal_4294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C ( clk ), .D ( new_AGEMA_signal_4295 ), .Q ( new_AGEMA_signal_4296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C ( clk ), .D ( new_AGEMA_signal_4303 ), .Q ( new_AGEMA_signal_4304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C ( clk ), .D ( new_AGEMA_signal_4311 ), .Q ( new_AGEMA_signal_4312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C ( clk ), .D ( new_AGEMA_signal_4313 ), .Q ( new_AGEMA_signal_4314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C ( clk ), .D ( new_AGEMA_signal_4315 ), .Q ( new_AGEMA_signal_4316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C ( clk ), .D ( new_AGEMA_signal_4319 ), .Q ( new_AGEMA_signal_4320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C ( clk ), .D ( new_AGEMA_signal_4323 ), .Q ( new_AGEMA_signal_4324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C ( clk ), .D ( new_AGEMA_signal_4331 ), .Q ( new_AGEMA_signal_4332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C ( clk ), .D ( new_AGEMA_signal_4339 ), .Q ( new_AGEMA_signal_4340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C ( clk ), .D ( new_AGEMA_signal_4341 ), .Q ( new_AGEMA_signal_4342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C ( clk ), .D ( new_AGEMA_signal_4343 ), .Q ( new_AGEMA_signal_4344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C ( clk ), .D ( new_AGEMA_signal_4349 ), .Q ( new_AGEMA_signal_4350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C ( clk ), .D ( new_AGEMA_signal_4355 ), .Q ( new_AGEMA_signal_4356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C ( clk ), .D ( new_AGEMA_signal_4359 ), .Q ( new_AGEMA_signal_4360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C ( clk ), .D ( new_AGEMA_signal_4363 ), .Q ( new_AGEMA_signal_4364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C ( clk ), .D ( new_AGEMA_signal_4371 ), .Q ( new_AGEMA_signal_4372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C ( clk ), .D ( new_AGEMA_signal_4379 ), .Q ( new_AGEMA_signal_4380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C ( clk ), .D ( new_AGEMA_signal_4383 ), .Q ( new_AGEMA_signal_4384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C ( clk ), .D ( new_AGEMA_signal_4387 ), .Q ( new_AGEMA_signal_4388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C ( clk ), .D ( new_AGEMA_signal_4393 ), .Q ( new_AGEMA_signal_4394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C ( clk ), .D ( new_AGEMA_signal_4399 ), .Q ( new_AGEMA_signal_4400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C ( clk ), .D ( new_AGEMA_signal_4405 ), .Q ( new_AGEMA_signal_4406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C ( clk ), .D ( new_AGEMA_signal_4411 ), .Q ( new_AGEMA_signal_4412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C ( clk ), .D ( new_AGEMA_signal_4417 ), .Q ( new_AGEMA_signal_4418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C ( clk ), .D ( new_AGEMA_signal_4423 ), .Q ( new_AGEMA_signal_4424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C ( clk ), .D ( new_AGEMA_signal_4429 ), .Q ( new_AGEMA_signal_4430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C ( clk ), .D ( new_AGEMA_signal_4435 ), .Q ( new_AGEMA_signal_4436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C ( clk ), .D ( new_AGEMA_signal_4441 ), .Q ( new_AGEMA_signal_4442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C ( clk ), .D ( new_AGEMA_signal_4447 ), .Q ( new_AGEMA_signal_4448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C ( clk ), .D ( new_AGEMA_signal_4451 ), .Q ( new_AGEMA_signal_4452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C ( clk ), .D ( new_AGEMA_signal_4455 ), .Q ( new_AGEMA_signal_4456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C ( clk ), .D ( new_AGEMA_signal_4463 ), .Q ( new_AGEMA_signal_4464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C ( clk ), .D ( new_AGEMA_signal_4471 ), .Q ( new_AGEMA_signal_4472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C ( clk ), .D ( new_AGEMA_signal_4475 ), .Q ( new_AGEMA_signal_4476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C ( clk ), .D ( new_AGEMA_signal_4479 ), .Q ( new_AGEMA_signal_4480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C ( clk ), .D ( new_AGEMA_signal_4485 ), .Q ( new_AGEMA_signal_4486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C ( clk ), .D ( new_AGEMA_signal_4491 ), .Q ( new_AGEMA_signal_4492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C ( clk ), .D ( new_AGEMA_signal_4499 ), .Q ( new_AGEMA_signal_4500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C ( clk ), .D ( new_AGEMA_signal_4507 ), .Q ( new_AGEMA_signal_4508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C ( clk ), .D ( new_AGEMA_signal_4509 ), .Q ( new_AGEMA_signal_4510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C ( clk ), .D ( new_AGEMA_signal_4511 ), .Q ( new_AGEMA_signal_4512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C ( clk ), .D ( new_AGEMA_signal_4517 ), .Q ( new_AGEMA_signal_4518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C ( clk ), .D ( new_AGEMA_signal_4523 ), .Q ( new_AGEMA_signal_4524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C ( clk ), .D ( new_AGEMA_signal_4525 ), .Q ( new_AGEMA_signal_4526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C ( clk ), .D ( new_AGEMA_signal_4527 ), .Q ( new_AGEMA_signal_4528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C ( clk ), .D ( new_AGEMA_signal_4529 ), .Q ( new_AGEMA_signal_4530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C ( clk ), .D ( new_AGEMA_signal_4531 ), .Q ( new_AGEMA_signal_4532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C ( clk ), .D ( new_AGEMA_signal_4537 ), .Q ( new_AGEMA_signal_4538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C ( clk ), .D ( new_AGEMA_signal_4543 ), .Q ( new_AGEMA_signal_4544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C ( clk ), .D ( new_AGEMA_signal_4549 ), .Q ( new_AGEMA_signal_4550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C ( clk ), .D ( new_AGEMA_signal_4555 ), .Q ( new_AGEMA_signal_4556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C ( clk ), .D ( new_AGEMA_signal_4563 ), .Q ( new_AGEMA_signal_4564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C ( clk ), .D ( new_AGEMA_signal_4571 ), .Q ( new_AGEMA_signal_4572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C ( clk ), .D ( new_AGEMA_signal_4579 ), .Q ( new_AGEMA_signal_4580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C ( clk ), .D ( new_AGEMA_signal_4587 ), .Q ( new_AGEMA_signal_4588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C ( clk ), .D ( new_AGEMA_signal_4593 ), .Q ( new_AGEMA_signal_4594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C ( clk ), .D ( new_AGEMA_signal_4599 ), .Q ( new_AGEMA_signal_4600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C ( clk ), .D ( new_AGEMA_signal_4605 ), .Q ( new_AGEMA_signal_4606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C ( clk ), .D ( new_AGEMA_signal_4611 ), .Q ( new_AGEMA_signal_4612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C ( clk ), .D ( new_AGEMA_signal_4613 ), .Q ( new_AGEMA_signal_4614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C ( clk ), .D ( new_AGEMA_signal_4615 ), .Q ( new_AGEMA_signal_4616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C ( clk ), .D ( new_AGEMA_signal_4619 ), .Q ( new_AGEMA_signal_4620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C ( clk ), .D ( new_AGEMA_signal_4623 ), .Q ( new_AGEMA_signal_4624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C ( clk ), .D ( new_AGEMA_signal_4627 ), .Q ( new_AGEMA_signal_4628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C ( clk ), .D ( new_AGEMA_signal_4631 ), .Q ( new_AGEMA_signal_4632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C ( clk ), .D ( new_AGEMA_signal_4635 ), .Q ( new_AGEMA_signal_4636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C ( clk ), .D ( new_AGEMA_signal_4639 ), .Q ( new_AGEMA_signal_4640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C ( clk ), .D ( new_AGEMA_signal_4641 ), .Q ( new_AGEMA_signal_4642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C ( clk ), .D ( new_AGEMA_signal_4643 ), .Q ( new_AGEMA_signal_4644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C ( clk ), .D ( new_AGEMA_signal_4647 ), .Q ( new_AGEMA_signal_4648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C ( clk ), .D ( new_AGEMA_signal_4653 ), .Q ( new_AGEMA_signal_4654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C ( clk ), .D ( new_AGEMA_signal_4661 ), .Q ( new_AGEMA_signal_4662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C ( clk ), .D ( new_AGEMA_signal_4665 ), .Q ( new_AGEMA_signal_4666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C ( clk ), .D ( new_AGEMA_signal_4673 ), .Q ( new_AGEMA_signal_4674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C ( clk ), .D ( new_AGEMA_signal_4681 ), .Q ( new_AGEMA_signal_4682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C ( clk ), .D ( new_AGEMA_signal_4689 ), .Q ( new_AGEMA_signal_4690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C ( clk ), .D ( new_AGEMA_signal_4697 ), .Q ( new_AGEMA_signal_4698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C ( clk ), .D ( new_AGEMA_signal_4705 ), .Q ( new_AGEMA_signal_4706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C ( clk ), .D ( new_AGEMA_signal_4713 ), .Q ( new_AGEMA_signal_4714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C ( clk ), .D ( new_AGEMA_signal_4721 ), .Q ( new_AGEMA_signal_4722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C ( clk ), .D ( new_AGEMA_signal_4729 ), .Q ( new_AGEMA_signal_4730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C ( clk ), .D ( new_AGEMA_signal_4735 ), .Q ( new_AGEMA_signal_4736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C ( clk ), .D ( new_AGEMA_signal_4741 ), .Q ( new_AGEMA_signal_4742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C ( clk ), .D ( new_AGEMA_signal_4751 ), .Q ( new_AGEMA_signal_4752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C ( clk ), .D ( new_AGEMA_signal_4761 ), .Q ( new_AGEMA_signal_4762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C ( clk ), .D ( new_AGEMA_signal_4769 ), .Q ( new_AGEMA_signal_4770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C ( clk ), .D ( new_AGEMA_signal_4777 ), .Q ( new_AGEMA_signal_4778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C ( clk ), .D ( new_AGEMA_signal_4785 ), .Q ( new_AGEMA_signal_4786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C ( clk ), .D ( new_AGEMA_signal_4793 ), .Q ( new_AGEMA_signal_4794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C ( clk ), .D ( new_AGEMA_signal_4801 ), .Q ( new_AGEMA_signal_4802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C ( clk ), .D ( new_AGEMA_signal_4809 ), .Q ( new_AGEMA_signal_4810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C ( clk ), .D ( new_AGEMA_signal_4817 ), .Q ( new_AGEMA_signal_4818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C ( clk ), .D ( new_AGEMA_signal_4821 ), .Q ( new_AGEMA_signal_4822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C ( clk ), .D ( new_AGEMA_signal_4827 ), .Q ( new_AGEMA_signal_4828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C ( clk ), .D ( new_AGEMA_signal_4833 ), .Q ( new_AGEMA_signal_4834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C ( clk ), .D ( new_AGEMA_signal_4837 ), .Q ( new_AGEMA_signal_4838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C ( clk ), .D ( new_AGEMA_signal_4841 ), .Q ( new_AGEMA_signal_4842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C ( clk ), .D ( new_AGEMA_signal_4851 ), .Q ( new_AGEMA_signal_4852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C ( clk ), .D ( new_AGEMA_signal_4861 ), .Q ( new_AGEMA_signal_4862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C ( clk ), .D ( new_AGEMA_signal_4869 ), .Q ( new_AGEMA_signal_4870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C ( clk ), .D ( new_AGEMA_signal_4877 ), .Q ( new_AGEMA_signal_4878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C ( clk ), .D ( new_AGEMA_signal_4881 ), .Q ( new_AGEMA_signal_4882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C ( clk ), .D ( new_AGEMA_signal_4885 ), .Q ( new_AGEMA_signal_4886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C ( clk ), .D ( new_AGEMA_signal_4897 ), .Q ( new_AGEMA_signal_4898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C ( clk ), .D ( new_AGEMA_signal_4905 ), .Q ( new_AGEMA_signal_4906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C ( clk ), .D ( new_AGEMA_signal_4913 ), .Q ( new_AGEMA_signal_4914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C ( clk ), .D ( new_AGEMA_signal_4921 ), .Q ( new_AGEMA_signal_4922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C ( clk ), .D ( new_AGEMA_signal_4927 ), .Q ( new_AGEMA_signal_4928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C ( clk ), .D ( new_AGEMA_signal_4933 ), .Q ( new_AGEMA_signal_4934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C ( clk ), .D ( new_AGEMA_signal_4937 ), .Q ( new_AGEMA_signal_4938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C ( clk ), .D ( new_AGEMA_signal_4941 ), .Q ( new_AGEMA_signal_4942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C ( clk ), .D ( new_AGEMA_signal_4949 ), .Q ( new_AGEMA_signal_4950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C ( clk ), .D ( new_AGEMA_signal_4957 ), .Q ( new_AGEMA_signal_4958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C ( clk ), .D ( new_AGEMA_signal_4965 ), .Q ( new_AGEMA_signal_4966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C ( clk ), .D ( new_AGEMA_signal_4971 ), .Q ( new_AGEMA_signal_4972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C ( clk ), .D ( new_AGEMA_signal_4977 ), .Q ( new_AGEMA_signal_4978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C ( clk ), .D ( new_AGEMA_signal_4983 ), .Q ( new_AGEMA_signal_4984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C ( clk ), .D ( new_AGEMA_signal_4989 ), .Q ( new_AGEMA_signal_4990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C ( clk ), .D ( new_AGEMA_signal_4995 ), .Q ( new_AGEMA_signal_4996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C ( clk ), .D ( new_AGEMA_signal_5011 ), .Q ( new_AGEMA_signal_5012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C ( clk ), .D ( new_AGEMA_signal_5019 ), .Q ( new_AGEMA_signal_5020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C ( clk ), .D ( new_AGEMA_signal_5025 ), .Q ( new_AGEMA_signal_5026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C ( clk ), .D ( new_AGEMA_signal_5031 ), .Q ( new_AGEMA_signal_5032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C ( clk ), .D ( new_AGEMA_signal_5047 ), .Q ( new_AGEMA_signal_5048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C ( clk ), .D ( new_AGEMA_signal_5055 ), .Q ( new_AGEMA_signal_5056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C ( clk ), .D ( new_AGEMA_signal_5063 ), .Q ( new_AGEMA_signal_5064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C ( clk ), .D ( new_AGEMA_signal_5071 ), .Q ( new_AGEMA_signal_5072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C ( clk ), .D ( new_AGEMA_signal_5081 ), .Q ( new_AGEMA_signal_5082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C ( clk ), .D ( new_AGEMA_signal_5091 ), .Q ( new_AGEMA_signal_5092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C ( clk ), .D ( new_AGEMA_signal_5099 ), .Q ( new_AGEMA_signal_5100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C ( clk ), .D ( new_AGEMA_signal_5107 ), .Q ( new_AGEMA_signal_5108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C ( clk ), .D ( new_AGEMA_signal_5113 ), .Q ( new_AGEMA_signal_5114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C ( clk ), .D ( new_AGEMA_signal_5119 ), .Q ( new_AGEMA_signal_5120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C ( clk ), .D ( new_AGEMA_signal_5133 ), .Q ( new_AGEMA_signal_5134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C ( clk ), .D ( new_AGEMA_signal_5139 ), .Q ( new_AGEMA_signal_5140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C ( clk ), .D ( new_AGEMA_signal_5147 ), .Q ( new_AGEMA_signal_5148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C ( clk ), .D ( new_AGEMA_signal_5155 ), .Q ( new_AGEMA_signal_5156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C ( clk ), .D ( new_AGEMA_signal_5161 ), .Q ( new_AGEMA_signal_5162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C ( clk ), .D ( new_AGEMA_signal_5167 ), .Q ( new_AGEMA_signal_5168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C ( clk ), .D ( new_AGEMA_signal_5179 ), .Q ( new_AGEMA_signal_5180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C ( clk ), .D ( new_AGEMA_signal_5187 ), .Q ( new_AGEMA_signal_5188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C ( clk ), .D ( new_AGEMA_signal_5201 ), .Q ( new_AGEMA_signal_5202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C ( clk ), .D ( new_AGEMA_signal_5207 ), .Q ( new_AGEMA_signal_5208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C ( clk ), .D ( new_AGEMA_signal_5213 ), .Q ( new_AGEMA_signal_5214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C ( clk ), .D ( new_AGEMA_signal_5219 ), .Q ( new_AGEMA_signal_5220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C ( clk ), .D ( new_AGEMA_signal_5267 ), .Q ( new_AGEMA_signal_5268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C ( clk ), .D ( new_AGEMA_signal_5277 ), .Q ( new_AGEMA_signal_5278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C ( clk ), .D ( new_AGEMA_signal_5325 ), .Q ( new_AGEMA_signal_5326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C ( clk ), .D ( new_AGEMA_signal_5333 ), .Q ( new_AGEMA_signal_5334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C ( clk ), .D ( new_AGEMA_signal_5353 ), .Q ( new_AGEMA_signal_5354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C ( clk ), .D ( new_AGEMA_signal_5361 ), .Q ( new_AGEMA_signal_5362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C ( clk ), .D ( new_AGEMA_signal_5369 ), .Q ( new_AGEMA_signal_5370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C ( clk ), .D ( new_AGEMA_signal_5377 ), .Q ( new_AGEMA_signal_5378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C ( clk ), .D ( new_AGEMA_signal_5405 ), .Q ( new_AGEMA_signal_5406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C ( clk ), .D ( new_AGEMA_signal_5413 ), .Q ( new_AGEMA_signal_5414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C ( clk ), .D ( new_AGEMA_signal_5447 ), .Q ( new_AGEMA_signal_5448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C ( clk ), .D ( new_AGEMA_signal_5459 ), .Q ( new_AGEMA_signal_5460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C ( clk ), .D ( new_AGEMA_signal_5473 ), .Q ( new_AGEMA_signal_5474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C ( clk ), .D ( new_AGEMA_signal_5487 ), .Q ( new_AGEMA_signal_5488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C ( clk ), .D ( new_AGEMA_signal_5517 ), .Q ( new_AGEMA_signal_5518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C ( clk ), .D ( new_AGEMA_signal_5531 ), .Q ( new_AGEMA_signal_5532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C ( clk ), .D ( new_AGEMA_signal_5589 ), .Q ( new_AGEMA_signal_5590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C ( clk ), .D ( new_AGEMA_signal_5605 ), .Q ( new_AGEMA_signal_5606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C ( clk ), .D ( new_AGEMA_signal_5633 ), .Q ( new_AGEMA_signal_5634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C ( clk ), .D ( new_AGEMA_signal_5649 ), .Q ( new_AGEMA_signal_5650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C ( clk ), .D ( new_AGEMA_signal_5731 ), .Q ( new_AGEMA_signal_5732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C ( clk ), .D ( new_AGEMA_signal_5747 ), .Q ( new_AGEMA_signal_5748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C ( clk ), .D ( new_AGEMA_signal_5785 ), .Q ( new_AGEMA_signal_5786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C ( clk ), .D ( new_AGEMA_signal_5803 ), .Q ( new_AGEMA_signal_5804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C ( clk ), .D ( new_AGEMA_signal_5885 ), .Q ( new_AGEMA_signal_5886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C ( clk ), .D ( new_AGEMA_signal_5905 ), .Q ( new_AGEMA_signal_5906 ) ) ;

    /* cells in depth 13 */
    buf_clk new_AGEMA_reg_buffer_2831 ( .C ( clk ), .D ( new_AGEMA_signal_4648 ), .Q ( new_AGEMA_signal_4649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C ( clk ), .D ( new_AGEMA_signal_4654 ), .Q ( new_AGEMA_signal_4655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C ( clk ), .D ( new_AGEMA_signal_4620 ), .Q ( new_AGEMA_signal_4657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C ( clk ), .D ( new_AGEMA_signal_4624 ), .Q ( new_AGEMA_signal_4659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C ( clk ), .D ( new_AGEMA_signal_4662 ), .Q ( new_AGEMA_signal_4663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C ( clk ), .D ( new_AGEMA_signal_4666 ), .Q ( new_AGEMA_signal_4667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C ( clk ), .D ( new_AGEMA_signal_4674 ), .Q ( new_AGEMA_signal_4675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C ( clk ), .D ( new_AGEMA_signal_4682 ), .Q ( new_AGEMA_signal_4683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C ( clk ), .D ( new_AGEMA_signal_4690 ), .Q ( new_AGEMA_signal_4691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C ( clk ), .D ( new_AGEMA_signal_4698 ), .Q ( new_AGEMA_signal_4699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C ( clk ), .D ( new_AGEMA_signal_4706 ), .Q ( new_AGEMA_signal_4707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C ( clk ), .D ( new_AGEMA_signal_4714 ), .Q ( new_AGEMA_signal_4715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C ( clk ), .D ( new_AGEMA_signal_4722 ), .Q ( new_AGEMA_signal_4723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C ( clk ), .D ( new_AGEMA_signal_4730 ), .Q ( new_AGEMA_signal_4731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C ( clk ), .D ( new_AGEMA_signal_4736 ), .Q ( new_AGEMA_signal_4737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C ( clk ), .D ( new_AGEMA_signal_4742 ), .Q ( new_AGEMA_signal_4743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C ( clk ), .D ( new_AGEMA_signal_4752 ), .Q ( new_AGEMA_signal_4753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C ( clk ), .D ( new_AGEMA_signal_4762 ), .Q ( new_AGEMA_signal_4763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C ( clk ), .D ( new_AGEMA_signal_4770 ), .Q ( new_AGEMA_signal_4771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C ( clk ), .D ( new_AGEMA_signal_4778 ), .Q ( new_AGEMA_signal_4779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C ( clk ), .D ( new_AGEMA_signal_4786 ), .Q ( new_AGEMA_signal_4787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C ( clk ), .D ( new_AGEMA_signal_4794 ), .Q ( new_AGEMA_signal_4795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C ( clk ), .D ( new_AGEMA_signal_4802 ), .Q ( new_AGEMA_signal_4803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C ( clk ), .D ( new_AGEMA_signal_4810 ), .Q ( new_AGEMA_signal_4811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C ( clk ), .D ( new_AGEMA_signal_4342 ), .Q ( new_AGEMA_signal_4813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C ( clk ), .D ( new_AGEMA_signal_4344 ), .Q ( new_AGEMA_signal_4815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C ( clk ), .D ( new_AGEMA_signal_4818 ), .Q ( new_AGEMA_signal_4819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C ( clk ), .D ( new_AGEMA_signal_4822 ), .Q ( new_AGEMA_signal_4823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C ( clk ), .D ( new_AGEMA_signal_4828 ), .Q ( new_AGEMA_signal_4829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C ( clk ), .D ( new_AGEMA_signal_4834 ), .Q ( new_AGEMA_signal_4835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C ( clk ), .D ( new_AGEMA_signal_4838 ), .Q ( new_AGEMA_signal_4839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C ( clk ), .D ( new_AGEMA_signal_4842 ), .Q ( new_AGEMA_signal_4843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C ( clk ), .D ( new_AGEMA_signal_4852 ), .Q ( new_AGEMA_signal_4853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C ( clk ), .D ( new_AGEMA_signal_4862 ), .Q ( new_AGEMA_signal_4863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C ( clk ), .D ( new_AGEMA_signal_4870 ), .Q ( new_AGEMA_signal_4871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C ( clk ), .D ( new_AGEMA_signal_4878 ), .Q ( new_AGEMA_signal_4879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C ( clk ), .D ( new_AGEMA_signal_4882 ), .Q ( new_AGEMA_signal_4883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C ( clk ), .D ( new_AGEMA_signal_4886 ), .Q ( new_AGEMA_signal_4887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C ( clk ), .D ( n2509 ), .Q ( new_AGEMA_signal_4889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C ( clk ), .D ( new_AGEMA_signal_1757 ), .Q ( new_AGEMA_signal_4891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C ( clk ), .D ( new_AGEMA_signal_4898 ), .Q ( new_AGEMA_signal_4899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C ( clk ), .D ( new_AGEMA_signal_4906 ), .Q ( new_AGEMA_signal_4907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C ( clk ), .D ( new_AGEMA_signal_4914 ), .Q ( new_AGEMA_signal_4915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C ( clk ), .D ( new_AGEMA_signal_4922 ), .Q ( new_AGEMA_signal_4923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C ( clk ), .D ( new_AGEMA_signal_4928 ), .Q ( new_AGEMA_signal_4929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C ( clk ), .D ( new_AGEMA_signal_4934 ), .Q ( new_AGEMA_signal_4935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C ( clk ), .D ( new_AGEMA_signal_4938 ), .Q ( new_AGEMA_signal_4939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C ( clk ), .D ( new_AGEMA_signal_4942 ), .Q ( new_AGEMA_signal_4943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C ( clk ), .D ( new_AGEMA_signal_4950 ), .Q ( new_AGEMA_signal_4951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C ( clk ), .D ( new_AGEMA_signal_4958 ), .Q ( new_AGEMA_signal_4959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C ( clk ), .D ( n2802 ), .Q ( new_AGEMA_signal_4961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C ( clk ), .D ( new_AGEMA_signal_1723 ), .Q ( new_AGEMA_signal_4963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C ( clk ), .D ( new_AGEMA_signal_4966 ), .Q ( new_AGEMA_signal_4967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C ( clk ), .D ( new_AGEMA_signal_4972 ), .Q ( new_AGEMA_signal_4973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C ( clk ), .D ( new_AGEMA_signal_4978 ), .Q ( new_AGEMA_signal_4979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C ( clk ), .D ( new_AGEMA_signal_4984 ), .Q ( new_AGEMA_signal_4985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C ( clk ), .D ( new_AGEMA_signal_4990 ), .Q ( new_AGEMA_signal_4991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C ( clk ), .D ( new_AGEMA_signal_4996 ), .Q ( new_AGEMA_signal_4997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C ( clk ), .D ( new_AGEMA_signal_4642 ), .Q ( new_AGEMA_signal_5001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C ( clk ), .D ( new_AGEMA_signal_4644 ), .Q ( new_AGEMA_signal_5005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C ( clk ), .D ( new_AGEMA_signal_5012 ), .Q ( new_AGEMA_signal_5013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C ( clk ), .D ( new_AGEMA_signal_5020 ), .Q ( new_AGEMA_signal_5021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C ( clk ), .D ( new_AGEMA_signal_5026 ), .Q ( new_AGEMA_signal_5027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C ( clk ), .D ( new_AGEMA_signal_5032 ), .Q ( new_AGEMA_signal_5033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C ( clk ), .D ( n2072 ), .Q ( new_AGEMA_signal_5037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C ( clk ), .D ( new_AGEMA_signal_1676 ), .Q ( new_AGEMA_signal_5041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C ( clk ), .D ( new_AGEMA_signal_5048 ), .Q ( new_AGEMA_signal_5049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C ( clk ), .D ( new_AGEMA_signal_5056 ), .Q ( new_AGEMA_signal_5057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C ( clk ), .D ( new_AGEMA_signal_5064 ), .Q ( new_AGEMA_signal_5065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C ( clk ), .D ( new_AGEMA_signal_5072 ), .Q ( new_AGEMA_signal_5073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C ( clk ), .D ( new_AGEMA_signal_5082 ), .Q ( new_AGEMA_signal_5083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C ( clk ), .D ( new_AGEMA_signal_5092 ), .Q ( new_AGEMA_signal_5093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C ( clk ), .D ( new_AGEMA_signal_5100 ), .Q ( new_AGEMA_signal_5101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C ( clk ), .D ( new_AGEMA_signal_5108 ), .Q ( new_AGEMA_signal_5109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C ( clk ), .D ( new_AGEMA_signal_5114 ), .Q ( new_AGEMA_signal_5115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C ( clk ), .D ( new_AGEMA_signal_5120 ), .Q ( new_AGEMA_signal_5121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C ( clk ), .D ( n2276 ), .Q ( new_AGEMA_signal_5125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C ( clk ), .D ( new_AGEMA_signal_1692 ), .Q ( new_AGEMA_signal_5129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C ( clk ), .D ( new_AGEMA_signal_5134 ), .Q ( new_AGEMA_signal_5135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C ( clk ), .D ( new_AGEMA_signal_5140 ), .Q ( new_AGEMA_signal_5141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C ( clk ), .D ( new_AGEMA_signal_5148 ), .Q ( new_AGEMA_signal_5149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C ( clk ), .D ( new_AGEMA_signal_5156 ), .Q ( new_AGEMA_signal_5157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C ( clk ), .D ( new_AGEMA_signal_5162 ), .Q ( new_AGEMA_signal_5163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C ( clk ), .D ( new_AGEMA_signal_5168 ), .Q ( new_AGEMA_signal_5169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C ( clk ), .D ( new_AGEMA_signal_5180 ), .Q ( new_AGEMA_signal_5181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C ( clk ), .D ( new_AGEMA_signal_5188 ), .Q ( new_AGEMA_signal_5189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C ( clk ), .D ( n2622 ), .Q ( new_AGEMA_signal_5193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C ( clk ), .D ( new_AGEMA_signal_1715 ), .Q ( new_AGEMA_signal_5197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C ( clk ), .D ( new_AGEMA_signal_5202 ), .Q ( new_AGEMA_signal_5203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C ( clk ), .D ( new_AGEMA_signal_5208 ), .Q ( new_AGEMA_signal_5209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C ( clk ), .D ( new_AGEMA_signal_5214 ), .Q ( new_AGEMA_signal_5215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C ( clk ), .D ( new_AGEMA_signal_5220 ), .Q ( new_AGEMA_signal_5221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C ( clk ), .D ( n2804 ), .Q ( new_AGEMA_signal_5225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C ( clk ), .D ( new_AGEMA_signal_1722 ), .Q ( new_AGEMA_signal_5229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C ( clk ), .D ( n1990 ), .Q ( new_AGEMA_signal_5233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C ( clk ), .D ( new_AGEMA_signal_1590 ), .Q ( new_AGEMA_signal_5239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C ( clk ), .D ( n2078 ), .Q ( new_AGEMA_signal_5253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C ( clk ), .D ( new_AGEMA_signal_1678 ), .Q ( new_AGEMA_signal_5259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C ( clk ), .D ( new_AGEMA_signal_5268 ), .Q ( new_AGEMA_signal_5269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C ( clk ), .D ( new_AGEMA_signal_5278 ), .Q ( new_AGEMA_signal_5279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C ( clk ), .D ( n2128 ), .Q ( new_AGEMA_signal_5285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C ( clk ), .D ( new_AGEMA_signal_1735 ), .Q ( new_AGEMA_signal_5291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C ( clk ), .D ( n2148 ), .Q ( new_AGEMA_signal_5297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_5303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C ( clk ), .D ( new_AGEMA_signal_5326 ), .Q ( new_AGEMA_signal_5327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C ( clk ), .D ( new_AGEMA_signal_5334 ), .Q ( new_AGEMA_signal_5335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C ( clk ), .D ( n2306 ), .Q ( new_AGEMA_signal_5341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C ( clk ), .D ( new_AGEMA_signal_1621 ), .Q ( new_AGEMA_signal_5347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C ( clk ), .D ( new_AGEMA_signal_5354 ), .Q ( new_AGEMA_signal_5355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C ( clk ), .D ( new_AGEMA_signal_5362 ), .Q ( new_AGEMA_signal_5363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C ( clk ), .D ( new_AGEMA_signal_5370 ), .Q ( new_AGEMA_signal_5371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C ( clk ), .D ( new_AGEMA_signal_5378 ), .Q ( new_AGEMA_signal_5379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C ( clk ), .D ( new_AGEMA_signal_5406 ), .Q ( new_AGEMA_signal_5407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C ( clk ), .D ( new_AGEMA_signal_5414 ), .Q ( new_AGEMA_signal_5415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C ( clk ), .D ( n1999 ), .Q ( new_AGEMA_signal_5429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C ( clk ), .D ( new_AGEMA_signal_1671 ), .Q ( new_AGEMA_signal_5437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C ( clk ), .D ( new_AGEMA_signal_5448 ), .Q ( new_AGEMA_signal_5449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C ( clk ), .D ( new_AGEMA_signal_5460 ), .Q ( new_AGEMA_signal_5461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C ( clk ), .D ( new_AGEMA_signal_5474 ), .Q ( new_AGEMA_signal_5475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C ( clk ), .D ( new_AGEMA_signal_5488 ), .Q ( new_AGEMA_signal_5489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C ( clk ), .D ( n2205 ), .Q ( new_AGEMA_signal_5497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C ( clk ), .D ( new_AGEMA_signal_1741 ), .Q ( new_AGEMA_signal_5505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C ( clk ), .D ( new_AGEMA_signal_5518 ), .Q ( new_AGEMA_signal_5519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C ( clk ), .D ( new_AGEMA_signal_5532 ), .Q ( new_AGEMA_signal_5533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C ( clk ), .D ( n2516 ), .Q ( new_AGEMA_signal_5541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C ( clk ), .D ( new_AGEMA_signal_1704 ), .Q ( new_AGEMA_signal_5549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C ( clk ), .D ( n2808 ), .Q ( new_AGEMA_signal_5557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C ( clk ), .D ( new_AGEMA_signal_1719 ), .Q ( new_AGEMA_signal_5565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C ( clk ), .D ( new_AGEMA_signal_5590 ), .Q ( new_AGEMA_signal_5591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C ( clk ), .D ( new_AGEMA_signal_5606 ), .Q ( new_AGEMA_signal_5607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C ( clk ), .D ( new_AGEMA_signal_5634 ), .Q ( new_AGEMA_signal_5635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C ( clk ), .D ( new_AGEMA_signal_5650 ), .Q ( new_AGEMA_signal_5651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C ( clk ), .D ( n2527 ), .Q ( new_AGEMA_signal_5661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C ( clk ), .D ( new_AGEMA_signal_1758 ), .Q ( new_AGEMA_signal_5671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C ( clk ), .D ( new_AGEMA_signal_5732 ), .Q ( new_AGEMA_signal_5733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C ( clk ), .D ( new_AGEMA_signal_5748 ), .Q ( new_AGEMA_signal_5749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C ( clk ), .D ( new_AGEMA_signal_5786 ), .Q ( new_AGEMA_signal_5787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C ( clk ), .D ( new_AGEMA_signal_5804 ), .Q ( new_AGEMA_signal_5805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C ( clk ), .D ( new_AGEMA_signal_5886 ), .Q ( new_AGEMA_signal_5887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C ( clk ), .D ( new_AGEMA_signal_5906 ), .Q ( new_AGEMA_signal_5907 ) ) ;

    /* cells in depth 14 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2002 ( .a ({new_AGEMA_signal_4296, new_AGEMA_signal_4294}), .b ({new_AGEMA_signal_1667, n1933}), .clk ( clk ), .r ( Fresh[723] ), .c ({new_AGEMA_signal_1726, n1935}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2054 ( .a ({new_AGEMA_signal_1668, n1958}), .b ({new_AGEMA_signal_4312, new_AGEMA_signal_4304}), .clk ( clk ), .r ( Fresh[724] ), .c ({new_AGEMA_signal_1727, n1959}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2109 ( .a ({new_AGEMA_signal_1670, n1982}), .b ({new_AGEMA_signal_4316, new_AGEMA_signal_4314}), .clk ( clk ), .r ( Fresh[725] ), .c ({new_AGEMA_signal_1728, n1983}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2149 ( .a ({new_AGEMA_signal_4324, new_AGEMA_signal_4320}), .b ({new_AGEMA_signal_1672, n2011}), .clk ( clk ), .r ( Fresh[726] ), .c ({new_AGEMA_signal_1729, n2014}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2166 ( .a ({new_AGEMA_signal_4340, new_AGEMA_signal_4332}), .b ({new_AGEMA_signal_1596, n2025}), .clk ( clk ), .r ( Fresh[727] ), .c ({new_AGEMA_signal_1673, n2029}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2180 ( .a ({new_AGEMA_signal_4344, new_AGEMA_signal_4342}), .b ({new_AGEMA_signal_1674, n2036}), .clk ( clk ), .r ( Fresh[728] ), .c ({new_AGEMA_signal_1731, n2037}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2197 ( .a ({new_AGEMA_signal_4356, new_AGEMA_signal_4350}), .b ({new_AGEMA_signal_1675, n2049}), .clk ( clk ), .r ( Fresh[729] ), .c ({new_AGEMA_signal_1732, n2052}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2219 ( .a ({new_AGEMA_signal_1677, n2067}), .b ({new_AGEMA_signal_4364, new_AGEMA_signal_4360}), .clk ( clk ), .r ( Fresh[730] ), .c ({new_AGEMA_signal_1733, n2070}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2258 ( .a ({new_AGEMA_signal_1679, n2097}), .b ({new_AGEMA_signal_1680, n2096}), .clk ( clk ), .r ( Fresh[731] ), .c ({new_AGEMA_signal_1734, n2098}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2287 ( .a ({new_AGEMA_signal_1682, n2124}), .b ({new_AGEMA_signal_4380, new_AGEMA_signal_4372}), .clk ( clk ), .r ( Fresh[732] ), .c ({new_AGEMA_signal_1736, n2125}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2311 ( .a ({new_AGEMA_signal_4388, new_AGEMA_signal_4384}), .b ({new_AGEMA_signal_1683, n2142}), .clk ( clk ), .r ( Fresh[733] ), .c ({new_AGEMA_signal_1737, n2145}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2333 ( .a ({new_AGEMA_signal_1684, n2168}), .b ({new_AGEMA_signal_1685, n2167}), .clk ( clk ), .r ( Fresh[734] ), .c ({new_AGEMA_signal_1738, n2169}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2350 ( .a ({new_AGEMA_signal_1686, n2184}), .b ({new_AGEMA_signal_4400, new_AGEMA_signal_4394}), .clk ( clk ), .r ( Fresh[735] ), .c ({new_AGEMA_signal_1739, n2185}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2365 ( .a ({new_AGEMA_signal_1687, n2197}), .b ({new_AGEMA_signal_4412, new_AGEMA_signal_4406}), .clk ( clk ), .r ( Fresh[736] ), .c ({new_AGEMA_signal_1740, n2198}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2396 ( .a ({new_AGEMA_signal_1689, n2232}), .b ({new_AGEMA_signal_1615, n2231}), .clk ( clk ), .r ( Fresh[737] ), .c ({new_AGEMA_signal_1742, n2312}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2404 ( .a ({new_AGEMA_signal_1743, n2239}), .b ({new_AGEMA_signal_4424, new_AGEMA_signal_4418}), .clk ( clk ), .r ( Fresh[738] ), .c ({new_AGEMA_signal_1781, n2258}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2415 ( .a ({new_AGEMA_signal_1691, n2250}), .b ({new_AGEMA_signal_4436, new_AGEMA_signal_4430}), .clk ( clk ), .r ( Fresh[739] ), .c ({new_AGEMA_signal_1744, n2251}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2440 ( .a ({new_AGEMA_signal_4448, new_AGEMA_signal_4442}), .b ({new_AGEMA_signal_1693, n2272}), .clk ( clk ), .r ( Fresh[740] ), .c ({new_AGEMA_signal_1745, n2274}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2469 ( .a ({new_AGEMA_signal_4456, new_AGEMA_signal_4452}), .b ({new_AGEMA_signal_1694, n2296}), .clk ( clk ), .r ( Fresh[741] ), .c ({new_AGEMA_signal_1746, n2302}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2490 ( .a ({new_AGEMA_signal_1695, n2324}), .b ({new_AGEMA_signal_4472, new_AGEMA_signal_4464}), .clk ( clk ), .r ( Fresh[742] ), .c ({new_AGEMA_signal_1747, n2339}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2503 ( .a ({new_AGEMA_signal_1696, n2337}), .b ({new_AGEMA_signal_4480, new_AGEMA_signal_4476}), .clk ( clk ), .r ( Fresh[743] ), .c ({new_AGEMA_signal_1748, n2338}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2515 ( .a ({new_AGEMA_signal_1697, n2350}), .b ({new_AGEMA_signal_4492, new_AGEMA_signal_4486}), .clk ( clk ), .r ( Fresh[744] ), .c ({new_AGEMA_signal_1749, n2351}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2529 ( .a ({new_AGEMA_signal_4508, new_AGEMA_signal_4500}), .b ({new_AGEMA_signal_1698, n2362}), .clk ( clk ), .r ( Fresh[745] ), .c ({new_AGEMA_signal_1750, n2365}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2551 ( .a ({new_AGEMA_signal_1629, n2389}), .b ({new_AGEMA_signal_4512, new_AGEMA_signal_4510}), .clk ( clk ), .r ( Fresh[746] ), .c ({new_AGEMA_signal_1699, n2399}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2560 ( .a ({new_AGEMA_signal_1700, n2397}), .b ({new_AGEMA_signal_4524, new_AGEMA_signal_4518}), .clk ( clk ), .r ( Fresh[747] ), .c ({new_AGEMA_signal_1751, n2398}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2572 ( .a ({new_AGEMA_signal_1631, n2411}), .b ({new_AGEMA_signal_4528, new_AGEMA_signal_4526}), .clk ( clk ), .r ( Fresh[748] ), .c ({new_AGEMA_signal_1701, n2423}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2581 ( .a ({new_AGEMA_signal_4532, new_AGEMA_signal_4530}), .b ({new_AGEMA_signal_1634, n2420}), .clk ( clk ), .r ( Fresh[749] ), .c ({new_AGEMA_signal_1702, n2422}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2596 ( .a ({new_AGEMA_signal_1703, n2440}), .b ({new_AGEMA_signal_4544, new_AGEMA_signal_4538}), .clk ( clk ), .r ( Fresh[750] ), .c ({new_AGEMA_signal_1753, n2441}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2623 ( .a ({new_AGEMA_signal_1639, n2471}), .b ({new_AGEMA_signal_4556, new_AGEMA_signal_4550}), .clk ( clk ), .r ( Fresh[751] ), .c ({new_AGEMA_signal_1705, n2479}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2637 ( .a ({new_AGEMA_signal_1706, n2485}), .b ({new_AGEMA_signal_4572, new_AGEMA_signal_4564}), .clk ( clk ), .r ( Fresh[752] ), .c ({new_AGEMA_signal_1755, n2512}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2652 ( .a ({new_AGEMA_signal_1641, n2502}), .b ({new_AGEMA_signal_1707, n2501}), .clk ( clk ), .r ( Fresh[753] ), .c ({new_AGEMA_signal_1756, n2510}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2686 ( .a ({new_AGEMA_signal_1710, n2550}), .b ({new_AGEMA_signal_1711, n2549}), .clk ( clk ), .r ( Fresh[754] ), .c ({new_AGEMA_signal_1759, n2552}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2702 ( .a ({new_AGEMA_signal_4588, new_AGEMA_signal_4580}), .b ({new_AGEMA_signal_1712, n2569}), .clk ( clk ), .r ( Fresh[755] ), .c ({new_AGEMA_signal_1760, n2593}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2713 ( .a ({new_AGEMA_signal_4600, new_AGEMA_signal_4594}), .b ({new_AGEMA_signal_1713, n2584}), .clk ( clk ), .r ( Fresh[756] ), .c ({new_AGEMA_signal_1761, n2589}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2730 ( .a ({new_AGEMA_signal_4612, new_AGEMA_signal_4606}), .b ({new_AGEMA_signal_1650, n2606}), .clk ( clk ), .r ( Fresh[757] ), .c ({new_AGEMA_signal_1714, n2608}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2748 ( .a ({new_AGEMA_signal_4616, new_AGEMA_signal_4614}), .b ({new_AGEMA_signal_1716, n2634}), .clk ( clk ), .r ( Fresh[758] ), .c ({new_AGEMA_signal_1763, n2636}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2762 ( .a ({new_AGEMA_signal_4624, new_AGEMA_signal_4620}), .b ({new_AGEMA_signal_1717, n2657}), .clk ( clk ), .r ( Fresh[759] ), .c ({new_AGEMA_signal_1764, n2659}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2784 ( .a ({new_AGEMA_signal_4632, new_AGEMA_signal_4628}), .b ({new_AGEMA_signal_1718, n2697}), .clk ( clk ), .r ( Fresh[760] ), .c ({new_AGEMA_signal_1765, n2702}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2811 ( .a ({new_AGEMA_signal_1720, n2747}), .b ({new_AGEMA_signal_1721, n2746}), .clk ( clk ), .r ( Fresh[761] ), .c ({new_AGEMA_signal_1766, n2806}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2839 ( .a ({new_AGEMA_signal_4640, new_AGEMA_signal_4636}), .b ({new_AGEMA_signal_1665, n2799}), .clk ( clk ), .r ( Fresh[762] ), .c ({new_AGEMA_signal_1724, n2801}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2853 ( .a ({new_AGEMA_signal_4644, new_AGEMA_signal_4642}), .b ({new_AGEMA_signal_1725, n2827}), .clk ( clk ), .r ( Fresh[763] ), .c ({new_AGEMA_signal_1768, n2829}) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C ( clk ), .D ( new_AGEMA_signal_4649 ), .Q ( new_AGEMA_signal_4650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C ( clk ), .D ( new_AGEMA_signal_4655 ), .Q ( new_AGEMA_signal_4656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C ( clk ), .D ( new_AGEMA_signal_4657 ), .Q ( new_AGEMA_signal_4658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C ( clk ), .D ( new_AGEMA_signal_4659 ), .Q ( new_AGEMA_signal_4660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C ( clk ), .D ( new_AGEMA_signal_4663 ), .Q ( new_AGEMA_signal_4664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C ( clk ), .D ( new_AGEMA_signal_4667 ), .Q ( new_AGEMA_signal_4668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C ( clk ), .D ( new_AGEMA_signal_4675 ), .Q ( new_AGEMA_signal_4676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C ( clk ), .D ( new_AGEMA_signal_4683 ), .Q ( new_AGEMA_signal_4684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C ( clk ), .D ( new_AGEMA_signal_4691 ), .Q ( new_AGEMA_signal_4692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C ( clk ), .D ( new_AGEMA_signal_4699 ), .Q ( new_AGEMA_signal_4700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C ( clk ), .D ( new_AGEMA_signal_4707 ), .Q ( new_AGEMA_signal_4708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C ( clk ), .D ( new_AGEMA_signal_4715 ), .Q ( new_AGEMA_signal_4716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C ( clk ), .D ( new_AGEMA_signal_4723 ), .Q ( new_AGEMA_signal_4724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C ( clk ), .D ( new_AGEMA_signal_4731 ), .Q ( new_AGEMA_signal_4732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C ( clk ), .D ( new_AGEMA_signal_4737 ), .Q ( new_AGEMA_signal_4738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C ( clk ), .D ( new_AGEMA_signal_4743 ), .Q ( new_AGEMA_signal_4744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C ( clk ), .D ( new_AGEMA_signal_4753 ), .Q ( new_AGEMA_signal_4754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C ( clk ), .D ( new_AGEMA_signal_4763 ), .Q ( new_AGEMA_signal_4764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C ( clk ), .D ( new_AGEMA_signal_4771 ), .Q ( new_AGEMA_signal_4772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C ( clk ), .D ( new_AGEMA_signal_4779 ), .Q ( new_AGEMA_signal_4780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C ( clk ), .D ( new_AGEMA_signal_4787 ), .Q ( new_AGEMA_signal_4788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C ( clk ), .D ( new_AGEMA_signal_4795 ), .Q ( new_AGEMA_signal_4796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C ( clk ), .D ( new_AGEMA_signal_4803 ), .Q ( new_AGEMA_signal_4804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C ( clk ), .D ( new_AGEMA_signal_4811 ), .Q ( new_AGEMA_signal_4812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C ( clk ), .D ( new_AGEMA_signal_4813 ), .Q ( new_AGEMA_signal_4814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C ( clk ), .D ( new_AGEMA_signal_4815 ), .Q ( new_AGEMA_signal_4816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C ( clk ), .D ( new_AGEMA_signal_4819 ), .Q ( new_AGEMA_signal_4820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C ( clk ), .D ( new_AGEMA_signal_4823 ), .Q ( new_AGEMA_signal_4824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C ( clk ), .D ( new_AGEMA_signal_4829 ), .Q ( new_AGEMA_signal_4830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C ( clk ), .D ( new_AGEMA_signal_4835 ), .Q ( new_AGEMA_signal_4836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C ( clk ), .D ( new_AGEMA_signal_4839 ), .Q ( new_AGEMA_signal_4840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C ( clk ), .D ( new_AGEMA_signal_4843 ), .Q ( new_AGEMA_signal_4844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C ( clk ), .D ( new_AGEMA_signal_4853 ), .Q ( new_AGEMA_signal_4854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C ( clk ), .D ( new_AGEMA_signal_4863 ), .Q ( new_AGEMA_signal_4864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C ( clk ), .D ( new_AGEMA_signal_4871 ), .Q ( new_AGEMA_signal_4872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C ( clk ), .D ( new_AGEMA_signal_4879 ), .Q ( new_AGEMA_signal_4880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C ( clk ), .D ( new_AGEMA_signal_4883 ), .Q ( new_AGEMA_signal_4884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C ( clk ), .D ( new_AGEMA_signal_4887 ), .Q ( new_AGEMA_signal_4888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C ( clk ), .D ( new_AGEMA_signal_4889 ), .Q ( new_AGEMA_signal_4890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C ( clk ), .D ( new_AGEMA_signal_4891 ), .Q ( new_AGEMA_signal_4892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C ( clk ), .D ( new_AGEMA_signal_4899 ), .Q ( new_AGEMA_signal_4900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C ( clk ), .D ( new_AGEMA_signal_4907 ), .Q ( new_AGEMA_signal_4908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C ( clk ), .D ( new_AGEMA_signal_4915 ), .Q ( new_AGEMA_signal_4916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C ( clk ), .D ( new_AGEMA_signal_4923 ), .Q ( new_AGEMA_signal_4924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C ( clk ), .D ( new_AGEMA_signal_4929 ), .Q ( new_AGEMA_signal_4930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C ( clk ), .D ( new_AGEMA_signal_4935 ), .Q ( new_AGEMA_signal_4936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C ( clk ), .D ( new_AGEMA_signal_4939 ), .Q ( new_AGEMA_signal_4940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C ( clk ), .D ( new_AGEMA_signal_4943 ), .Q ( new_AGEMA_signal_4944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C ( clk ), .D ( new_AGEMA_signal_4951 ), .Q ( new_AGEMA_signal_4952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C ( clk ), .D ( new_AGEMA_signal_4959 ), .Q ( new_AGEMA_signal_4960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C ( clk ), .D ( new_AGEMA_signal_4961 ), .Q ( new_AGEMA_signal_4962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C ( clk ), .D ( new_AGEMA_signal_4963 ), .Q ( new_AGEMA_signal_4964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C ( clk ), .D ( new_AGEMA_signal_4967 ), .Q ( new_AGEMA_signal_4968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C ( clk ), .D ( new_AGEMA_signal_4973 ), .Q ( new_AGEMA_signal_4974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C ( clk ), .D ( new_AGEMA_signal_4979 ), .Q ( new_AGEMA_signal_4980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C ( clk ), .D ( new_AGEMA_signal_4985 ), .Q ( new_AGEMA_signal_4986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C ( clk ), .D ( new_AGEMA_signal_4991 ), .Q ( new_AGEMA_signal_4992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C ( clk ), .D ( new_AGEMA_signal_4997 ), .Q ( new_AGEMA_signal_4998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C ( clk ), .D ( new_AGEMA_signal_5001 ), .Q ( new_AGEMA_signal_5002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C ( clk ), .D ( new_AGEMA_signal_5005 ), .Q ( new_AGEMA_signal_5006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C ( clk ), .D ( new_AGEMA_signal_5013 ), .Q ( new_AGEMA_signal_5014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C ( clk ), .D ( new_AGEMA_signal_5021 ), .Q ( new_AGEMA_signal_5022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C ( clk ), .D ( new_AGEMA_signal_5027 ), .Q ( new_AGEMA_signal_5028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C ( clk ), .D ( new_AGEMA_signal_5033 ), .Q ( new_AGEMA_signal_5034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C ( clk ), .D ( new_AGEMA_signal_5037 ), .Q ( new_AGEMA_signal_5038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C ( clk ), .D ( new_AGEMA_signal_5041 ), .Q ( new_AGEMA_signal_5042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C ( clk ), .D ( new_AGEMA_signal_5049 ), .Q ( new_AGEMA_signal_5050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C ( clk ), .D ( new_AGEMA_signal_5057 ), .Q ( new_AGEMA_signal_5058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C ( clk ), .D ( new_AGEMA_signal_5065 ), .Q ( new_AGEMA_signal_5066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C ( clk ), .D ( new_AGEMA_signal_5073 ), .Q ( new_AGEMA_signal_5074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C ( clk ), .D ( new_AGEMA_signal_5083 ), .Q ( new_AGEMA_signal_5084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C ( clk ), .D ( new_AGEMA_signal_5093 ), .Q ( new_AGEMA_signal_5094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C ( clk ), .D ( new_AGEMA_signal_5101 ), .Q ( new_AGEMA_signal_5102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C ( clk ), .D ( new_AGEMA_signal_5109 ), .Q ( new_AGEMA_signal_5110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C ( clk ), .D ( new_AGEMA_signal_5115 ), .Q ( new_AGEMA_signal_5116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C ( clk ), .D ( new_AGEMA_signal_5121 ), .Q ( new_AGEMA_signal_5122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C ( clk ), .D ( new_AGEMA_signal_5125 ), .Q ( new_AGEMA_signal_5126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C ( clk ), .D ( new_AGEMA_signal_5129 ), .Q ( new_AGEMA_signal_5130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C ( clk ), .D ( new_AGEMA_signal_5135 ), .Q ( new_AGEMA_signal_5136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C ( clk ), .D ( new_AGEMA_signal_5141 ), .Q ( new_AGEMA_signal_5142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C ( clk ), .D ( new_AGEMA_signal_5149 ), .Q ( new_AGEMA_signal_5150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C ( clk ), .D ( new_AGEMA_signal_5157 ), .Q ( new_AGEMA_signal_5158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C ( clk ), .D ( new_AGEMA_signal_5163 ), .Q ( new_AGEMA_signal_5164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C ( clk ), .D ( new_AGEMA_signal_5169 ), .Q ( new_AGEMA_signal_5170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C ( clk ), .D ( new_AGEMA_signal_5181 ), .Q ( new_AGEMA_signal_5182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C ( clk ), .D ( new_AGEMA_signal_5189 ), .Q ( new_AGEMA_signal_5190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C ( clk ), .D ( new_AGEMA_signal_5193 ), .Q ( new_AGEMA_signal_5194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C ( clk ), .D ( new_AGEMA_signal_5197 ), .Q ( new_AGEMA_signal_5198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C ( clk ), .D ( new_AGEMA_signal_5203 ), .Q ( new_AGEMA_signal_5204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C ( clk ), .D ( new_AGEMA_signal_5209 ), .Q ( new_AGEMA_signal_5210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C ( clk ), .D ( new_AGEMA_signal_5215 ), .Q ( new_AGEMA_signal_5216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C ( clk ), .D ( new_AGEMA_signal_5221 ), .Q ( new_AGEMA_signal_5222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C ( clk ), .D ( new_AGEMA_signal_5225 ), .Q ( new_AGEMA_signal_5226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C ( clk ), .D ( new_AGEMA_signal_5229 ), .Q ( new_AGEMA_signal_5230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C ( clk ), .D ( new_AGEMA_signal_5233 ), .Q ( new_AGEMA_signal_5234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C ( clk ), .D ( new_AGEMA_signal_5239 ), .Q ( new_AGEMA_signal_5240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C ( clk ), .D ( new_AGEMA_signal_5253 ), .Q ( new_AGEMA_signal_5254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C ( clk ), .D ( new_AGEMA_signal_5259 ), .Q ( new_AGEMA_signal_5260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C ( clk ), .D ( new_AGEMA_signal_5269 ), .Q ( new_AGEMA_signal_5270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C ( clk ), .D ( new_AGEMA_signal_5279 ), .Q ( new_AGEMA_signal_5280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C ( clk ), .D ( new_AGEMA_signal_5285 ), .Q ( new_AGEMA_signal_5286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C ( clk ), .D ( new_AGEMA_signal_5291 ), .Q ( new_AGEMA_signal_5292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C ( clk ), .D ( new_AGEMA_signal_5297 ), .Q ( new_AGEMA_signal_5298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C ( clk ), .D ( new_AGEMA_signal_5303 ), .Q ( new_AGEMA_signal_5304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C ( clk ), .D ( new_AGEMA_signal_5327 ), .Q ( new_AGEMA_signal_5328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C ( clk ), .D ( new_AGEMA_signal_5335 ), .Q ( new_AGEMA_signal_5336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C ( clk ), .D ( new_AGEMA_signal_5341 ), .Q ( new_AGEMA_signal_5342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C ( clk ), .D ( new_AGEMA_signal_5347 ), .Q ( new_AGEMA_signal_5348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C ( clk ), .D ( new_AGEMA_signal_5355 ), .Q ( new_AGEMA_signal_5356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C ( clk ), .D ( new_AGEMA_signal_5363 ), .Q ( new_AGEMA_signal_5364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C ( clk ), .D ( new_AGEMA_signal_5371 ), .Q ( new_AGEMA_signal_5372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C ( clk ), .D ( new_AGEMA_signal_5379 ), .Q ( new_AGEMA_signal_5380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C ( clk ), .D ( new_AGEMA_signal_5407 ), .Q ( new_AGEMA_signal_5408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C ( clk ), .D ( new_AGEMA_signal_5415 ), .Q ( new_AGEMA_signal_5416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C ( clk ), .D ( new_AGEMA_signal_5429 ), .Q ( new_AGEMA_signal_5430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C ( clk ), .D ( new_AGEMA_signal_5437 ), .Q ( new_AGEMA_signal_5438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C ( clk ), .D ( new_AGEMA_signal_5449 ), .Q ( new_AGEMA_signal_5450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C ( clk ), .D ( new_AGEMA_signal_5461 ), .Q ( new_AGEMA_signal_5462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C ( clk ), .D ( new_AGEMA_signal_5475 ), .Q ( new_AGEMA_signal_5476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C ( clk ), .D ( new_AGEMA_signal_5489 ), .Q ( new_AGEMA_signal_5490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C ( clk ), .D ( new_AGEMA_signal_5497 ), .Q ( new_AGEMA_signal_5498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C ( clk ), .D ( new_AGEMA_signal_5505 ), .Q ( new_AGEMA_signal_5506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C ( clk ), .D ( new_AGEMA_signal_5519 ), .Q ( new_AGEMA_signal_5520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C ( clk ), .D ( new_AGEMA_signal_5533 ), .Q ( new_AGEMA_signal_5534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C ( clk ), .D ( new_AGEMA_signal_5541 ), .Q ( new_AGEMA_signal_5542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C ( clk ), .D ( new_AGEMA_signal_5549 ), .Q ( new_AGEMA_signal_5550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C ( clk ), .D ( new_AGEMA_signal_5557 ), .Q ( new_AGEMA_signal_5558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C ( clk ), .D ( new_AGEMA_signal_5565 ), .Q ( new_AGEMA_signal_5566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C ( clk ), .D ( new_AGEMA_signal_5591 ), .Q ( new_AGEMA_signal_5592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C ( clk ), .D ( new_AGEMA_signal_5607 ), .Q ( new_AGEMA_signal_5608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C ( clk ), .D ( new_AGEMA_signal_5635 ), .Q ( new_AGEMA_signal_5636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C ( clk ), .D ( new_AGEMA_signal_5651 ), .Q ( new_AGEMA_signal_5652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C ( clk ), .D ( new_AGEMA_signal_5661 ), .Q ( new_AGEMA_signal_5662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C ( clk ), .D ( new_AGEMA_signal_5671 ), .Q ( new_AGEMA_signal_5672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C ( clk ), .D ( new_AGEMA_signal_5733 ), .Q ( new_AGEMA_signal_5734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C ( clk ), .D ( new_AGEMA_signal_5749 ), .Q ( new_AGEMA_signal_5750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C ( clk ), .D ( new_AGEMA_signal_5787 ), .Q ( new_AGEMA_signal_5788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C ( clk ), .D ( new_AGEMA_signal_5805 ), .Q ( new_AGEMA_signal_5806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C ( clk ), .D ( new_AGEMA_signal_5887 ), .Q ( new_AGEMA_signal_5888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C ( clk ), .D ( new_AGEMA_signal_5907 ), .Q ( new_AGEMA_signal_5908 ) ) ;

    /* cells in depth 15 */
    buf_clk new_AGEMA_reg_buffer_3151 ( .C ( clk ), .D ( new_AGEMA_signal_4968 ), .Q ( new_AGEMA_signal_4969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C ( clk ), .D ( new_AGEMA_signal_4974 ), .Q ( new_AGEMA_signal_4975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C ( clk ), .D ( new_AGEMA_signal_4980 ), .Q ( new_AGEMA_signal_4981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C ( clk ), .D ( new_AGEMA_signal_4986 ), .Q ( new_AGEMA_signal_4987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C ( clk ), .D ( new_AGEMA_signal_4992 ), .Q ( new_AGEMA_signal_4993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C ( clk ), .D ( new_AGEMA_signal_4998 ), .Q ( new_AGEMA_signal_4999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C ( clk ), .D ( new_AGEMA_signal_5002 ), .Q ( new_AGEMA_signal_5003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C ( clk ), .D ( new_AGEMA_signal_5006 ), .Q ( new_AGEMA_signal_5007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C ( clk ), .D ( new_AGEMA_signal_5014 ), .Q ( new_AGEMA_signal_5015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C ( clk ), .D ( new_AGEMA_signal_5022 ), .Q ( new_AGEMA_signal_5023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C ( clk ), .D ( new_AGEMA_signal_5028 ), .Q ( new_AGEMA_signal_5029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C ( clk ), .D ( new_AGEMA_signal_5034 ), .Q ( new_AGEMA_signal_5035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C ( clk ), .D ( new_AGEMA_signal_5038 ), .Q ( new_AGEMA_signal_5039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C ( clk ), .D ( new_AGEMA_signal_5042 ), .Q ( new_AGEMA_signal_5043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C ( clk ), .D ( new_AGEMA_signal_5050 ), .Q ( new_AGEMA_signal_5051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C ( clk ), .D ( new_AGEMA_signal_5058 ), .Q ( new_AGEMA_signal_5059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C ( clk ), .D ( new_AGEMA_signal_5066 ), .Q ( new_AGEMA_signal_5067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C ( clk ), .D ( new_AGEMA_signal_5074 ), .Q ( new_AGEMA_signal_5075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C ( clk ), .D ( new_AGEMA_signal_5084 ), .Q ( new_AGEMA_signal_5085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C ( clk ), .D ( new_AGEMA_signal_5094 ), .Q ( new_AGEMA_signal_5095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C ( clk ), .D ( new_AGEMA_signal_5102 ), .Q ( new_AGEMA_signal_5103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C ( clk ), .D ( new_AGEMA_signal_5110 ), .Q ( new_AGEMA_signal_5111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C ( clk ), .D ( new_AGEMA_signal_5116 ), .Q ( new_AGEMA_signal_5117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C ( clk ), .D ( new_AGEMA_signal_5122 ), .Q ( new_AGEMA_signal_5123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C ( clk ), .D ( new_AGEMA_signal_5126 ), .Q ( new_AGEMA_signal_5127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C ( clk ), .D ( new_AGEMA_signal_5130 ), .Q ( new_AGEMA_signal_5131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C ( clk ), .D ( new_AGEMA_signal_5136 ), .Q ( new_AGEMA_signal_5137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C ( clk ), .D ( new_AGEMA_signal_5142 ), .Q ( new_AGEMA_signal_5143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C ( clk ), .D ( new_AGEMA_signal_5150 ), .Q ( new_AGEMA_signal_5151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C ( clk ), .D ( new_AGEMA_signal_5158 ), .Q ( new_AGEMA_signal_5159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C ( clk ), .D ( new_AGEMA_signal_5164 ), .Q ( new_AGEMA_signal_5165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C ( clk ), .D ( new_AGEMA_signal_5170 ), .Q ( new_AGEMA_signal_5171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C ( clk ), .D ( n2512 ), .Q ( new_AGEMA_signal_5173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C ( clk ), .D ( new_AGEMA_signal_1755 ), .Q ( new_AGEMA_signal_5175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C ( clk ), .D ( new_AGEMA_signal_5182 ), .Q ( new_AGEMA_signal_5183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C ( clk ), .D ( new_AGEMA_signal_5190 ), .Q ( new_AGEMA_signal_5191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C ( clk ), .D ( new_AGEMA_signal_5194 ), .Q ( new_AGEMA_signal_5195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C ( clk ), .D ( new_AGEMA_signal_5198 ), .Q ( new_AGEMA_signal_5199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C ( clk ), .D ( new_AGEMA_signal_5204 ), .Q ( new_AGEMA_signal_5205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C ( clk ), .D ( new_AGEMA_signal_5210 ), .Q ( new_AGEMA_signal_5211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C ( clk ), .D ( new_AGEMA_signal_5216 ), .Q ( new_AGEMA_signal_5217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C ( clk ), .D ( new_AGEMA_signal_5222 ), .Q ( new_AGEMA_signal_5223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C ( clk ), .D ( new_AGEMA_signal_5226 ), .Q ( new_AGEMA_signal_5227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C ( clk ), .D ( new_AGEMA_signal_5230 ), .Q ( new_AGEMA_signal_5231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C ( clk ), .D ( new_AGEMA_signal_5234 ), .Q ( new_AGEMA_signal_5235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C ( clk ), .D ( new_AGEMA_signal_5240 ), .Q ( new_AGEMA_signal_5241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C ( clk ), .D ( n2037 ), .Q ( new_AGEMA_signal_5245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C ( clk ), .D ( new_AGEMA_signal_1731 ), .Q ( new_AGEMA_signal_5249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C ( clk ), .D ( new_AGEMA_signal_5254 ), .Q ( new_AGEMA_signal_5255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C ( clk ), .D ( new_AGEMA_signal_5260 ), .Q ( new_AGEMA_signal_5261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C ( clk ), .D ( new_AGEMA_signal_5270 ), .Q ( new_AGEMA_signal_5271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C ( clk ), .D ( new_AGEMA_signal_5280 ), .Q ( new_AGEMA_signal_5281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C ( clk ), .D ( new_AGEMA_signal_5286 ), .Q ( new_AGEMA_signal_5287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C ( clk ), .D ( new_AGEMA_signal_5292 ), .Q ( new_AGEMA_signal_5293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C ( clk ), .D ( new_AGEMA_signal_5298 ), .Q ( new_AGEMA_signal_5299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C ( clk ), .D ( new_AGEMA_signal_5304 ), .Q ( new_AGEMA_signal_5305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C ( clk ), .D ( n2198 ), .Q ( new_AGEMA_signal_5309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C ( clk ), .D ( new_AGEMA_signal_1740 ), .Q ( new_AGEMA_signal_5313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C ( clk ), .D ( n2258 ), .Q ( new_AGEMA_signal_5317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C ( clk ), .D ( new_AGEMA_signal_1781 ), .Q ( new_AGEMA_signal_5321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C ( clk ), .D ( new_AGEMA_signal_5328 ), .Q ( new_AGEMA_signal_5329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C ( clk ), .D ( new_AGEMA_signal_5336 ), .Q ( new_AGEMA_signal_5337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C ( clk ), .D ( new_AGEMA_signal_5342 ), .Q ( new_AGEMA_signal_5343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C ( clk ), .D ( new_AGEMA_signal_5348 ), .Q ( new_AGEMA_signal_5349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C ( clk ), .D ( new_AGEMA_signal_5356 ), .Q ( new_AGEMA_signal_5357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C ( clk ), .D ( new_AGEMA_signal_5364 ), .Q ( new_AGEMA_signal_5365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C ( clk ), .D ( new_AGEMA_signal_5372 ), .Q ( new_AGEMA_signal_5373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C ( clk ), .D ( new_AGEMA_signal_5380 ), .Q ( new_AGEMA_signal_5381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C ( clk ), .D ( n2593 ), .Q ( new_AGEMA_signal_5389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C ( clk ), .D ( new_AGEMA_signal_1760 ), .Q ( new_AGEMA_signal_5393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C ( clk ), .D ( n2636 ), .Q ( new_AGEMA_signal_5397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_5401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C ( clk ), .D ( new_AGEMA_signal_5408 ), .Q ( new_AGEMA_signal_5409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C ( clk ), .D ( new_AGEMA_signal_5416 ), .Q ( new_AGEMA_signal_5417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C ( clk ), .D ( n2806 ), .Q ( new_AGEMA_signal_5421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_5425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C ( clk ), .D ( new_AGEMA_signal_5430 ), .Q ( new_AGEMA_signal_5431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C ( clk ), .D ( new_AGEMA_signal_5438 ), .Q ( new_AGEMA_signal_5439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C ( clk ), .D ( new_AGEMA_signal_5450 ), .Q ( new_AGEMA_signal_5451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C ( clk ), .D ( new_AGEMA_signal_5462 ), .Q ( new_AGEMA_signal_5463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C ( clk ), .D ( new_AGEMA_signal_5476 ), .Q ( new_AGEMA_signal_5477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C ( clk ), .D ( new_AGEMA_signal_5490 ), .Q ( new_AGEMA_signal_5491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C ( clk ), .D ( new_AGEMA_signal_5498 ), .Q ( new_AGEMA_signal_5499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C ( clk ), .D ( new_AGEMA_signal_5506 ), .Q ( new_AGEMA_signal_5507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C ( clk ), .D ( new_AGEMA_signal_5520 ), .Q ( new_AGEMA_signal_5521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C ( clk ), .D ( new_AGEMA_signal_5534 ), .Q ( new_AGEMA_signal_5535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C ( clk ), .D ( new_AGEMA_signal_5542 ), .Q ( new_AGEMA_signal_5543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C ( clk ), .D ( new_AGEMA_signal_5550 ), .Q ( new_AGEMA_signal_5551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C ( clk ), .D ( new_AGEMA_signal_5558 ), .Q ( new_AGEMA_signal_5559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C ( clk ), .D ( new_AGEMA_signal_5566 ), .Q ( new_AGEMA_signal_5567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C ( clk ), .D ( new_AGEMA_signal_5592 ), .Q ( new_AGEMA_signal_5593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C ( clk ), .D ( new_AGEMA_signal_5608 ), .Q ( new_AGEMA_signal_5609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C ( clk ), .D ( new_AGEMA_signal_5636 ), .Q ( new_AGEMA_signal_5637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C ( clk ), .D ( new_AGEMA_signal_5652 ), .Q ( new_AGEMA_signal_5653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C ( clk ), .D ( new_AGEMA_signal_5662 ), .Q ( new_AGEMA_signal_5663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C ( clk ), .D ( new_AGEMA_signal_5672 ), .Q ( new_AGEMA_signal_5673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C ( clk ), .D ( n2829 ), .Q ( new_AGEMA_signal_5689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C ( clk ), .D ( new_AGEMA_signal_1768 ), .Q ( new_AGEMA_signal_5697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C ( clk ), .D ( new_AGEMA_signal_5734 ), .Q ( new_AGEMA_signal_5735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C ( clk ), .D ( new_AGEMA_signal_5750 ), .Q ( new_AGEMA_signal_5751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C ( clk ), .D ( n2312 ), .Q ( new_AGEMA_signal_5761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C ( clk ), .D ( new_AGEMA_signal_1742 ), .Q ( new_AGEMA_signal_5771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C ( clk ), .D ( new_AGEMA_signal_5788 ), .Q ( new_AGEMA_signal_5789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C ( clk ), .D ( new_AGEMA_signal_5806 ), .Q ( new_AGEMA_signal_5807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C ( clk ), .D ( new_AGEMA_signal_5888 ), .Q ( new_AGEMA_signal_5889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C ( clk ), .D ( new_AGEMA_signal_5908 ), .Q ( new_AGEMA_signal_5909 ) ) ;

    /* cells in depth 16 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2003 ( .a ({new_AGEMA_signal_4656, new_AGEMA_signal_4650}), .b ({new_AGEMA_signal_1726, n1935}), .clk ( clk ), .r ( Fresh[764] ), .c ({new_AGEMA_signal_1769, n1941}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2059 ( .a ({new_AGEMA_signal_1727, n1959}), .b ({new_AGEMA_signal_4660, new_AGEMA_signal_4658}), .clk ( clk ), .r ( Fresh[765] ), .c ({new_AGEMA_signal_1770, n1960}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2110 ( .a ({new_AGEMA_signal_4668, new_AGEMA_signal_4664}), .b ({new_AGEMA_signal_1728, n1983}), .clk ( clk ), .r ( Fresh[766] ), .c ({new_AGEMA_signal_1771, n1988}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2153 ( .a ({new_AGEMA_signal_1729, n2014}), .b ({new_AGEMA_signal_4684, new_AGEMA_signal_4676}), .clk ( clk ), .r ( Fresh[767] ), .c ({new_AGEMA_signal_1772, n2015}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2169 ( .a ({new_AGEMA_signal_1673, n2029}), .b ({new_AGEMA_signal_4700, new_AGEMA_signal_4692}), .clk ( clk ), .r ( Fresh[768] ), .c ({new_AGEMA_signal_1730, n2030}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2200 ( .a ({new_AGEMA_signal_1732, n2052}), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4708}), .clk ( clk ), .r ( Fresh[769] ), .c ({new_AGEMA_signal_1774, n2053}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2222 ( .a ({new_AGEMA_signal_1733, n2070}), .b ({new_AGEMA_signal_4732, new_AGEMA_signal_4724}), .clk ( clk ), .r ( Fresh[770] ), .c ({new_AGEMA_signal_1775, n2071}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2259 ( .a ({new_AGEMA_signal_4744, new_AGEMA_signal_4738}), .b ({new_AGEMA_signal_1734, n2098}), .clk ( clk ), .r ( Fresh[771] ), .c ({new_AGEMA_signal_1776, n2103}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2288 ( .a ({new_AGEMA_signal_4764, new_AGEMA_signal_4754}), .b ({new_AGEMA_signal_1736, n2125}), .clk ( clk ), .r ( Fresh[772] ), .c ({new_AGEMA_signal_1777, n2126}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2314 ( .a ({new_AGEMA_signal_1737, n2145}), .b ({new_AGEMA_signal_4780, new_AGEMA_signal_4772}), .clk ( clk ), .r ( Fresh[773] ), .c ({new_AGEMA_signal_1778, n2146}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2334 ( .a ({new_AGEMA_signal_4796, new_AGEMA_signal_4788}), .b ({new_AGEMA_signal_1738, n2169}), .clk ( clk ), .r ( Fresh[774] ), .c ({new_AGEMA_signal_1779, n2173}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2351 ( .a ({new_AGEMA_signal_4812, new_AGEMA_signal_4804}), .b ({new_AGEMA_signal_1739, n2185}), .clk ( clk ), .r ( Fresh[775] ), .c ({new_AGEMA_signal_1780, n2187}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2416 ( .a ({new_AGEMA_signal_4816, new_AGEMA_signal_4814}), .b ({new_AGEMA_signal_1744, n2251}), .clk ( clk ), .r ( Fresh[776] ), .c ({new_AGEMA_signal_1782, n2256}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2441 ( .a ({new_AGEMA_signal_1745, n2274}), .b ({new_AGEMA_signal_4824, new_AGEMA_signal_4820}), .clk ( clk ), .r ( Fresh[777] ), .c ({new_AGEMA_signal_1783, n2275}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2474 ( .a ({new_AGEMA_signal_1746, n2302}), .b ({new_AGEMA_signal_4836, new_AGEMA_signal_4830}), .clk ( clk ), .r ( Fresh[778] ), .c ({new_AGEMA_signal_1784, n2303}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2504 ( .a ({new_AGEMA_signal_1747, n2339}), .b ({new_AGEMA_signal_1748, n2338}), .clk ( clk ), .r ( Fresh[779] ), .c ({new_AGEMA_signal_1785, n2382}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2516 ( .a ({new_AGEMA_signal_1749, n2351}), .b ({new_AGEMA_signal_4844, new_AGEMA_signal_4840}), .clk ( clk ), .r ( Fresh[780] ), .c ({new_AGEMA_signal_1786, n2380}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2531 ( .a ({new_AGEMA_signal_1750, n2365}), .b ({new_AGEMA_signal_4864, new_AGEMA_signal_4854}), .clk ( clk ), .r ( Fresh[781] ), .c ({new_AGEMA_signal_1787, n2366}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2561 ( .a ({new_AGEMA_signal_1699, n2399}), .b ({new_AGEMA_signal_1751, n2398}), .clk ( clk ), .r ( Fresh[782] ), .c ({new_AGEMA_signal_1788, n2425}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2582 ( .a ({new_AGEMA_signal_1701, n2423}), .b ({new_AGEMA_signal_1702, n2422}), .clk ( clk ), .r ( Fresh[783] ), .c ({new_AGEMA_signal_1752, n2424}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2597 ( .a ({new_AGEMA_signal_4880, new_AGEMA_signal_4872}), .b ({new_AGEMA_signal_1753, n2441}), .clk ( clk ), .r ( Fresh[784] ), .c ({new_AGEMA_signal_1789, n2451}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2631 ( .a ({new_AGEMA_signal_1705, n2479}), .b ({new_AGEMA_signal_4888, new_AGEMA_signal_4884}), .clk ( clk ), .r ( Fresh[785] ), .c ({new_AGEMA_signal_1754, n2514}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2658 ( .a ({new_AGEMA_signal_1756, n2510}), .b ({new_AGEMA_signal_4892, new_AGEMA_signal_4890}), .clk ( clk ), .r ( Fresh[786] ), .c ({new_AGEMA_signal_1790, n2511}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2688 ( .a ({new_AGEMA_signal_1759, n2552}), .b ({new_AGEMA_signal_4908, new_AGEMA_signal_4900}), .clk ( clk ), .r ( Fresh[787] ), .c ({new_AGEMA_signal_1791, n2671}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2716 ( .a ({new_AGEMA_signal_1761, n2589}), .b ({new_AGEMA_signal_4924, new_AGEMA_signal_4916}), .clk ( clk ), .r ( Fresh[788] ), .c ({new_AGEMA_signal_1792, n2590}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2731 ( .a ({new_AGEMA_signal_1714, n2608}), .b ({new_AGEMA_signal_4936, new_AGEMA_signal_4930}), .clk ( clk ), .r ( Fresh[789] ), .c ({new_AGEMA_signal_1762, n2623}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2763 ( .a ({new_AGEMA_signal_4944, new_AGEMA_signal_4940}), .b ({new_AGEMA_signal_1764, n2659}), .clk ( clk ), .r ( Fresh[790] ), .c ({new_AGEMA_signal_1794, n2667}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2786 ( .a ({new_AGEMA_signal_1765, n2702}), .b ({new_AGEMA_signal_4960, new_AGEMA_signal_4952}), .clk ( clk ), .r ( Fresh[791] ), .c ({new_AGEMA_signal_1795, n2703}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) U2840 ( .s ({new_AGEMA_signal_4824, new_AGEMA_signal_4820}), .b ({new_AGEMA_signal_4964, new_AGEMA_signal_4962}), .a ({new_AGEMA_signal_1724, n2801}), .clk ( clk ), .r ( Fresh[792] ), .c ({new_AGEMA_signal_1767, n2803}) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C ( clk ), .D ( new_AGEMA_signal_4969 ), .Q ( new_AGEMA_signal_4970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C ( clk ), .D ( new_AGEMA_signal_4975 ), .Q ( new_AGEMA_signal_4976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C ( clk ), .D ( new_AGEMA_signal_4981 ), .Q ( new_AGEMA_signal_4982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C ( clk ), .D ( new_AGEMA_signal_4987 ), .Q ( new_AGEMA_signal_4988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C ( clk ), .D ( new_AGEMA_signal_4993 ), .Q ( new_AGEMA_signal_4994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C ( clk ), .D ( new_AGEMA_signal_4999 ), .Q ( new_AGEMA_signal_5000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C ( clk ), .D ( new_AGEMA_signal_5003 ), .Q ( new_AGEMA_signal_5004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C ( clk ), .D ( new_AGEMA_signal_5007 ), .Q ( new_AGEMA_signal_5008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C ( clk ), .D ( new_AGEMA_signal_5015 ), .Q ( new_AGEMA_signal_5016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C ( clk ), .D ( new_AGEMA_signal_5023 ), .Q ( new_AGEMA_signal_5024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C ( clk ), .D ( new_AGEMA_signal_5029 ), .Q ( new_AGEMA_signal_5030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C ( clk ), .D ( new_AGEMA_signal_5035 ), .Q ( new_AGEMA_signal_5036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C ( clk ), .D ( new_AGEMA_signal_5039 ), .Q ( new_AGEMA_signal_5040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C ( clk ), .D ( new_AGEMA_signal_5043 ), .Q ( new_AGEMA_signal_5044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C ( clk ), .D ( new_AGEMA_signal_5051 ), .Q ( new_AGEMA_signal_5052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C ( clk ), .D ( new_AGEMA_signal_5059 ), .Q ( new_AGEMA_signal_5060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C ( clk ), .D ( new_AGEMA_signal_5067 ), .Q ( new_AGEMA_signal_5068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C ( clk ), .D ( new_AGEMA_signal_5075 ), .Q ( new_AGEMA_signal_5076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C ( clk ), .D ( new_AGEMA_signal_5085 ), .Q ( new_AGEMA_signal_5086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C ( clk ), .D ( new_AGEMA_signal_5095 ), .Q ( new_AGEMA_signal_5096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C ( clk ), .D ( new_AGEMA_signal_5103 ), .Q ( new_AGEMA_signal_5104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C ( clk ), .D ( new_AGEMA_signal_5111 ), .Q ( new_AGEMA_signal_5112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C ( clk ), .D ( new_AGEMA_signal_5117 ), .Q ( new_AGEMA_signal_5118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C ( clk ), .D ( new_AGEMA_signal_5123 ), .Q ( new_AGEMA_signal_5124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C ( clk ), .D ( new_AGEMA_signal_5127 ), .Q ( new_AGEMA_signal_5128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C ( clk ), .D ( new_AGEMA_signal_5131 ), .Q ( new_AGEMA_signal_5132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C ( clk ), .D ( new_AGEMA_signal_5137 ), .Q ( new_AGEMA_signal_5138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C ( clk ), .D ( new_AGEMA_signal_5143 ), .Q ( new_AGEMA_signal_5144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C ( clk ), .D ( new_AGEMA_signal_5151 ), .Q ( new_AGEMA_signal_5152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C ( clk ), .D ( new_AGEMA_signal_5159 ), .Q ( new_AGEMA_signal_5160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C ( clk ), .D ( new_AGEMA_signal_5165 ), .Q ( new_AGEMA_signal_5166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C ( clk ), .D ( new_AGEMA_signal_5171 ), .Q ( new_AGEMA_signal_5172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C ( clk ), .D ( new_AGEMA_signal_5173 ), .Q ( new_AGEMA_signal_5174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C ( clk ), .D ( new_AGEMA_signal_5175 ), .Q ( new_AGEMA_signal_5176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C ( clk ), .D ( new_AGEMA_signal_5183 ), .Q ( new_AGEMA_signal_5184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C ( clk ), .D ( new_AGEMA_signal_5191 ), .Q ( new_AGEMA_signal_5192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C ( clk ), .D ( new_AGEMA_signal_5195 ), .Q ( new_AGEMA_signal_5196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C ( clk ), .D ( new_AGEMA_signal_5199 ), .Q ( new_AGEMA_signal_5200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C ( clk ), .D ( new_AGEMA_signal_5205 ), .Q ( new_AGEMA_signal_5206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C ( clk ), .D ( new_AGEMA_signal_5211 ), .Q ( new_AGEMA_signal_5212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C ( clk ), .D ( new_AGEMA_signal_5217 ), .Q ( new_AGEMA_signal_5218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C ( clk ), .D ( new_AGEMA_signal_5223 ), .Q ( new_AGEMA_signal_5224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C ( clk ), .D ( new_AGEMA_signal_5227 ), .Q ( new_AGEMA_signal_5228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C ( clk ), .D ( new_AGEMA_signal_5231 ), .Q ( new_AGEMA_signal_5232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C ( clk ), .D ( new_AGEMA_signal_5235 ), .Q ( new_AGEMA_signal_5236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C ( clk ), .D ( new_AGEMA_signal_5241 ), .Q ( new_AGEMA_signal_5242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C ( clk ), .D ( new_AGEMA_signal_5245 ), .Q ( new_AGEMA_signal_5246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C ( clk ), .D ( new_AGEMA_signal_5249 ), .Q ( new_AGEMA_signal_5250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C ( clk ), .D ( new_AGEMA_signal_5255 ), .Q ( new_AGEMA_signal_5256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C ( clk ), .D ( new_AGEMA_signal_5261 ), .Q ( new_AGEMA_signal_5262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C ( clk ), .D ( new_AGEMA_signal_5271 ), .Q ( new_AGEMA_signal_5272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C ( clk ), .D ( new_AGEMA_signal_5281 ), .Q ( new_AGEMA_signal_5282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C ( clk ), .D ( new_AGEMA_signal_5287 ), .Q ( new_AGEMA_signal_5288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C ( clk ), .D ( new_AGEMA_signal_5293 ), .Q ( new_AGEMA_signal_5294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C ( clk ), .D ( new_AGEMA_signal_5299 ), .Q ( new_AGEMA_signal_5300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C ( clk ), .D ( new_AGEMA_signal_5305 ), .Q ( new_AGEMA_signal_5306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C ( clk ), .D ( new_AGEMA_signal_5309 ), .Q ( new_AGEMA_signal_5310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C ( clk ), .D ( new_AGEMA_signal_5313 ), .Q ( new_AGEMA_signal_5314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C ( clk ), .D ( new_AGEMA_signal_5317 ), .Q ( new_AGEMA_signal_5318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C ( clk ), .D ( new_AGEMA_signal_5321 ), .Q ( new_AGEMA_signal_5322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C ( clk ), .D ( new_AGEMA_signal_5329 ), .Q ( new_AGEMA_signal_5330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C ( clk ), .D ( new_AGEMA_signal_5337 ), .Q ( new_AGEMA_signal_5338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C ( clk ), .D ( new_AGEMA_signal_5343 ), .Q ( new_AGEMA_signal_5344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C ( clk ), .D ( new_AGEMA_signal_5349 ), .Q ( new_AGEMA_signal_5350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C ( clk ), .D ( new_AGEMA_signal_5357 ), .Q ( new_AGEMA_signal_5358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C ( clk ), .D ( new_AGEMA_signal_5365 ), .Q ( new_AGEMA_signal_5366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C ( clk ), .D ( new_AGEMA_signal_5373 ), .Q ( new_AGEMA_signal_5374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C ( clk ), .D ( new_AGEMA_signal_5381 ), .Q ( new_AGEMA_signal_5382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C ( clk ), .D ( new_AGEMA_signal_5389 ), .Q ( new_AGEMA_signal_5390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C ( clk ), .D ( new_AGEMA_signal_5393 ), .Q ( new_AGEMA_signal_5394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C ( clk ), .D ( new_AGEMA_signal_5397 ), .Q ( new_AGEMA_signal_5398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C ( clk ), .D ( new_AGEMA_signal_5401 ), .Q ( new_AGEMA_signal_5402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C ( clk ), .D ( new_AGEMA_signal_5409 ), .Q ( new_AGEMA_signal_5410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C ( clk ), .D ( new_AGEMA_signal_5417 ), .Q ( new_AGEMA_signal_5418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C ( clk ), .D ( new_AGEMA_signal_5421 ), .Q ( new_AGEMA_signal_5422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C ( clk ), .D ( new_AGEMA_signal_5425 ), .Q ( new_AGEMA_signal_5426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C ( clk ), .D ( new_AGEMA_signal_5431 ), .Q ( new_AGEMA_signal_5432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C ( clk ), .D ( new_AGEMA_signal_5439 ), .Q ( new_AGEMA_signal_5440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C ( clk ), .D ( new_AGEMA_signal_5451 ), .Q ( new_AGEMA_signal_5452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C ( clk ), .D ( new_AGEMA_signal_5463 ), .Q ( new_AGEMA_signal_5464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C ( clk ), .D ( new_AGEMA_signal_5477 ), .Q ( new_AGEMA_signal_5478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C ( clk ), .D ( new_AGEMA_signal_5491 ), .Q ( new_AGEMA_signal_5492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C ( clk ), .D ( new_AGEMA_signal_5499 ), .Q ( new_AGEMA_signal_5500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C ( clk ), .D ( new_AGEMA_signal_5507 ), .Q ( new_AGEMA_signal_5508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C ( clk ), .D ( new_AGEMA_signal_5521 ), .Q ( new_AGEMA_signal_5522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C ( clk ), .D ( new_AGEMA_signal_5535 ), .Q ( new_AGEMA_signal_5536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C ( clk ), .D ( new_AGEMA_signal_5543 ), .Q ( new_AGEMA_signal_5544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C ( clk ), .D ( new_AGEMA_signal_5551 ), .Q ( new_AGEMA_signal_5552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C ( clk ), .D ( new_AGEMA_signal_5559 ), .Q ( new_AGEMA_signal_5560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C ( clk ), .D ( new_AGEMA_signal_5567 ), .Q ( new_AGEMA_signal_5568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C ( clk ), .D ( new_AGEMA_signal_5593 ), .Q ( new_AGEMA_signal_5594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C ( clk ), .D ( new_AGEMA_signal_5609 ), .Q ( new_AGEMA_signal_5610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C ( clk ), .D ( new_AGEMA_signal_5637 ), .Q ( new_AGEMA_signal_5638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C ( clk ), .D ( new_AGEMA_signal_5653 ), .Q ( new_AGEMA_signal_5654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C ( clk ), .D ( new_AGEMA_signal_5663 ), .Q ( new_AGEMA_signal_5664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C ( clk ), .D ( new_AGEMA_signal_5673 ), .Q ( new_AGEMA_signal_5674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C ( clk ), .D ( new_AGEMA_signal_5689 ), .Q ( new_AGEMA_signal_5690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C ( clk ), .D ( new_AGEMA_signal_5697 ), .Q ( new_AGEMA_signal_5698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C ( clk ), .D ( new_AGEMA_signal_5735 ), .Q ( new_AGEMA_signal_5736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C ( clk ), .D ( new_AGEMA_signal_5751 ), .Q ( new_AGEMA_signal_5752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C ( clk ), .D ( new_AGEMA_signal_5761 ), .Q ( new_AGEMA_signal_5762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C ( clk ), .D ( new_AGEMA_signal_5771 ), .Q ( new_AGEMA_signal_5772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C ( clk ), .D ( new_AGEMA_signal_5789 ), .Q ( new_AGEMA_signal_5790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C ( clk ), .D ( new_AGEMA_signal_5807 ), .Q ( new_AGEMA_signal_5808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C ( clk ), .D ( new_AGEMA_signal_5889 ), .Q ( new_AGEMA_signal_5890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C ( clk ), .D ( new_AGEMA_signal_5909 ), .Q ( new_AGEMA_signal_5910 ) ) ;

    /* cells in depth 17 */
    buf_clk new_AGEMA_reg_buffer_3419 ( .C ( clk ), .D ( new_AGEMA_signal_5236 ), .Q ( new_AGEMA_signal_5237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C ( clk ), .D ( new_AGEMA_signal_5242 ), .Q ( new_AGEMA_signal_5243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C ( clk ), .D ( new_AGEMA_signal_5246 ), .Q ( new_AGEMA_signal_5247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C ( clk ), .D ( new_AGEMA_signal_5250 ), .Q ( new_AGEMA_signal_5251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C ( clk ), .D ( new_AGEMA_signal_5256 ), .Q ( new_AGEMA_signal_5257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C ( clk ), .D ( new_AGEMA_signal_5262 ), .Q ( new_AGEMA_signal_5263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C ( clk ), .D ( new_AGEMA_signal_5272 ), .Q ( new_AGEMA_signal_5273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C ( clk ), .D ( new_AGEMA_signal_5282 ), .Q ( new_AGEMA_signal_5283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C ( clk ), .D ( new_AGEMA_signal_5288 ), .Q ( new_AGEMA_signal_5289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C ( clk ), .D ( new_AGEMA_signal_5294 ), .Q ( new_AGEMA_signal_5295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C ( clk ), .D ( new_AGEMA_signal_5300 ), .Q ( new_AGEMA_signal_5301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C ( clk ), .D ( new_AGEMA_signal_5306 ), .Q ( new_AGEMA_signal_5307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C ( clk ), .D ( new_AGEMA_signal_5310 ), .Q ( new_AGEMA_signal_5311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C ( clk ), .D ( new_AGEMA_signal_5314 ), .Q ( new_AGEMA_signal_5315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C ( clk ), .D ( new_AGEMA_signal_5318 ), .Q ( new_AGEMA_signal_5319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C ( clk ), .D ( new_AGEMA_signal_5322 ), .Q ( new_AGEMA_signal_5323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C ( clk ), .D ( new_AGEMA_signal_5330 ), .Q ( new_AGEMA_signal_5331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C ( clk ), .D ( new_AGEMA_signal_5338 ), .Q ( new_AGEMA_signal_5339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C ( clk ), .D ( new_AGEMA_signal_5344 ), .Q ( new_AGEMA_signal_5345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C ( clk ), .D ( new_AGEMA_signal_5350 ), .Q ( new_AGEMA_signal_5351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C ( clk ), .D ( new_AGEMA_signal_5358 ), .Q ( new_AGEMA_signal_5359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C ( clk ), .D ( new_AGEMA_signal_5366 ), .Q ( new_AGEMA_signal_5367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C ( clk ), .D ( new_AGEMA_signal_5374 ), .Q ( new_AGEMA_signal_5375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C ( clk ), .D ( new_AGEMA_signal_5382 ), .Q ( new_AGEMA_signal_5383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C ( clk ), .D ( n2514 ), .Q ( new_AGEMA_signal_5385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C ( clk ), .D ( new_AGEMA_signal_1754 ), .Q ( new_AGEMA_signal_5387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C ( clk ), .D ( new_AGEMA_signal_5390 ), .Q ( new_AGEMA_signal_5391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C ( clk ), .D ( new_AGEMA_signal_5394 ), .Q ( new_AGEMA_signal_5395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C ( clk ), .D ( new_AGEMA_signal_5398 ), .Q ( new_AGEMA_signal_5399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C ( clk ), .D ( new_AGEMA_signal_5402 ), .Q ( new_AGEMA_signal_5403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C ( clk ), .D ( new_AGEMA_signal_5410 ), .Q ( new_AGEMA_signal_5411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C ( clk ), .D ( new_AGEMA_signal_5418 ), .Q ( new_AGEMA_signal_5419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C ( clk ), .D ( new_AGEMA_signal_5422 ), .Q ( new_AGEMA_signal_5423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C ( clk ), .D ( new_AGEMA_signal_5426 ), .Q ( new_AGEMA_signal_5427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C ( clk ), .D ( new_AGEMA_signal_5432 ), .Q ( new_AGEMA_signal_5433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C ( clk ), .D ( new_AGEMA_signal_5440 ), .Q ( new_AGEMA_signal_5441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C ( clk ), .D ( new_AGEMA_signal_5452 ), .Q ( new_AGEMA_signal_5453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C ( clk ), .D ( new_AGEMA_signal_5464 ), .Q ( new_AGEMA_signal_5465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C ( clk ), .D ( new_AGEMA_signal_5478 ), .Q ( new_AGEMA_signal_5479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C ( clk ), .D ( new_AGEMA_signal_5492 ), .Q ( new_AGEMA_signal_5493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C ( clk ), .D ( new_AGEMA_signal_5500 ), .Q ( new_AGEMA_signal_5501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C ( clk ), .D ( new_AGEMA_signal_5508 ), .Q ( new_AGEMA_signal_5509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C ( clk ), .D ( new_AGEMA_signal_5522 ), .Q ( new_AGEMA_signal_5523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C ( clk ), .D ( new_AGEMA_signal_5536 ), .Q ( new_AGEMA_signal_5537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C ( clk ), .D ( new_AGEMA_signal_5544 ), .Q ( new_AGEMA_signal_5545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C ( clk ), .D ( new_AGEMA_signal_5552 ), .Q ( new_AGEMA_signal_5553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C ( clk ), .D ( new_AGEMA_signal_5560 ), .Q ( new_AGEMA_signal_5561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C ( clk ), .D ( new_AGEMA_signal_5568 ), .Q ( new_AGEMA_signal_5569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C ( clk ), .D ( new_AGEMA_signal_5594 ), .Q ( new_AGEMA_signal_5595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C ( clk ), .D ( new_AGEMA_signal_5610 ), .Q ( new_AGEMA_signal_5611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C ( clk ), .D ( new_AGEMA_signal_5638 ), .Q ( new_AGEMA_signal_5639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C ( clk ), .D ( new_AGEMA_signal_5654 ), .Q ( new_AGEMA_signal_5655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C ( clk ), .D ( new_AGEMA_signal_5664 ), .Q ( new_AGEMA_signal_5665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C ( clk ), .D ( new_AGEMA_signal_5674 ), .Q ( new_AGEMA_signal_5675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C ( clk ), .D ( new_AGEMA_signal_5690 ), .Q ( new_AGEMA_signal_5691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C ( clk ), .D ( new_AGEMA_signal_5698 ), .Q ( new_AGEMA_signal_5699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C ( clk ), .D ( new_AGEMA_signal_5736 ), .Q ( new_AGEMA_signal_5737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C ( clk ), .D ( new_AGEMA_signal_5752 ), .Q ( new_AGEMA_signal_5753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C ( clk ), .D ( new_AGEMA_signal_5762 ), .Q ( new_AGEMA_signal_5763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C ( clk ), .D ( new_AGEMA_signal_5772 ), .Q ( new_AGEMA_signal_5773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C ( clk ), .D ( new_AGEMA_signal_5790 ), .Q ( new_AGEMA_signal_5791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C ( clk ), .D ( new_AGEMA_signal_5808 ), .Q ( new_AGEMA_signal_5809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C ( clk ), .D ( n2671 ), .Q ( new_AGEMA_signal_5825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C ( clk ), .D ( new_AGEMA_signal_1791 ), .Q ( new_AGEMA_signal_5833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C ( clk ), .D ( new_AGEMA_signal_5890 ), .Q ( new_AGEMA_signal_5891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C ( clk ), .D ( new_AGEMA_signal_5910 ), .Q ( new_AGEMA_signal_5911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C ( clk ), .D ( n2380 ), .Q ( new_AGEMA_signal_5937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C ( clk ), .D ( new_AGEMA_signal_1786 ), .Q ( new_AGEMA_signal_5949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C ( clk ), .D ( n2382 ), .Q ( new_AGEMA_signal_5961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C ( clk ), .D ( new_AGEMA_signal_1785 ), .Q ( new_AGEMA_signal_5975 ) ) ;

    /* cells in depth 18 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2016 ( .a ({new_AGEMA_signal_1769, n1941}), .b ({new_AGEMA_signal_4976, new_AGEMA_signal_4970}), .clk ( clk ), .r ( Fresh[793] ), .c ({new_AGEMA_signal_1797, n2019}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2060 ( .a ({new_AGEMA_signal_4988, new_AGEMA_signal_4982}), .b ({new_AGEMA_signal_1770, n1960}), .clk ( clk ), .r ( Fresh[794] ), .c ({new_AGEMA_signal_1798, n2002}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2116 ( .a ({new_AGEMA_signal_1771, n1988}), .b ({new_AGEMA_signal_5000, new_AGEMA_signal_4994}), .clk ( clk ), .r ( Fresh[795] ), .c ({new_AGEMA_signal_1799, n1989}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2154 ( .a ({new_AGEMA_signal_5008, new_AGEMA_signal_5004}), .b ({new_AGEMA_signal_1772, n2015}), .clk ( clk ), .r ( Fresh[796] ), .c ({new_AGEMA_signal_1800, n2016}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2170 ( .a ({new_AGEMA_signal_5024, new_AGEMA_signal_5016}), .b ({new_AGEMA_signal_1730, n2030}), .clk ( clk ), .r ( Fresh[797] ), .c ({new_AGEMA_signal_1773, n2038}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2201 ( .a ({new_AGEMA_signal_5036, new_AGEMA_signal_5030}), .b ({new_AGEMA_signal_1774, n2053}), .clk ( clk ), .r ( Fresh[798] ), .c ({new_AGEMA_signal_1802, n2111}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2223 ( .a ({new_AGEMA_signal_5044, new_AGEMA_signal_5040}), .b ({new_AGEMA_signal_1775, n2071}), .clk ( clk ), .r ( Fresh[799] ), .c ({new_AGEMA_signal_1803, n2079}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2263 ( .a ({new_AGEMA_signal_1776, n2103}), .b ({new_AGEMA_signal_5060, new_AGEMA_signal_5052}), .clk ( clk ), .r ( Fresh[800] ), .c ({new_AGEMA_signal_1804, n2104}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2289 ( .a ({new_AGEMA_signal_5076, new_AGEMA_signal_5068}), .b ({new_AGEMA_signal_1777, n2126}), .clk ( clk ), .r ( Fresh[801] ), .c ({new_AGEMA_signal_1805, n2127}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2315 ( .a ({new_AGEMA_signal_5008, new_AGEMA_signal_5004}), .b ({new_AGEMA_signal_1778, n2146}), .clk ( clk ), .r ( Fresh[802] ), .c ({new_AGEMA_signal_1806, n2147}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2336 ( .a ({new_AGEMA_signal_1779, n2173}), .b ({new_AGEMA_signal_5096, new_AGEMA_signal_5086}), .clk ( clk ), .r ( Fresh[803] ), .c ({new_AGEMA_signal_1807, n2208}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2352 ( .a ({new_AGEMA_signal_1780, n2187}), .b ({new_AGEMA_signal_5112, new_AGEMA_signal_5104}), .clk ( clk ), .r ( Fresh[804] ), .c ({new_AGEMA_signal_1808, n2199}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2420 ( .a ({new_AGEMA_signal_1782, n2256}), .b ({new_AGEMA_signal_5124, new_AGEMA_signal_5118}), .clk ( clk ), .r ( Fresh[805] ), .c ({new_AGEMA_signal_1809, n2257}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2442 ( .a ({new_AGEMA_signal_5132, new_AGEMA_signal_5128}), .b ({new_AGEMA_signal_1783, n2275}), .clk ( clk ), .r ( Fresh[806] ), .c ({new_AGEMA_signal_1810, n2281}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2475 ( .a ({new_AGEMA_signal_5144, new_AGEMA_signal_5138}), .b ({new_AGEMA_signal_1784, n2303}), .clk ( clk ), .r ( Fresh[807] ), .c ({new_AGEMA_signal_1811, n2305}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2532 ( .a ({new_AGEMA_signal_5160, new_AGEMA_signal_5152}), .b ({new_AGEMA_signal_1787, n2366}), .clk ( clk ), .r ( Fresh[808] ), .c ({new_AGEMA_signal_1812, n2368}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2583 ( .a ({new_AGEMA_signal_1788, n2425}), .b ({new_AGEMA_signal_1752, n2424}), .clk ( clk ), .r ( Fresh[809] ), .c ({new_AGEMA_signal_1813, n2426}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2605 ( .a ({new_AGEMA_signal_1789, n2451}), .b ({new_AGEMA_signal_5172, new_AGEMA_signal_5166}), .clk ( clk ), .r ( Fresh[810] ), .c ({new_AGEMA_signal_1814, n2457}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2659 ( .a ({new_AGEMA_signal_5176, new_AGEMA_signal_5174}), .b ({new_AGEMA_signal_1790, n2511}), .clk ( clk ), .r ( Fresh[811] ), .c ({new_AGEMA_signal_1815, n2513}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2717 ( .a ({new_AGEMA_signal_5192, new_AGEMA_signal_5184}), .b ({new_AGEMA_signal_1792, n2590}), .clk ( clk ), .r ( Fresh[812] ), .c ({new_AGEMA_signal_1816, n2592}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2741 ( .a ({new_AGEMA_signal_1762, n2623}), .b ({new_AGEMA_signal_5200, new_AGEMA_signal_5196}), .clk ( clk ), .r ( Fresh[813] ), .c ({new_AGEMA_signal_1793, n2637}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2767 ( .a ({new_AGEMA_signal_1794, n2667}), .b ({new_AGEMA_signal_5212, new_AGEMA_signal_5206}), .clk ( clk ), .r ( Fresh[814] ), .c ({new_AGEMA_signal_1818, n2668}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2787 ( .a ({new_AGEMA_signal_5224, new_AGEMA_signal_5218}), .b ({new_AGEMA_signal_1795, n2703}), .clk ( clk ), .r ( Fresh[815] ), .c ({new_AGEMA_signal_1819, n2705}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2841 ( .a ({new_AGEMA_signal_5232, new_AGEMA_signal_5228}), .b ({new_AGEMA_signal_1767, n2803}), .clk ( clk ), .r ( Fresh[816] ), .c ({new_AGEMA_signal_1796, n2805}) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C ( clk ), .D ( new_AGEMA_signal_5237 ), .Q ( new_AGEMA_signal_5238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C ( clk ), .D ( new_AGEMA_signal_5243 ), .Q ( new_AGEMA_signal_5244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C ( clk ), .D ( new_AGEMA_signal_5247 ), .Q ( new_AGEMA_signal_5248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C ( clk ), .D ( new_AGEMA_signal_5251 ), .Q ( new_AGEMA_signal_5252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C ( clk ), .D ( new_AGEMA_signal_5257 ), .Q ( new_AGEMA_signal_5258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C ( clk ), .D ( new_AGEMA_signal_5263 ), .Q ( new_AGEMA_signal_5264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C ( clk ), .D ( new_AGEMA_signal_5273 ), .Q ( new_AGEMA_signal_5274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C ( clk ), .D ( new_AGEMA_signal_5283 ), .Q ( new_AGEMA_signal_5284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C ( clk ), .D ( new_AGEMA_signal_5289 ), .Q ( new_AGEMA_signal_5290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C ( clk ), .D ( new_AGEMA_signal_5295 ), .Q ( new_AGEMA_signal_5296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C ( clk ), .D ( new_AGEMA_signal_5301 ), .Q ( new_AGEMA_signal_5302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C ( clk ), .D ( new_AGEMA_signal_5307 ), .Q ( new_AGEMA_signal_5308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C ( clk ), .D ( new_AGEMA_signal_5311 ), .Q ( new_AGEMA_signal_5312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C ( clk ), .D ( new_AGEMA_signal_5315 ), .Q ( new_AGEMA_signal_5316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C ( clk ), .D ( new_AGEMA_signal_5319 ), .Q ( new_AGEMA_signal_5320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C ( clk ), .D ( new_AGEMA_signal_5323 ), .Q ( new_AGEMA_signal_5324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C ( clk ), .D ( new_AGEMA_signal_5331 ), .Q ( new_AGEMA_signal_5332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C ( clk ), .D ( new_AGEMA_signal_5339 ), .Q ( new_AGEMA_signal_5340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C ( clk ), .D ( new_AGEMA_signal_5345 ), .Q ( new_AGEMA_signal_5346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C ( clk ), .D ( new_AGEMA_signal_5351 ), .Q ( new_AGEMA_signal_5352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C ( clk ), .D ( new_AGEMA_signal_5359 ), .Q ( new_AGEMA_signal_5360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C ( clk ), .D ( new_AGEMA_signal_5367 ), .Q ( new_AGEMA_signal_5368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C ( clk ), .D ( new_AGEMA_signal_5375 ), .Q ( new_AGEMA_signal_5376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C ( clk ), .D ( new_AGEMA_signal_5383 ), .Q ( new_AGEMA_signal_5384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C ( clk ), .D ( new_AGEMA_signal_5385 ), .Q ( new_AGEMA_signal_5386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C ( clk ), .D ( new_AGEMA_signal_5387 ), .Q ( new_AGEMA_signal_5388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C ( clk ), .D ( new_AGEMA_signal_5391 ), .Q ( new_AGEMA_signal_5392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C ( clk ), .D ( new_AGEMA_signal_5395 ), .Q ( new_AGEMA_signal_5396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C ( clk ), .D ( new_AGEMA_signal_5399 ), .Q ( new_AGEMA_signal_5400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C ( clk ), .D ( new_AGEMA_signal_5403 ), .Q ( new_AGEMA_signal_5404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C ( clk ), .D ( new_AGEMA_signal_5411 ), .Q ( new_AGEMA_signal_5412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C ( clk ), .D ( new_AGEMA_signal_5419 ), .Q ( new_AGEMA_signal_5420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C ( clk ), .D ( new_AGEMA_signal_5423 ), .Q ( new_AGEMA_signal_5424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C ( clk ), .D ( new_AGEMA_signal_5427 ), .Q ( new_AGEMA_signal_5428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C ( clk ), .D ( new_AGEMA_signal_5433 ), .Q ( new_AGEMA_signal_5434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C ( clk ), .D ( new_AGEMA_signal_5441 ), .Q ( new_AGEMA_signal_5442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C ( clk ), .D ( new_AGEMA_signal_5453 ), .Q ( new_AGEMA_signal_5454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C ( clk ), .D ( new_AGEMA_signal_5465 ), .Q ( new_AGEMA_signal_5466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C ( clk ), .D ( new_AGEMA_signal_5479 ), .Q ( new_AGEMA_signal_5480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C ( clk ), .D ( new_AGEMA_signal_5493 ), .Q ( new_AGEMA_signal_5494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C ( clk ), .D ( new_AGEMA_signal_5501 ), .Q ( new_AGEMA_signal_5502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C ( clk ), .D ( new_AGEMA_signal_5509 ), .Q ( new_AGEMA_signal_5510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C ( clk ), .D ( new_AGEMA_signal_5523 ), .Q ( new_AGEMA_signal_5524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C ( clk ), .D ( new_AGEMA_signal_5537 ), .Q ( new_AGEMA_signal_5538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C ( clk ), .D ( new_AGEMA_signal_5545 ), .Q ( new_AGEMA_signal_5546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C ( clk ), .D ( new_AGEMA_signal_5553 ), .Q ( new_AGEMA_signal_5554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C ( clk ), .D ( new_AGEMA_signal_5561 ), .Q ( new_AGEMA_signal_5562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C ( clk ), .D ( new_AGEMA_signal_5569 ), .Q ( new_AGEMA_signal_5570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C ( clk ), .D ( new_AGEMA_signal_5595 ), .Q ( new_AGEMA_signal_5596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C ( clk ), .D ( new_AGEMA_signal_5611 ), .Q ( new_AGEMA_signal_5612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C ( clk ), .D ( new_AGEMA_signal_5639 ), .Q ( new_AGEMA_signal_5640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C ( clk ), .D ( new_AGEMA_signal_5655 ), .Q ( new_AGEMA_signal_5656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C ( clk ), .D ( new_AGEMA_signal_5665 ), .Q ( new_AGEMA_signal_5666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C ( clk ), .D ( new_AGEMA_signal_5675 ), .Q ( new_AGEMA_signal_5676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C ( clk ), .D ( new_AGEMA_signal_5691 ), .Q ( new_AGEMA_signal_5692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C ( clk ), .D ( new_AGEMA_signal_5699 ), .Q ( new_AGEMA_signal_5700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C ( clk ), .D ( new_AGEMA_signal_5737 ), .Q ( new_AGEMA_signal_5738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C ( clk ), .D ( new_AGEMA_signal_5753 ), .Q ( new_AGEMA_signal_5754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C ( clk ), .D ( new_AGEMA_signal_5763 ), .Q ( new_AGEMA_signal_5764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C ( clk ), .D ( new_AGEMA_signal_5773 ), .Q ( new_AGEMA_signal_5774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C ( clk ), .D ( new_AGEMA_signal_5791 ), .Q ( new_AGEMA_signal_5792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C ( clk ), .D ( new_AGEMA_signal_5809 ), .Q ( new_AGEMA_signal_5810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C ( clk ), .D ( new_AGEMA_signal_5825 ), .Q ( new_AGEMA_signal_5826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C ( clk ), .D ( new_AGEMA_signal_5833 ), .Q ( new_AGEMA_signal_5834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C ( clk ), .D ( new_AGEMA_signal_5891 ), .Q ( new_AGEMA_signal_5892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C ( clk ), .D ( new_AGEMA_signal_5911 ), .Q ( new_AGEMA_signal_5912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C ( clk ), .D ( new_AGEMA_signal_5937 ), .Q ( new_AGEMA_signal_5938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C ( clk ), .D ( new_AGEMA_signal_5949 ), .Q ( new_AGEMA_signal_5950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C ( clk ), .D ( new_AGEMA_signal_5961 ), .Q ( new_AGEMA_signal_5962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C ( clk ), .D ( new_AGEMA_signal_5975 ), .Q ( new_AGEMA_signal_5976 ) ) ;

    /* cells in depth 19 */
    buf_clk new_AGEMA_reg_buffer_3617 ( .C ( clk ), .D ( new_AGEMA_signal_5434 ), .Q ( new_AGEMA_signal_5435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C ( clk ), .D ( new_AGEMA_signal_5442 ), .Q ( new_AGEMA_signal_5443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C ( clk ), .D ( new_AGEMA_signal_5454 ), .Q ( new_AGEMA_signal_5455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C ( clk ), .D ( new_AGEMA_signal_5466 ), .Q ( new_AGEMA_signal_5467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C ( clk ), .D ( new_AGEMA_signal_5480 ), .Q ( new_AGEMA_signal_5481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C ( clk ), .D ( new_AGEMA_signal_5494 ), .Q ( new_AGEMA_signal_5495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C ( clk ), .D ( new_AGEMA_signal_5502 ), .Q ( new_AGEMA_signal_5503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C ( clk ), .D ( new_AGEMA_signal_5510 ), .Q ( new_AGEMA_signal_5511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C ( clk ), .D ( new_AGEMA_signal_5524 ), .Q ( new_AGEMA_signal_5525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C ( clk ), .D ( new_AGEMA_signal_5538 ), .Q ( new_AGEMA_signal_5539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C ( clk ), .D ( new_AGEMA_signal_5546 ), .Q ( new_AGEMA_signal_5547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C ( clk ), .D ( new_AGEMA_signal_5554 ), .Q ( new_AGEMA_signal_5555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C ( clk ), .D ( new_AGEMA_signal_5562 ), .Q ( new_AGEMA_signal_5563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C ( clk ), .D ( new_AGEMA_signal_5570 ), .Q ( new_AGEMA_signal_5571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C ( clk ), .D ( n2002 ), .Q ( new_AGEMA_signal_5573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C ( clk ), .D ( new_AGEMA_signal_1798 ), .Q ( new_AGEMA_signal_5577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C ( clk ), .D ( new_AGEMA_signal_5596 ), .Q ( new_AGEMA_signal_5597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C ( clk ), .D ( new_AGEMA_signal_5612 ), .Q ( new_AGEMA_signal_5613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C ( clk ), .D ( n2208 ), .Q ( new_AGEMA_signal_5617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C ( clk ), .D ( new_AGEMA_signal_1807 ), .Q ( new_AGEMA_signal_5621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C ( clk ), .D ( new_AGEMA_signal_5640 ), .Q ( new_AGEMA_signal_5641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C ( clk ), .D ( new_AGEMA_signal_5656 ), .Q ( new_AGEMA_signal_5657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C ( clk ), .D ( new_AGEMA_signal_5666 ), .Q ( new_AGEMA_signal_5667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C ( clk ), .D ( new_AGEMA_signal_5676 ), .Q ( new_AGEMA_signal_5677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C ( clk ), .D ( n2668 ), .Q ( new_AGEMA_signal_5681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C ( clk ), .D ( new_AGEMA_signal_1818 ), .Q ( new_AGEMA_signal_5685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C ( clk ), .D ( new_AGEMA_signal_5692 ), .Q ( new_AGEMA_signal_5693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C ( clk ), .D ( new_AGEMA_signal_5700 ), .Q ( new_AGEMA_signal_5701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C ( clk ), .D ( n2016 ), .Q ( new_AGEMA_signal_5705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C ( clk ), .D ( new_AGEMA_signal_1800 ), .Q ( new_AGEMA_signal_5711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C ( clk ), .D ( n2111 ), .Q ( new_AGEMA_signal_5717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C ( clk ), .D ( new_AGEMA_signal_1802 ), .Q ( new_AGEMA_signal_5723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C ( clk ), .D ( new_AGEMA_signal_5738 ), .Q ( new_AGEMA_signal_5739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C ( clk ), .D ( new_AGEMA_signal_5754 ), .Q ( new_AGEMA_signal_5755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C ( clk ), .D ( new_AGEMA_signal_5764 ), .Q ( new_AGEMA_signal_5765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C ( clk ), .D ( new_AGEMA_signal_5774 ), .Q ( new_AGEMA_signal_5775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C ( clk ), .D ( new_AGEMA_signal_5792 ), .Q ( new_AGEMA_signal_5793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C ( clk ), .D ( new_AGEMA_signal_5810 ), .Q ( new_AGEMA_signal_5811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C ( clk ), .D ( new_AGEMA_signal_5826 ), .Q ( new_AGEMA_signal_5827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C ( clk ), .D ( new_AGEMA_signal_5834 ), .Q ( new_AGEMA_signal_5835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C ( clk ), .D ( n2019 ), .Q ( new_AGEMA_signal_5849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C ( clk ), .D ( new_AGEMA_signal_1797 ), .Q ( new_AGEMA_signal_5857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C ( clk ), .D ( new_AGEMA_signal_5892 ), .Q ( new_AGEMA_signal_5893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C ( clk ), .D ( new_AGEMA_signal_5912 ), .Q ( new_AGEMA_signal_5913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C ( clk ), .D ( new_AGEMA_signal_5938 ), .Q ( new_AGEMA_signal_5939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C ( clk ), .D ( new_AGEMA_signal_5950 ), .Q ( new_AGEMA_signal_5951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C ( clk ), .D ( new_AGEMA_signal_5962 ), .Q ( new_AGEMA_signal_5963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C ( clk ), .D ( new_AGEMA_signal_5976 ), .Q ( new_AGEMA_signal_5977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C ( clk ), .D ( n2426 ), .Q ( new_AGEMA_signal_5989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C ( clk ), .D ( new_AGEMA_signal_1813 ), .Q ( new_AGEMA_signal_6003 ) ) ;

    /* cells in depth 20 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2117 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5238}), .b ({new_AGEMA_signal_1799, n1989}), .clk ( clk ), .r ( Fresh[817] ), .c ({new_AGEMA_signal_1821, n2000}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2181 ( .a ({new_AGEMA_signal_1773, n2038}), .b ({new_AGEMA_signal_5252, new_AGEMA_signal_5248}), .clk ( clk ), .r ( Fresh[818] ), .c ({new_AGEMA_signal_1801, n2113}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2231 ( .a ({new_AGEMA_signal_1803, n2079}), .b ({new_AGEMA_signal_5264, new_AGEMA_signal_5258}), .clk ( clk ), .r ( Fresh[819] ), .c ({new_AGEMA_signal_1822, n2109}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2264 ( .a ({new_AGEMA_signal_5284, new_AGEMA_signal_5274}), .b ({new_AGEMA_signal_1804, n2104}), .clk ( clk ), .r ( Fresh[820] ), .c ({new_AGEMA_signal_1823, n2107}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2290 ( .a ({new_AGEMA_signal_5296, new_AGEMA_signal_5290}), .b ({new_AGEMA_signal_1805, n2127}), .clk ( clk ), .r ( Fresh[821] ), .c ({new_AGEMA_signal_1824, n2212}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2316 ( .a ({new_AGEMA_signal_5308, new_AGEMA_signal_5302}), .b ({new_AGEMA_signal_1806, n2147}), .clk ( clk ), .r ( Fresh[822] ), .c ({new_AGEMA_signal_1825, n2149}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2366 ( .a ({new_AGEMA_signal_1808, n2199}), .b ({new_AGEMA_signal_5316, new_AGEMA_signal_5312}), .clk ( clk ), .r ( Fresh[823] ), .c ({new_AGEMA_signal_1826, n2206}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2421 ( .a ({new_AGEMA_signal_5324, new_AGEMA_signal_5320}), .b ({new_AGEMA_signal_1809, n2257}), .clk ( clk ), .r ( Fresh[824] ), .c ({new_AGEMA_signal_1827, n2310}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2447 ( .a ({new_AGEMA_signal_1810, n2281}), .b ({new_AGEMA_signal_5340, new_AGEMA_signal_5332}), .clk ( clk ), .r ( Fresh[825] ), .c ({new_AGEMA_signal_1828, n2308}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2476 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5346}), .b ({new_AGEMA_signal_1811, n2305}), .clk ( clk ), .r ( Fresh[826] ), .c ({new_AGEMA_signal_1829, n2307}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2533 ( .a ({new_AGEMA_signal_5368, new_AGEMA_signal_5360}), .b ({new_AGEMA_signal_1812, n2368}), .clk ( clk ), .r ( Fresh[827] ), .c ({new_AGEMA_signal_1830, n2370}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2611 ( .a ({new_AGEMA_signal_1814, n2457}), .b ({new_AGEMA_signal_5384, new_AGEMA_signal_5376}), .clk ( clk ), .r ( Fresh[828] ), .c ({new_AGEMA_signal_1831, n2530}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2660 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5386}), .b ({new_AGEMA_signal_1815, n2513}), .clk ( clk ), .r ( Fresh[829] ), .c ({new_AGEMA_signal_1832, n2515}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2718 ( .a ({new_AGEMA_signal_5396, new_AGEMA_signal_5392}), .b ({new_AGEMA_signal_1816, n2592}), .clk ( clk ), .r ( Fresh[830] ), .c ({new_AGEMA_signal_1833, n2639}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2749 ( .a ({new_AGEMA_signal_1793, n2637}), .b ({new_AGEMA_signal_5404, new_AGEMA_signal_5400}), .clk ( clk ), .r ( Fresh[831] ), .c ({new_AGEMA_signal_1817, n2638}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2788 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5412}), .b ({new_AGEMA_signal_1819, n2705}), .clk ( clk ), .r ( Fresh[832] ), .c ({new_AGEMA_signal_1834, n2832}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2842 ( .a ({new_AGEMA_signal_5428, new_AGEMA_signal_5424}), .b ({new_AGEMA_signal_1796, n2805}), .clk ( clk ), .r ( Fresh[833] ), .c ({new_AGEMA_signal_1820, n2807}) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C ( clk ), .D ( new_AGEMA_signal_5435 ), .Q ( new_AGEMA_signal_5436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C ( clk ), .D ( new_AGEMA_signal_5443 ), .Q ( new_AGEMA_signal_5444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C ( clk ), .D ( new_AGEMA_signal_5455 ), .Q ( new_AGEMA_signal_5456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C ( clk ), .D ( new_AGEMA_signal_5467 ), .Q ( new_AGEMA_signal_5468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C ( clk ), .D ( new_AGEMA_signal_5481 ), .Q ( new_AGEMA_signal_5482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C ( clk ), .D ( new_AGEMA_signal_5495 ), .Q ( new_AGEMA_signal_5496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C ( clk ), .D ( new_AGEMA_signal_5503 ), .Q ( new_AGEMA_signal_5504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C ( clk ), .D ( new_AGEMA_signal_5511 ), .Q ( new_AGEMA_signal_5512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C ( clk ), .D ( new_AGEMA_signal_5525 ), .Q ( new_AGEMA_signal_5526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C ( clk ), .D ( new_AGEMA_signal_5539 ), .Q ( new_AGEMA_signal_5540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C ( clk ), .D ( new_AGEMA_signal_5547 ), .Q ( new_AGEMA_signal_5548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C ( clk ), .D ( new_AGEMA_signal_5555 ), .Q ( new_AGEMA_signal_5556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C ( clk ), .D ( new_AGEMA_signal_5563 ), .Q ( new_AGEMA_signal_5564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C ( clk ), .D ( new_AGEMA_signal_5571 ), .Q ( new_AGEMA_signal_5572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C ( clk ), .D ( new_AGEMA_signal_5573 ), .Q ( new_AGEMA_signal_5574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C ( clk ), .D ( new_AGEMA_signal_5577 ), .Q ( new_AGEMA_signal_5578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C ( clk ), .D ( new_AGEMA_signal_5597 ), .Q ( new_AGEMA_signal_5598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C ( clk ), .D ( new_AGEMA_signal_5613 ), .Q ( new_AGEMA_signal_5614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C ( clk ), .D ( new_AGEMA_signal_5617 ), .Q ( new_AGEMA_signal_5618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C ( clk ), .D ( new_AGEMA_signal_5621 ), .Q ( new_AGEMA_signal_5622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C ( clk ), .D ( new_AGEMA_signal_5641 ), .Q ( new_AGEMA_signal_5642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C ( clk ), .D ( new_AGEMA_signal_5657 ), .Q ( new_AGEMA_signal_5658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C ( clk ), .D ( new_AGEMA_signal_5667 ), .Q ( new_AGEMA_signal_5668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C ( clk ), .D ( new_AGEMA_signal_5677 ), .Q ( new_AGEMA_signal_5678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C ( clk ), .D ( new_AGEMA_signal_5681 ), .Q ( new_AGEMA_signal_5682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C ( clk ), .D ( new_AGEMA_signal_5685 ), .Q ( new_AGEMA_signal_5686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C ( clk ), .D ( new_AGEMA_signal_5693 ), .Q ( new_AGEMA_signal_5694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C ( clk ), .D ( new_AGEMA_signal_5701 ), .Q ( new_AGEMA_signal_5702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C ( clk ), .D ( new_AGEMA_signal_5705 ), .Q ( new_AGEMA_signal_5706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C ( clk ), .D ( new_AGEMA_signal_5711 ), .Q ( new_AGEMA_signal_5712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C ( clk ), .D ( new_AGEMA_signal_5717 ), .Q ( new_AGEMA_signal_5718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C ( clk ), .D ( new_AGEMA_signal_5723 ), .Q ( new_AGEMA_signal_5724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C ( clk ), .D ( new_AGEMA_signal_5739 ), .Q ( new_AGEMA_signal_5740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C ( clk ), .D ( new_AGEMA_signal_5755 ), .Q ( new_AGEMA_signal_5756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C ( clk ), .D ( new_AGEMA_signal_5765 ), .Q ( new_AGEMA_signal_5766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C ( clk ), .D ( new_AGEMA_signal_5775 ), .Q ( new_AGEMA_signal_5776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C ( clk ), .D ( new_AGEMA_signal_5793 ), .Q ( new_AGEMA_signal_5794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C ( clk ), .D ( new_AGEMA_signal_5811 ), .Q ( new_AGEMA_signal_5812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C ( clk ), .D ( new_AGEMA_signal_5827 ), .Q ( new_AGEMA_signal_5828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C ( clk ), .D ( new_AGEMA_signal_5835 ), .Q ( new_AGEMA_signal_5836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C ( clk ), .D ( new_AGEMA_signal_5849 ), .Q ( new_AGEMA_signal_5850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C ( clk ), .D ( new_AGEMA_signal_5857 ), .Q ( new_AGEMA_signal_5858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C ( clk ), .D ( new_AGEMA_signal_5893 ), .Q ( new_AGEMA_signal_5894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C ( clk ), .D ( new_AGEMA_signal_5913 ), .Q ( new_AGEMA_signal_5914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C ( clk ), .D ( new_AGEMA_signal_5939 ), .Q ( new_AGEMA_signal_5940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C ( clk ), .D ( new_AGEMA_signal_5951 ), .Q ( new_AGEMA_signal_5952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C ( clk ), .D ( new_AGEMA_signal_5963 ), .Q ( new_AGEMA_signal_5964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C ( clk ), .D ( new_AGEMA_signal_5977 ), .Q ( new_AGEMA_signal_5978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C ( clk ), .D ( new_AGEMA_signal_5989 ), .Q ( new_AGEMA_signal_5990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C ( clk ), .D ( new_AGEMA_signal_6003 ), .Q ( new_AGEMA_signal_6004 ) ) ;

    /* cells in depth 21 */
    buf_clk new_AGEMA_reg_buffer_3757 ( .C ( clk ), .D ( new_AGEMA_signal_5574 ), .Q ( new_AGEMA_signal_5575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C ( clk ), .D ( new_AGEMA_signal_5578 ), .Q ( new_AGEMA_signal_5579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C ( clk ), .D ( n2109 ), .Q ( new_AGEMA_signal_5581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_5583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C ( clk ), .D ( new_AGEMA_signal_5598 ), .Q ( new_AGEMA_signal_5599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C ( clk ), .D ( new_AGEMA_signal_5614 ), .Q ( new_AGEMA_signal_5615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C ( clk ), .D ( new_AGEMA_signal_5618 ), .Q ( new_AGEMA_signal_5619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C ( clk ), .D ( new_AGEMA_signal_5622 ), .Q ( new_AGEMA_signal_5623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C ( clk ), .D ( n2310 ), .Q ( new_AGEMA_signal_5625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C ( clk ), .D ( new_AGEMA_signal_1827 ), .Q ( new_AGEMA_signal_5627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C ( clk ), .D ( new_AGEMA_signal_5642 ), .Q ( new_AGEMA_signal_5643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C ( clk ), .D ( new_AGEMA_signal_5658 ), .Q ( new_AGEMA_signal_5659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C ( clk ), .D ( new_AGEMA_signal_5668 ), .Q ( new_AGEMA_signal_5669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C ( clk ), .D ( new_AGEMA_signal_5678 ), .Q ( new_AGEMA_signal_5679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C ( clk ), .D ( new_AGEMA_signal_5682 ), .Q ( new_AGEMA_signal_5683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C ( clk ), .D ( new_AGEMA_signal_5686 ), .Q ( new_AGEMA_signal_5687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C ( clk ), .D ( new_AGEMA_signal_5694 ), .Q ( new_AGEMA_signal_5695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C ( clk ), .D ( new_AGEMA_signal_5702 ), .Q ( new_AGEMA_signal_5703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C ( clk ), .D ( new_AGEMA_signal_5706 ), .Q ( new_AGEMA_signal_5707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C ( clk ), .D ( new_AGEMA_signal_5712 ), .Q ( new_AGEMA_signal_5713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C ( clk ), .D ( new_AGEMA_signal_5718 ), .Q ( new_AGEMA_signal_5719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C ( clk ), .D ( new_AGEMA_signal_5724 ), .Q ( new_AGEMA_signal_5725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C ( clk ), .D ( new_AGEMA_signal_5740 ), .Q ( new_AGEMA_signal_5741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C ( clk ), .D ( new_AGEMA_signal_5756 ), .Q ( new_AGEMA_signal_5757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C ( clk ), .D ( new_AGEMA_signal_5766 ), .Q ( new_AGEMA_signal_5767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C ( clk ), .D ( new_AGEMA_signal_5776 ), .Q ( new_AGEMA_signal_5777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C ( clk ), .D ( new_AGEMA_signal_5794 ), .Q ( new_AGEMA_signal_5795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C ( clk ), .D ( new_AGEMA_signal_5812 ), .Q ( new_AGEMA_signal_5813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C ( clk ), .D ( n2530 ), .Q ( new_AGEMA_signal_5817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C ( clk ), .D ( new_AGEMA_signal_1831 ), .Q ( new_AGEMA_signal_5821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C ( clk ), .D ( new_AGEMA_signal_5828 ), .Q ( new_AGEMA_signal_5829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C ( clk ), .D ( new_AGEMA_signal_5836 ), .Q ( new_AGEMA_signal_5837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C ( clk ), .D ( n2832 ), .Q ( new_AGEMA_signal_5841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C ( clk ), .D ( new_AGEMA_signal_1834 ), .Q ( new_AGEMA_signal_5845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C ( clk ), .D ( new_AGEMA_signal_5850 ), .Q ( new_AGEMA_signal_5851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C ( clk ), .D ( new_AGEMA_signal_5858 ), .Q ( new_AGEMA_signal_5859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C ( clk ), .D ( n2113 ), .Q ( new_AGEMA_signal_5865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C ( clk ), .D ( new_AGEMA_signal_1801 ), .Q ( new_AGEMA_signal_5871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C ( clk ), .D ( new_AGEMA_signal_5894 ), .Q ( new_AGEMA_signal_5895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C ( clk ), .D ( new_AGEMA_signal_5914 ), .Q ( new_AGEMA_signal_5915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C ( clk ), .D ( n2212 ), .Q ( new_AGEMA_signal_5921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C ( clk ), .D ( new_AGEMA_signal_1824 ), .Q ( new_AGEMA_signal_5929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C ( clk ), .D ( new_AGEMA_signal_5940 ), .Q ( new_AGEMA_signal_5941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C ( clk ), .D ( new_AGEMA_signal_5952 ), .Q ( new_AGEMA_signal_5953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C ( clk ), .D ( new_AGEMA_signal_5964 ), .Q ( new_AGEMA_signal_5965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C ( clk ), .D ( new_AGEMA_signal_5978 ), .Q ( new_AGEMA_signal_5979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C ( clk ), .D ( new_AGEMA_signal_5990 ), .Q ( new_AGEMA_signal_5991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C ( clk ), .D ( new_AGEMA_signal_6004 ), .Q ( new_AGEMA_signal_6005 ) ) ;

    /* cells in depth 22 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2129 ( .a ({new_AGEMA_signal_1821, n2000}), .b ({new_AGEMA_signal_5444, new_AGEMA_signal_5436}), .clk ( clk ), .r ( Fresh[834] ), .c ({new_AGEMA_signal_1836, n2001}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2267 ( .a ({new_AGEMA_signal_1823, n2107}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5456}), .clk ( clk ), .r ( Fresh[835] ), .c ({new_AGEMA_signal_1837, n2108}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2317 ( .a ({new_AGEMA_signal_5496, new_AGEMA_signal_5482}), .b ({new_AGEMA_signal_1825, n2149}), .clk ( clk ), .r ( Fresh[836] ), .c ({new_AGEMA_signal_1838, n2153}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2374 ( .a ({new_AGEMA_signal_1826, n2206}), .b ({new_AGEMA_signal_5512, new_AGEMA_signal_5504}), .clk ( clk ), .r ( Fresh[837] ), .c ({new_AGEMA_signal_1839, n2207}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2477 ( .a ({new_AGEMA_signal_1828, n2308}), .b ({new_AGEMA_signal_1829, n2307}), .clk ( clk ), .r ( Fresh[838] ), .c ({new_AGEMA_signal_1840, n2309}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2535 ( .a ({new_AGEMA_signal_1830, n2370}), .b ({new_AGEMA_signal_5540, new_AGEMA_signal_5526}), .clk ( clk ), .r ( Fresh[839] ), .c ({new_AGEMA_signal_1841, n2373}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2661 ( .a ({new_AGEMA_signal_5556, new_AGEMA_signal_5548}), .b ({new_AGEMA_signal_1832, n2515}), .clk ( clk ), .r ( Fresh[840] ), .c ({new_AGEMA_signal_1842, n2528}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2750 ( .a ({new_AGEMA_signal_1833, n2639}), .b ({new_AGEMA_signal_1817, n2638}), .clk ( clk ), .r ( Fresh[841] ), .c ({new_AGEMA_signal_1843, n2669}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2843 ( .a ({new_AGEMA_signal_5572, new_AGEMA_signal_5564}), .b ({new_AGEMA_signal_1820, n2807}), .clk ( clk ), .r ( Fresh[842] ), .c ({new_AGEMA_signal_1835, n2830}) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C ( clk ), .D ( new_AGEMA_signal_5575 ), .Q ( new_AGEMA_signal_5576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C ( clk ), .D ( new_AGEMA_signal_5579 ), .Q ( new_AGEMA_signal_5580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C ( clk ), .D ( new_AGEMA_signal_5581 ), .Q ( new_AGEMA_signal_5582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C ( clk ), .D ( new_AGEMA_signal_5583 ), .Q ( new_AGEMA_signal_5584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C ( clk ), .D ( new_AGEMA_signal_5599 ), .Q ( new_AGEMA_signal_5600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C ( clk ), .D ( new_AGEMA_signal_5615 ), .Q ( new_AGEMA_signal_5616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C ( clk ), .D ( new_AGEMA_signal_5619 ), .Q ( new_AGEMA_signal_5620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C ( clk ), .D ( new_AGEMA_signal_5623 ), .Q ( new_AGEMA_signal_5624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C ( clk ), .D ( new_AGEMA_signal_5625 ), .Q ( new_AGEMA_signal_5626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C ( clk ), .D ( new_AGEMA_signal_5627 ), .Q ( new_AGEMA_signal_5628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C ( clk ), .D ( new_AGEMA_signal_5643 ), .Q ( new_AGEMA_signal_5644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C ( clk ), .D ( new_AGEMA_signal_5659 ), .Q ( new_AGEMA_signal_5660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C ( clk ), .D ( new_AGEMA_signal_5669 ), .Q ( new_AGEMA_signal_5670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C ( clk ), .D ( new_AGEMA_signal_5679 ), .Q ( new_AGEMA_signal_5680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C ( clk ), .D ( new_AGEMA_signal_5683 ), .Q ( new_AGEMA_signal_5684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C ( clk ), .D ( new_AGEMA_signal_5687 ), .Q ( new_AGEMA_signal_5688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C ( clk ), .D ( new_AGEMA_signal_5695 ), .Q ( new_AGEMA_signal_5696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C ( clk ), .D ( new_AGEMA_signal_5703 ), .Q ( new_AGEMA_signal_5704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C ( clk ), .D ( new_AGEMA_signal_5707 ), .Q ( new_AGEMA_signal_5708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C ( clk ), .D ( new_AGEMA_signal_5713 ), .Q ( new_AGEMA_signal_5714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C ( clk ), .D ( new_AGEMA_signal_5719 ), .Q ( new_AGEMA_signal_5720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C ( clk ), .D ( new_AGEMA_signal_5725 ), .Q ( new_AGEMA_signal_5726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C ( clk ), .D ( new_AGEMA_signal_5741 ), .Q ( new_AGEMA_signal_5742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C ( clk ), .D ( new_AGEMA_signal_5757 ), .Q ( new_AGEMA_signal_5758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C ( clk ), .D ( new_AGEMA_signal_5767 ), .Q ( new_AGEMA_signal_5768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C ( clk ), .D ( new_AGEMA_signal_5777 ), .Q ( new_AGEMA_signal_5778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C ( clk ), .D ( new_AGEMA_signal_5795 ), .Q ( new_AGEMA_signal_5796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C ( clk ), .D ( new_AGEMA_signal_5813 ), .Q ( new_AGEMA_signal_5814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C ( clk ), .D ( new_AGEMA_signal_5817 ), .Q ( new_AGEMA_signal_5818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C ( clk ), .D ( new_AGEMA_signal_5821 ), .Q ( new_AGEMA_signal_5822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C ( clk ), .D ( new_AGEMA_signal_5829 ), .Q ( new_AGEMA_signal_5830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C ( clk ), .D ( new_AGEMA_signal_5837 ), .Q ( new_AGEMA_signal_5838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C ( clk ), .D ( new_AGEMA_signal_5841 ), .Q ( new_AGEMA_signal_5842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C ( clk ), .D ( new_AGEMA_signal_5845 ), .Q ( new_AGEMA_signal_5846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C ( clk ), .D ( new_AGEMA_signal_5851 ), .Q ( new_AGEMA_signal_5852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C ( clk ), .D ( new_AGEMA_signal_5859 ), .Q ( new_AGEMA_signal_5860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C ( clk ), .D ( new_AGEMA_signal_5865 ), .Q ( new_AGEMA_signal_5866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C ( clk ), .D ( new_AGEMA_signal_5871 ), .Q ( new_AGEMA_signal_5872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C ( clk ), .D ( new_AGEMA_signal_5895 ), .Q ( new_AGEMA_signal_5896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C ( clk ), .D ( new_AGEMA_signal_5915 ), .Q ( new_AGEMA_signal_5916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C ( clk ), .D ( new_AGEMA_signal_5921 ), .Q ( new_AGEMA_signal_5922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C ( clk ), .D ( new_AGEMA_signal_5929 ), .Q ( new_AGEMA_signal_5930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C ( clk ), .D ( new_AGEMA_signal_5941 ), .Q ( new_AGEMA_signal_5942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C ( clk ), .D ( new_AGEMA_signal_5953 ), .Q ( new_AGEMA_signal_5954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C ( clk ), .D ( new_AGEMA_signal_5965 ), .Q ( new_AGEMA_signal_5966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C ( clk ), .D ( new_AGEMA_signal_5979 ), .Q ( new_AGEMA_signal_5980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C ( clk ), .D ( new_AGEMA_signal_5991 ), .Q ( new_AGEMA_signal_5992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C ( clk ), .D ( new_AGEMA_signal_6005 ), .Q ( new_AGEMA_signal_6006 ) ) ;

    /* cells in depth 23 */
    buf_clk new_AGEMA_reg_buffer_3891 ( .C ( clk ), .D ( new_AGEMA_signal_5708 ), .Q ( new_AGEMA_signal_5709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C ( clk ), .D ( new_AGEMA_signal_5714 ), .Q ( new_AGEMA_signal_5715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C ( clk ), .D ( new_AGEMA_signal_5720 ), .Q ( new_AGEMA_signal_5721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C ( clk ), .D ( new_AGEMA_signal_5726 ), .Q ( new_AGEMA_signal_5727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C ( clk ), .D ( new_AGEMA_signal_5742 ), .Q ( new_AGEMA_signal_5743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C ( clk ), .D ( new_AGEMA_signal_5758 ), .Q ( new_AGEMA_signal_5759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C ( clk ), .D ( new_AGEMA_signal_5768 ), .Q ( new_AGEMA_signal_5769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C ( clk ), .D ( new_AGEMA_signal_5778 ), .Q ( new_AGEMA_signal_5779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C ( clk ), .D ( new_AGEMA_signal_5796 ), .Q ( new_AGEMA_signal_5797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C ( clk ), .D ( new_AGEMA_signal_5814 ), .Q ( new_AGEMA_signal_5815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C ( clk ), .D ( new_AGEMA_signal_5818 ), .Q ( new_AGEMA_signal_5819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C ( clk ), .D ( new_AGEMA_signal_5822 ), .Q ( new_AGEMA_signal_5823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C ( clk ), .D ( new_AGEMA_signal_5830 ), .Q ( new_AGEMA_signal_5831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C ( clk ), .D ( new_AGEMA_signal_5838 ), .Q ( new_AGEMA_signal_5839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C ( clk ), .D ( new_AGEMA_signal_5842 ), .Q ( new_AGEMA_signal_5843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C ( clk ), .D ( new_AGEMA_signal_5846 ), .Q ( new_AGEMA_signal_5847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C ( clk ), .D ( new_AGEMA_signal_5852 ), .Q ( new_AGEMA_signal_5853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C ( clk ), .D ( new_AGEMA_signal_5860 ), .Q ( new_AGEMA_signal_5861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C ( clk ), .D ( new_AGEMA_signal_5866 ), .Q ( new_AGEMA_signal_5867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C ( clk ), .D ( new_AGEMA_signal_5872 ), .Q ( new_AGEMA_signal_5873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C ( clk ), .D ( new_AGEMA_signal_5896 ), .Q ( new_AGEMA_signal_5897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C ( clk ), .D ( new_AGEMA_signal_5916 ), .Q ( new_AGEMA_signal_5917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C ( clk ), .D ( new_AGEMA_signal_5922 ), .Q ( new_AGEMA_signal_5923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C ( clk ), .D ( new_AGEMA_signal_5930 ), .Q ( new_AGEMA_signal_5931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C ( clk ), .D ( new_AGEMA_signal_5942 ), .Q ( new_AGEMA_signal_5943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C ( clk ), .D ( new_AGEMA_signal_5954 ), .Q ( new_AGEMA_signal_5955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C ( clk ), .D ( new_AGEMA_signal_5966 ), .Q ( new_AGEMA_signal_5967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C ( clk ), .D ( new_AGEMA_signal_5980 ), .Q ( new_AGEMA_signal_5981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C ( clk ), .D ( new_AGEMA_signal_5992 ), .Q ( new_AGEMA_signal_5993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C ( clk ), .D ( new_AGEMA_signal_6006 ), .Q ( new_AGEMA_signal_6007 ) ) ;

    /* cells in depth 24 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2130 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5576}), .b ({new_AGEMA_signal_1836, n2001}), .clk ( clk ), .r ( Fresh[843] ), .c ({new_AGEMA_signal_1845, n2017}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2268 ( .a ({new_AGEMA_signal_5584, new_AGEMA_signal_5582}), .b ({new_AGEMA_signal_1837, n2108}), .clk ( clk ), .r ( Fresh[844] ), .c ({new_AGEMA_signal_1846, n2110}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2319 ( .a ({new_AGEMA_signal_1838, n2153}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5600}), .clk ( clk ), .r ( Fresh[845] ), .c ({new_AGEMA_signal_1847, n2154}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2375 ( .a ({new_AGEMA_signal_5624, new_AGEMA_signal_5620}), .b ({new_AGEMA_signal_1839, n2207}), .clk ( clk ), .r ( Fresh[846] ), .c ({new_AGEMA_signal_1848, n2209}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2478 ( .a ({new_AGEMA_signal_5628, new_AGEMA_signal_5626}), .b ({new_AGEMA_signal_1840, n2309}), .clk ( clk ), .r ( Fresh[847] ), .c ({new_AGEMA_signal_1849, n2311}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2537 ( .a ({new_AGEMA_signal_1841, n2373}), .b ({new_AGEMA_signal_5660, new_AGEMA_signal_5644}), .clk ( clk ), .r ( Fresh[848] ), .c ({new_AGEMA_signal_1850, n2374}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2672 ( .a ({new_AGEMA_signal_1842, n2528}), .b ({new_AGEMA_signal_5680, new_AGEMA_signal_5670}), .clk ( clk ), .r ( Fresh[849] ), .c ({new_AGEMA_signal_1851, n2529}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2768 ( .a ({new_AGEMA_signal_1843, n2669}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5684}), .clk ( clk ), .r ( Fresh[850] ), .c ({new_AGEMA_signal_1852, n2670}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2854 ( .a ({new_AGEMA_signal_1835, n2830}), .b ({new_AGEMA_signal_5704, new_AGEMA_signal_5696}), .clk ( clk ), .r ( Fresh[851] ), .c ({new_AGEMA_signal_1844, n2831}) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C ( clk ), .D ( new_AGEMA_signal_5709 ), .Q ( new_AGEMA_signal_5710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C ( clk ), .D ( new_AGEMA_signal_5715 ), .Q ( new_AGEMA_signal_5716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C ( clk ), .D ( new_AGEMA_signal_5721 ), .Q ( new_AGEMA_signal_5722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C ( clk ), .D ( new_AGEMA_signal_5727 ), .Q ( new_AGEMA_signal_5728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C ( clk ), .D ( new_AGEMA_signal_5743 ), .Q ( new_AGEMA_signal_5744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C ( clk ), .D ( new_AGEMA_signal_5759 ), .Q ( new_AGEMA_signal_5760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C ( clk ), .D ( new_AGEMA_signal_5769 ), .Q ( new_AGEMA_signal_5770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C ( clk ), .D ( new_AGEMA_signal_5779 ), .Q ( new_AGEMA_signal_5780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C ( clk ), .D ( new_AGEMA_signal_5797 ), .Q ( new_AGEMA_signal_5798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C ( clk ), .D ( new_AGEMA_signal_5815 ), .Q ( new_AGEMA_signal_5816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C ( clk ), .D ( new_AGEMA_signal_5819 ), .Q ( new_AGEMA_signal_5820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C ( clk ), .D ( new_AGEMA_signal_5823 ), .Q ( new_AGEMA_signal_5824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C ( clk ), .D ( new_AGEMA_signal_5831 ), .Q ( new_AGEMA_signal_5832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C ( clk ), .D ( new_AGEMA_signal_5839 ), .Q ( new_AGEMA_signal_5840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C ( clk ), .D ( new_AGEMA_signal_5843 ), .Q ( new_AGEMA_signal_5844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C ( clk ), .D ( new_AGEMA_signal_5847 ), .Q ( new_AGEMA_signal_5848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C ( clk ), .D ( new_AGEMA_signal_5853 ), .Q ( new_AGEMA_signal_5854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C ( clk ), .D ( new_AGEMA_signal_5861 ), .Q ( new_AGEMA_signal_5862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C ( clk ), .D ( new_AGEMA_signal_5867 ), .Q ( new_AGEMA_signal_5868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C ( clk ), .D ( new_AGEMA_signal_5873 ), .Q ( new_AGEMA_signal_5874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C ( clk ), .D ( new_AGEMA_signal_5897 ), .Q ( new_AGEMA_signal_5898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C ( clk ), .D ( new_AGEMA_signal_5917 ), .Q ( new_AGEMA_signal_5918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C ( clk ), .D ( new_AGEMA_signal_5923 ), .Q ( new_AGEMA_signal_5924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C ( clk ), .D ( new_AGEMA_signal_5931 ), .Q ( new_AGEMA_signal_5932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C ( clk ), .D ( new_AGEMA_signal_5943 ), .Q ( new_AGEMA_signal_5944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C ( clk ), .D ( new_AGEMA_signal_5955 ), .Q ( new_AGEMA_signal_5956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C ( clk ), .D ( new_AGEMA_signal_5967 ), .Q ( new_AGEMA_signal_5968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C ( clk ), .D ( new_AGEMA_signal_5981 ), .Q ( new_AGEMA_signal_5982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C ( clk ), .D ( new_AGEMA_signal_5993 ), .Q ( new_AGEMA_signal_5994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C ( clk ), .D ( new_AGEMA_signal_6007 ), .Q ( new_AGEMA_signal_6008 ) ) ;

    /* cells in depth 25 */
    buf_clk new_AGEMA_reg_buffer_4037 ( .C ( clk ), .D ( new_AGEMA_signal_5854 ), .Q ( new_AGEMA_signal_5855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C ( clk ), .D ( new_AGEMA_signal_5862 ), .Q ( new_AGEMA_signal_5863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C ( clk ), .D ( new_AGEMA_signal_5868 ), .Q ( new_AGEMA_signal_5869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C ( clk ), .D ( new_AGEMA_signal_5874 ), .Q ( new_AGEMA_signal_5875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C ( clk ), .D ( n2209 ), .Q ( new_AGEMA_signal_5877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C ( clk ), .D ( new_AGEMA_signal_1848 ), .Q ( new_AGEMA_signal_5879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C ( clk ), .D ( new_AGEMA_signal_5898 ), .Q ( new_AGEMA_signal_5899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C ( clk ), .D ( new_AGEMA_signal_5918 ), .Q ( new_AGEMA_signal_5919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C ( clk ), .D ( new_AGEMA_signal_5924 ), .Q ( new_AGEMA_signal_5925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C ( clk ), .D ( new_AGEMA_signal_5932 ), .Q ( new_AGEMA_signal_5933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C ( clk ), .D ( new_AGEMA_signal_5944 ), .Q ( new_AGEMA_signal_5945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C ( clk ), .D ( new_AGEMA_signal_5956 ), .Q ( new_AGEMA_signal_5957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C ( clk ), .D ( new_AGEMA_signal_5968 ), .Q ( new_AGEMA_signal_5969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C ( clk ), .D ( new_AGEMA_signal_5982 ), .Q ( new_AGEMA_signal_5983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C ( clk ), .D ( new_AGEMA_signal_5994 ), .Q ( new_AGEMA_signal_5995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C ( clk ), .D ( new_AGEMA_signal_6008 ), .Q ( new_AGEMA_signal_6009 ) ) ;

    /* cells in depth 26 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2155 ( .a ({new_AGEMA_signal_1845, n2017}), .b ({new_AGEMA_signal_5716, new_AGEMA_signal_5710}), .clk ( clk ), .r ( Fresh[852] ), .c ({new_AGEMA_signal_1854, n2018}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2269 ( .a ({new_AGEMA_signal_5728, new_AGEMA_signal_5722}), .b ({new_AGEMA_signal_1846, n2110}), .clk ( clk ), .r ( Fresh[853] ), .c ({new_AGEMA_signal_1855, n2112}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2320 ( .a ({new_AGEMA_signal_5760, new_AGEMA_signal_5744}), .b ({new_AGEMA_signal_1847, n2154}), .clk ( clk ), .r ( Fresh[854] ), .c ({new_AGEMA_signal_1856, n2210}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2479 ( .a ({new_AGEMA_signal_5780, new_AGEMA_signal_5770}), .b ({new_AGEMA_signal_1849, n2311}), .clk ( clk ), .r ( Fresh[855] ), .c ({new_AGEMA_signal_1857, N470}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2538 ( .a ({new_AGEMA_signal_5816, new_AGEMA_signal_5798}), .b ({new_AGEMA_signal_1850, n2374}), .clk ( clk ), .r ( Fresh[856] ), .c ({new_AGEMA_signal_1858, n2378}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2673 ( .a ({new_AGEMA_signal_5824, new_AGEMA_signal_5820}), .b ({new_AGEMA_signal_1851, n2529}), .clk ( clk ), .r ( Fresh[857] ), .c ({new_AGEMA_signal_1859, N639}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2769 ( .a ({new_AGEMA_signal_5840, new_AGEMA_signal_5832}), .b ({new_AGEMA_signal_1852, n2670}), .clk ( clk ), .r ( Fresh[858] ), .c ({new_AGEMA_signal_1860, N723}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2855 ( .a ({new_AGEMA_signal_5848, new_AGEMA_signal_5844}), .b ({new_AGEMA_signal_1844, n2831}), .clk ( clk ), .r ( Fresh[859] ), .c ({new_AGEMA_signal_1853, N789}) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C ( clk ), .D ( new_AGEMA_signal_5855 ), .Q ( new_AGEMA_signal_5856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C ( clk ), .D ( new_AGEMA_signal_5863 ), .Q ( new_AGEMA_signal_5864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C ( clk ), .D ( new_AGEMA_signal_5869 ), .Q ( new_AGEMA_signal_5870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C ( clk ), .D ( new_AGEMA_signal_5875 ), .Q ( new_AGEMA_signal_5876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C ( clk ), .D ( new_AGEMA_signal_5877 ), .Q ( new_AGEMA_signal_5878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C ( clk ), .D ( new_AGEMA_signal_5879 ), .Q ( new_AGEMA_signal_5880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C ( clk ), .D ( new_AGEMA_signal_5899 ), .Q ( new_AGEMA_signal_5900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C ( clk ), .D ( new_AGEMA_signal_5919 ), .Q ( new_AGEMA_signal_5920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C ( clk ), .D ( new_AGEMA_signal_5925 ), .Q ( new_AGEMA_signal_5926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C ( clk ), .D ( new_AGEMA_signal_5933 ), .Q ( new_AGEMA_signal_5934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C ( clk ), .D ( new_AGEMA_signal_5945 ), .Q ( new_AGEMA_signal_5946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C ( clk ), .D ( new_AGEMA_signal_5957 ), .Q ( new_AGEMA_signal_5958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C ( clk ), .D ( new_AGEMA_signal_5969 ), .Q ( new_AGEMA_signal_5970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C ( clk ), .D ( new_AGEMA_signal_5983 ), .Q ( new_AGEMA_signal_5984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C ( clk ), .D ( new_AGEMA_signal_5995 ), .Q ( new_AGEMA_signal_5996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C ( clk ), .D ( new_AGEMA_signal_6009 ), .Q ( new_AGEMA_signal_6010 ) ) ;

    /* cells in depth 27 */
    buf_clk new_AGEMA_reg_buffer_4109 ( .C ( clk ), .D ( new_AGEMA_signal_5926 ), .Q ( new_AGEMA_signal_5927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C ( clk ), .D ( new_AGEMA_signal_5934 ), .Q ( new_AGEMA_signal_5935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C ( clk ), .D ( new_AGEMA_signal_5946 ), .Q ( new_AGEMA_signal_5947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C ( clk ), .D ( new_AGEMA_signal_5958 ), .Q ( new_AGEMA_signal_5959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C ( clk ), .D ( new_AGEMA_signal_5970 ), .Q ( new_AGEMA_signal_5971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C ( clk ), .D ( new_AGEMA_signal_5984 ), .Q ( new_AGEMA_signal_5985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C ( clk ), .D ( new_AGEMA_signal_5996 ), .Q ( new_AGEMA_signal_5997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C ( clk ), .D ( new_AGEMA_signal_6010 ), .Q ( new_AGEMA_signal_6011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C ( clk ), .D ( N470 ), .Q ( new_AGEMA_signal_6049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C ( clk ), .D ( new_AGEMA_signal_1857 ), .Q ( new_AGEMA_signal_6057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C ( clk ), .D ( N639 ), .Q ( new_AGEMA_signal_6065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C ( clk ), .D ( new_AGEMA_signal_1859 ), .Q ( new_AGEMA_signal_6073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C ( clk ), .D ( N723 ), .Q ( new_AGEMA_signal_6081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C ( clk ), .D ( new_AGEMA_signal_1860 ), .Q ( new_AGEMA_signal_6089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C ( clk ), .D ( N789 ), .Q ( new_AGEMA_signal_6097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_6105 ) ) ;

    /* cells in depth 28 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2156 ( .a ({new_AGEMA_signal_5864, new_AGEMA_signal_5856}), .b ({new_AGEMA_signal_1854, n2018}), .clk ( clk ), .r ( Fresh[860] ), .c ({new_AGEMA_signal_1861, N169}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2270 ( .a ({new_AGEMA_signal_5876, new_AGEMA_signal_5870}), .b ({new_AGEMA_signal_1855, n2112}), .clk ( clk ), .r ( Fresh[861] ), .c ({new_AGEMA_signal_1862, N277}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2376 ( .a ({new_AGEMA_signal_1856, n2210}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5878}), .clk ( clk ), .r ( Fresh[862] ), .c ({new_AGEMA_signal_1863, n2211}) ) ;
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2540 ( .a ({new_AGEMA_signal_1858, n2378}), .b ({new_AGEMA_signal_5920, new_AGEMA_signal_5900}), .clk ( clk ), .r ( Fresh[863] ), .c ({new_AGEMA_signal_1864, n2379}) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C ( clk ), .D ( new_AGEMA_signal_5927 ), .Q ( new_AGEMA_signal_5928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C ( clk ), .D ( new_AGEMA_signal_5935 ), .Q ( new_AGEMA_signal_5936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C ( clk ), .D ( new_AGEMA_signal_5947 ), .Q ( new_AGEMA_signal_5948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C ( clk ), .D ( new_AGEMA_signal_5959 ), .Q ( new_AGEMA_signal_5960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C ( clk ), .D ( new_AGEMA_signal_5971 ), .Q ( new_AGEMA_signal_5972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C ( clk ), .D ( new_AGEMA_signal_5985 ), .Q ( new_AGEMA_signal_5986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C ( clk ), .D ( new_AGEMA_signal_5997 ), .Q ( new_AGEMA_signal_5998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C ( clk ), .D ( new_AGEMA_signal_6011 ), .Q ( new_AGEMA_signal_6012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C ( clk ), .D ( new_AGEMA_signal_6049 ), .Q ( new_AGEMA_signal_6050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C ( clk ), .D ( new_AGEMA_signal_6057 ), .Q ( new_AGEMA_signal_6058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C ( clk ), .D ( new_AGEMA_signal_6065 ), .Q ( new_AGEMA_signal_6066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C ( clk ), .D ( new_AGEMA_signal_6073 ), .Q ( new_AGEMA_signal_6074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C ( clk ), .D ( new_AGEMA_signal_6081 ), .Q ( new_AGEMA_signal_6082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C ( clk ), .D ( new_AGEMA_signal_6089 ), .Q ( new_AGEMA_signal_6090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C ( clk ), .D ( new_AGEMA_signal_6097 ), .Q ( new_AGEMA_signal_6098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C ( clk ), .D ( new_AGEMA_signal_6105 ), .Q ( new_AGEMA_signal_6106 ) ) ;

    /* cells in depth 29 */
    buf_clk new_AGEMA_reg_buffer_4155 ( .C ( clk ), .D ( new_AGEMA_signal_5972 ), .Q ( new_AGEMA_signal_5973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C ( clk ), .D ( new_AGEMA_signal_5986 ), .Q ( new_AGEMA_signal_5987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C ( clk ), .D ( new_AGEMA_signal_5998 ), .Q ( new_AGEMA_signal_5999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C ( clk ), .D ( new_AGEMA_signal_6012 ), .Q ( new_AGEMA_signal_6013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C ( clk ), .D ( N169 ), .Q ( new_AGEMA_signal_6017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C ( clk ), .D ( new_AGEMA_signal_1861 ), .Q ( new_AGEMA_signal_6023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C ( clk ), .D ( N277 ), .Q ( new_AGEMA_signal_6029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C ( clk ), .D ( new_AGEMA_signal_1862 ), .Q ( new_AGEMA_signal_6035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C ( clk ), .D ( new_AGEMA_signal_6050 ), .Q ( new_AGEMA_signal_6051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C ( clk ), .D ( new_AGEMA_signal_6058 ), .Q ( new_AGEMA_signal_6059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C ( clk ), .D ( new_AGEMA_signal_6066 ), .Q ( new_AGEMA_signal_6067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C ( clk ), .D ( new_AGEMA_signal_6074 ), .Q ( new_AGEMA_signal_6075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C ( clk ), .D ( new_AGEMA_signal_6082 ), .Q ( new_AGEMA_signal_6083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C ( clk ), .D ( new_AGEMA_signal_6090 ), .Q ( new_AGEMA_signal_6091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C ( clk ), .D ( new_AGEMA_signal_6098 ), .Q ( new_AGEMA_signal_6099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C ( clk ), .D ( new_AGEMA_signal_6106 ), .Q ( new_AGEMA_signal_6107 ) ) ;

    /* cells in depth 30 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2377 ( .a ({new_AGEMA_signal_5936, new_AGEMA_signal_5928}), .b ({new_AGEMA_signal_1863, n2211}), .clk ( clk ), .r ( Fresh[864] ), .c ({new_AGEMA_signal_1865, N379}) ) ;
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2541 ( .a ({new_AGEMA_signal_5960, new_AGEMA_signal_5948}), .b ({new_AGEMA_signal_1864, n2379}), .clk ( clk ), .r ( Fresh[865] ), .c ({new_AGEMA_signal_1866, n2381}) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C ( clk ), .D ( new_AGEMA_signal_5973 ), .Q ( new_AGEMA_signal_5974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C ( clk ), .D ( new_AGEMA_signal_5987 ), .Q ( new_AGEMA_signal_5988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C ( clk ), .D ( new_AGEMA_signal_5999 ), .Q ( new_AGEMA_signal_6000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C ( clk ), .D ( new_AGEMA_signal_6013 ), .Q ( new_AGEMA_signal_6014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C ( clk ), .D ( new_AGEMA_signal_6017 ), .Q ( new_AGEMA_signal_6018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C ( clk ), .D ( new_AGEMA_signal_6023 ), .Q ( new_AGEMA_signal_6024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C ( clk ), .D ( new_AGEMA_signal_6029 ), .Q ( new_AGEMA_signal_6030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C ( clk ), .D ( new_AGEMA_signal_6035 ), .Q ( new_AGEMA_signal_6036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C ( clk ), .D ( new_AGEMA_signal_6051 ), .Q ( new_AGEMA_signal_6052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C ( clk ), .D ( new_AGEMA_signal_6059 ), .Q ( new_AGEMA_signal_6060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C ( clk ), .D ( new_AGEMA_signal_6067 ), .Q ( new_AGEMA_signal_6068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C ( clk ), .D ( new_AGEMA_signal_6075 ), .Q ( new_AGEMA_signal_6076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C ( clk ), .D ( new_AGEMA_signal_6083 ), .Q ( new_AGEMA_signal_6084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C ( clk ), .D ( new_AGEMA_signal_6091 ), .Q ( new_AGEMA_signal_6092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C ( clk ), .D ( new_AGEMA_signal_6099 ), .Q ( new_AGEMA_signal_6100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C ( clk ), .D ( new_AGEMA_signal_6107 ), .Q ( new_AGEMA_signal_6108 ) ) ;

    /* cells in depth 31 */
    buf_clk new_AGEMA_reg_buffer_4183 ( .C ( clk ), .D ( new_AGEMA_signal_6000 ), .Q ( new_AGEMA_signal_6001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C ( clk ), .D ( new_AGEMA_signal_6014 ), .Q ( new_AGEMA_signal_6015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C ( clk ), .D ( new_AGEMA_signal_6018 ), .Q ( new_AGEMA_signal_6019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C ( clk ), .D ( new_AGEMA_signal_6024 ), .Q ( new_AGEMA_signal_6025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C ( clk ), .D ( new_AGEMA_signal_6030 ), .Q ( new_AGEMA_signal_6031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C ( clk ), .D ( new_AGEMA_signal_6036 ), .Q ( new_AGEMA_signal_6037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C ( clk ), .D ( N379 ), .Q ( new_AGEMA_signal_6041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_6045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C ( clk ), .D ( new_AGEMA_signal_6052 ), .Q ( new_AGEMA_signal_6053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C ( clk ), .D ( new_AGEMA_signal_6060 ), .Q ( new_AGEMA_signal_6061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C ( clk ), .D ( new_AGEMA_signal_6068 ), .Q ( new_AGEMA_signal_6069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C ( clk ), .D ( new_AGEMA_signal_6076 ), .Q ( new_AGEMA_signal_6077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C ( clk ), .D ( new_AGEMA_signal_6084 ), .Q ( new_AGEMA_signal_6085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C ( clk ), .D ( new_AGEMA_signal_6092 ), .Q ( new_AGEMA_signal_6093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C ( clk ), .D ( new_AGEMA_signal_6100 ), .Q ( new_AGEMA_signal_6101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C ( clk ), .D ( new_AGEMA_signal_6108 ), .Q ( new_AGEMA_signal_6109 ) ) ;

    /* cells in depth 32 */
    nor_HPC2 #(.security_order(1), .pipeline(1)) U2542 ( .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5974}), .b ({new_AGEMA_signal_1866, n2381}), .clk ( clk ), .r ( Fresh[866] ), .c ({new_AGEMA_signal_1867, n2427}) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C ( clk ), .D ( new_AGEMA_signal_6001 ), .Q ( new_AGEMA_signal_6002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C ( clk ), .D ( new_AGEMA_signal_6015 ), .Q ( new_AGEMA_signal_6016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C ( clk ), .D ( new_AGEMA_signal_6019 ), .Q ( new_AGEMA_signal_6020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C ( clk ), .D ( new_AGEMA_signal_6025 ), .Q ( new_AGEMA_signal_6026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C ( clk ), .D ( new_AGEMA_signal_6031 ), .Q ( new_AGEMA_signal_6032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C ( clk ), .D ( new_AGEMA_signal_6037 ), .Q ( new_AGEMA_signal_6038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C ( clk ), .D ( new_AGEMA_signal_6041 ), .Q ( new_AGEMA_signal_6042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C ( clk ), .D ( new_AGEMA_signal_6045 ), .Q ( new_AGEMA_signal_6046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C ( clk ), .D ( new_AGEMA_signal_6053 ), .Q ( new_AGEMA_signal_6054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C ( clk ), .D ( new_AGEMA_signal_6061 ), .Q ( new_AGEMA_signal_6062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C ( clk ), .D ( new_AGEMA_signal_6069 ), .Q ( new_AGEMA_signal_6070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C ( clk ), .D ( new_AGEMA_signal_6077 ), .Q ( new_AGEMA_signal_6078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C ( clk ), .D ( new_AGEMA_signal_6085 ), .Q ( new_AGEMA_signal_6086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C ( clk ), .D ( new_AGEMA_signal_6093 ), .Q ( new_AGEMA_signal_6094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C ( clk ), .D ( new_AGEMA_signal_6101 ), .Q ( new_AGEMA_signal_6102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C ( clk ), .D ( new_AGEMA_signal_6109 ), .Q ( new_AGEMA_signal_6110 ) ) ;

    /* cells in depth 33 */
    buf_clk new_AGEMA_reg_buffer_4203 ( .C ( clk ), .D ( new_AGEMA_signal_6020 ), .Q ( new_AGEMA_signal_6021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C ( clk ), .D ( new_AGEMA_signal_6026 ), .Q ( new_AGEMA_signal_6027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C ( clk ), .D ( new_AGEMA_signal_6032 ), .Q ( new_AGEMA_signal_6033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C ( clk ), .D ( new_AGEMA_signal_6038 ), .Q ( new_AGEMA_signal_6039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C ( clk ), .D ( new_AGEMA_signal_6042 ), .Q ( new_AGEMA_signal_6043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C ( clk ), .D ( new_AGEMA_signal_6046 ), .Q ( new_AGEMA_signal_6047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C ( clk ), .D ( new_AGEMA_signal_6054 ), .Q ( new_AGEMA_signal_6055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C ( clk ), .D ( new_AGEMA_signal_6062 ), .Q ( new_AGEMA_signal_6063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C ( clk ), .D ( new_AGEMA_signal_6070 ), .Q ( new_AGEMA_signal_6071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C ( clk ), .D ( new_AGEMA_signal_6078 ), .Q ( new_AGEMA_signal_6079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C ( clk ), .D ( new_AGEMA_signal_6086 ), .Q ( new_AGEMA_signal_6087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C ( clk ), .D ( new_AGEMA_signal_6094 ), .Q ( new_AGEMA_signal_6095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C ( clk ), .D ( new_AGEMA_signal_6102 ), .Q ( new_AGEMA_signal_6103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C ( clk ), .D ( new_AGEMA_signal_6110 ), .Q ( new_AGEMA_signal_6111 ) ) ;

    /* cells in depth 34 */
    nand_HPC2 #(.security_order(1), .pipeline(1)) U2584 ( .a ({new_AGEMA_signal_1867, n2427}), .b ({new_AGEMA_signal_6016, new_AGEMA_signal_6002}), .clk ( clk ), .r ( Fresh[867] ), .c ({new_AGEMA_signal_1868, N563}) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C ( clk ), .D ( new_AGEMA_signal_6021 ), .Q ( new_AGEMA_signal_6022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C ( clk ), .D ( new_AGEMA_signal_6027 ), .Q ( new_AGEMA_signal_6028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C ( clk ), .D ( new_AGEMA_signal_6033 ), .Q ( new_AGEMA_signal_6034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C ( clk ), .D ( new_AGEMA_signal_6039 ), .Q ( new_AGEMA_signal_6040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C ( clk ), .D ( new_AGEMA_signal_6043 ), .Q ( new_AGEMA_signal_6044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C ( clk ), .D ( new_AGEMA_signal_6047 ), .Q ( new_AGEMA_signal_6048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C ( clk ), .D ( new_AGEMA_signal_6055 ), .Q ( new_AGEMA_signal_6056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C ( clk ), .D ( new_AGEMA_signal_6063 ), .Q ( new_AGEMA_signal_6064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C ( clk ), .D ( new_AGEMA_signal_6071 ), .Q ( new_AGEMA_signal_6072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C ( clk ), .D ( new_AGEMA_signal_6079 ), .Q ( new_AGEMA_signal_6080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C ( clk ), .D ( new_AGEMA_signal_6087 ), .Q ( new_AGEMA_signal_6088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C ( clk ), .D ( new_AGEMA_signal_6095 ), .Q ( new_AGEMA_signal_6096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C ( clk ), .D ( new_AGEMA_signal_6103 ), .Q ( new_AGEMA_signal_6104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C ( clk ), .D ( new_AGEMA_signal_6111 ), .Q ( new_AGEMA_signal_6112 ) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_6028, new_AGEMA_signal_6022}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_6040, new_AGEMA_signal_6034}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_6048, new_AGEMA_signal_6044}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_6064, new_AGEMA_signal_6056}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_1868, N563}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_6080, new_AGEMA_signal_6072}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_6096, new_AGEMA_signal_6088}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_6112, new_AGEMA_signal_6104}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
