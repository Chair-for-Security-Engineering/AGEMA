/* modified netlist. Source: module SkinnyTop in file Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module SkinnyTop_GHPC_ANF_ClockGating_d1 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output Synch ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_943 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1485 ;
    wire signal_1487 ;
    wire signal_1489 ;
    wire signal_1491 ;
    wire signal_1493 ;
    wire signal_1495 ;
    wire signal_1497 ;
    wire signal_1499 ;
    wire signal_1501 ;
    wire signal_1503 ;
    wire signal_1505 ;
    wire signal_1507 ;
    wire signal_1509 ;
    wire signal_1511 ;
    wire signal_1513 ;
    wire signal_1515 ;
    wire signal_1517 ;
    wire signal_1519 ;
    wire signal_1521 ;
    wire signal_1523 ;
    wire signal_1525 ;
    wire signal_1527 ;
    wire signal_1529 ;
    wire signal_1531 ;
    wire signal_1533 ;
    wire signal_1535 ;
    wire signal_1537 ;
    wire signal_1539 ;
    wire signal_1541 ;
    wire signal_1543 ;
    wire signal_1545 ;
    wire signal_1547 ;
    wire signal_1549 ;
    wire signal_1551 ;
    wire signal_1553 ;
    wire signal_1555 ;
    wire signal_1557 ;
    wire signal_1559 ;
    wire signal_1561 ;
    wire signal_1563 ;
    wire signal_1565 ;
    wire signal_1567 ;
    wire signal_1569 ;
    wire signal_1571 ;
    wire signal_1573 ;
    wire signal_1575 ;
    wire signal_1577 ;
    wire signal_1579 ;
    wire signal_1581 ;
    wire signal_1583 ;
    wire signal_1585 ;
    wire signal_1587 ;
    wire signal_1589 ;
    wire signal_1591 ;
    wire signal_1593 ;
    wire signal_1595 ;
    wire signal_1597 ;
    wire signal_1599 ;
    wire signal_1601 ;
    wire signal_1603 ;
    wire signal_1605 ;
    wire signal_1607 ;
    wire signal_1609 ;
    wire signal_1611 ;
    wire signal_1676 ;

    /* cells in depth 0 */
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_769 ( .s (rst), .b ({signal_1164, signal_1163}), .a ({Key_s1[0], Key_s0[0]}), .c ({signal_1166, signal_1099}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_770 ( .s (rst), .b ({signal_1167, signal_1162}), .a ({Key_s1[1], Key_s0[1]}), .c ({signal_1169, signal_1098}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_771 ( .s (rst), .b ({signal_1170, signal_1161}), .a ({Key_s1[2], Key_s0[2]}), .c ({signal_1172, signal_1097}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_772 ( .s (rst), .b ({signal_1173, signal_1160}), .a ({Key_s1[3], Key_s0[3]}), .c ({signal_1175, signal_1096}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_773 ( .s (rst), .b ({signal_1176, signal_1159}), .a ({Key_s1[4], Key_s0[4]}), .c ({signal_1178, signal_1095}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_774 ( .s (rst), .b ({signal_1179, signal_1158}), .a ({Key_s1[5], Key_s0[5]}), .c ({signal_1181, signal_1094}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_775 ( .s (rst), .b ({signal_1182, signal_1157}), .a ({Key_s1[6], Key_s0[6]}), .c ({signal_1184, signal_1093}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_776 ( .s (rst), .b ({signal_1185, signal_1156}), .a ({Key_s1[7], Key_s0[7]}), .c ({signal_1187, signal_1092}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_777 ( .s (rst), .b ({signal_1188, signal_1155}), .a ({Key_s1[8], Key_s0[8]}), .c ({signal_1190, signal_1091}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_778 ( .s (rst), .b ({signal_1191, signal_1154}), .a ({Key_s1[9], Key_s0[9]}), .c ({signal_1193, signal_1090}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_779 ( .s (rst), .b ({signal_1194, signal_1153}), .a ({Key_s1[10], Key_s0[10]}), .c ({signal_1196, signal_1089}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_780 ( .s (rst), .b ({signal_1197, signal_1152}), .a ({Key_s1[11], Key_s0[11]}), .c ({signal_1199, signal_1088}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_781 ( .s (rst), .b ({signal_1200, signal_1151}), .a ({Key_s1[12], Key_s0[12]}), .c ({signal_1202, signal_1087}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_782 ( .s (rst), .b ({signal_1203, signal_1150}), .a ({Key_s1[13], Key_s0[13]}), .c ({signal_1205, signal_1086}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_783 ( .s (rst), .b ({signal_1206, signal_1149}), .a ({Key_s1[14], Key_s0[14]}), .c ({signal_1208, signal_1085}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_784 ( .s (rst), .b ({signal_1209, signal_1148}), .a ({Key_s1[15], Key_s0[15]}), .c ({signal_1211, signal_1084}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_785 ( .s (rst), .b ({signal_1212, signal_1147}), .a ({Key_s1[16], Key_s0[16]}), .c ({signal_1214, signal_1083}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_786 ( .s (rst), .b ({signal_1215, signal_1146}), .a ({Key_s1[17], Key_s0[17]}), .c ({signal_1217, signal_1082}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_787 ( .s (rst), .b ({signal_1218, signal_1145}), .a ({Key_s1[18], Key_s0[18]}), .c ({signal_1220, signal_1081}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_788 ( .s (rst), .b ({signal_1221, signal_1144}), .a ({Key_s1[19], Key_s0[19]}), .c ({signal_1223, signal_1080}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_789 ( .s (rst), .b ({signal_1224, signal_1143}), .a ({Key_s1[20], Key_s0[20]}), .c ({signal_1226, signal_1079}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_790 ( .s (rst), .b ({signal_1227, signal_1142}), .a ({Key_s1[21], Key_s0[21]}), .c ({signal_1229, signal_1078}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_791 ( .s (rst), .b ({signal_1230, signal_1141}), .a ({Key_s1[22], Key_s0[22]}), .c ({signal_1232, signal_1077}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_792 ( .s (rst), .b ({signal_1233, signal_1140}), .a ({Key_s1[23], Key_s0[23]}), .c ({signal_1235, signal_1076}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_793 ( .s (rst), .b ({signal_1236, signal_1139}), .a ({Key_s1[24], Key_s0[24]}), .c ({signal_1238, signal_1075}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_794 ( .s (rst), .b ({signal_1239, signal_1138}), .a ({Key_s1[25], Key_s0[25]}), .c ({signal_1241, signal_1074}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_795 ( .s (rst), .b ({signal_1242, signal_1137}), .a ({Key_s1[26], Key_s0[26]}), .c ({signal_1244, signal_1073}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_796 ( .s (rst), .b ({signal_1245, signal_1136}), .a ({Key_s1[27], Key_s0[27]}), .c ({signal_1247, signal_1072}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_797 ( .s (rst), .b ({signal_1248, signal_1135}), .a ({Key_s1[28], Key_s0[28]}), .c ({signal_1250, signal_1071}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_798 ( .s (rst), .b ({signal_1251, signal_1134}), .a ({Key_s1[29], Key_s0[29]}), .c ({signal_1253, signal_1070}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_799 ( .s (rst), .b ({signal_1254, signal_1133}), .a ({Key_s1[30], Key_s0[30]}), .c ({signal_1256, signal_1069}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_800 ( .s (rst), .b ({signal_1257, signal_1132}), .a ({Key_s1[31], Key_s0[31]}), .c ({signal_1259, signal_1068}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_801 ( .s (rst), .b ({signal_1260, signal_1131}), .a ({Key_s1[32], Key_s0[32]}), .c ({signal_1262, signal_1067}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_802 ( .s (rst), .b ({signal_1263, signal_1130}), .a ({Key_s1[33], Key_s0[33]}), .c ({signal_1265, signal_1066}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_803 ( .s (rst), .b ({signal_1266, signal_1129}), .a ({Key_s1[34], Key_s0[34]}), .c ({signal_1268, signal_1065}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_804 ( .s (rst), .b ({signal_1269, signal_1128}), .a ({Key_s1[35], Key_s0[35]}), .c ({signal_1271, signal_1064}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_805 ( .s (rst), .b ({signal_1272, signal_1127}), .a ({Key_s1[36], Key_s0[36]}), .c ({signal_1274, signal_1063}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_806 ( .s (rst), .b ({signal_1275, signal_1126}), .a ({Key_s1[37], Key_s0[37]}), .c ({signal_1277, signal_1062}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_807 ( .s (rst), .b ({signal_1278, signal_1125}), .a ({Key_s1[38], Key_s0[38]}), .c ({signal_1280, signal_1061}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_808 ( .s (rst), .b ({signal_1281, signal_1124}), .a ({Key_s1[39], Key_s0[39]}), .c ({signal_1283, signal_1060}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_809 ( .s (rst), .b ({signal_1284, signal_1123}), .a ({Key_s1[40], Key_s0[40]}), .c ({signal_1286, signal_1059}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_810 ( .s (rst), .b ({signal_1287, signal_1122}), .a ({Key_s1[41], Key_s0[41]}), .c ({signal_1289, signal_1058}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_811 ( .s (rst), .b ({signal_1290, signal_1121}), .a ({Key_s1[42], Key_s0[42]}), .c ({signal_1292, signal_1057}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_812 ( .s (rst), .b ({signal_1293, signal_1120}), .a ({Key_s1[43], Key_s0[43]}), .c ({signal_1295, signal_1056}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_813 ( .s (rst), .b ({signal_1296, signal_1119}), .a ({Key_s1[44], Key_s0[44]}), .c ({signal_1298, signal_1055}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_814 ( .s (rst), .b ({signal_1299, signal_1118}), .a ({Key_s1[45], Key_s0[45]}), .c ({signal_1301, signal_1054}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_815 ( .s (rst), .b ({signal_1302, signal_1117}), .a ({Key_s1[46], Key_s0[46]}), .c ({signal_1304, signal_1053}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_816 ( .s (rst), .b ({signal_1305, signal_1116}), .a ({Key_s1[47], Key_s0[47]}), .c ({signal_1307, signal_1052}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_817 ( .s (rst), .b ({signal_1308, signal_1115}), .a ({Key_s1[48], Key_s0[48]}), .c ({signal_1310, signal_1051}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_818 ( .s (rst), .b ({signal_1311, signal_1114}), .a ({Key_s1[49], Key_s0[49]}), .c ({signal_1313, signal_1050}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_819 ( .s (rst), .b ({signal_1314, signal_1113}), .a ({Key_s1[50], Key_s0[50]}), .c ({signal_1316, signal_1049}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_820 ( .s (rst), .b ({signal_1317, signal_1112}), .a ({Key_s1[51], Key_s0[51]}), .c ({signal_1319, signal_1048}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_821 ( .s (rst), .b ({signal_1320, signal_1111}), .a ({Key_s1[52], Key_s0[52]}), .c ({signal_1322, signal_1047}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_822 ( .s (rst), .b ({signal_1323, signal_1110}), .a ({Key_s1[53], Key_s0[53]}), .c ({signal_1325, signal_1046}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_823 ( .s (rst), .b ({signal_1326, signal_1109}), .a ({Key_s1[54], Key_s0[54]}), .c ({signal_1328, signal_1045}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_824 ( .s (rst), .b ({signal_1329, signal_1108}), .a ({Key_s1[55], Key_s0[55]}), .c ({signal_1331, signal_1044}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_825 ( .s (rst), .b ({signal_1332, signal_1107}), .a ({Key_s1[56], Key_s0[56]}), .c ({signal_1334, signal_1043}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_826 ( .s (rst), .b ({signal_1335, signal_1106}), .a ({Key_s1[57], Key_s0[57]}), .c ({signal_1337, signal_1042}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_827 ( .s (rst), .b ({signal_1338, signal_1105}), .a ({Key_s1[58], Key_s0[58]}), .c ({signal_1340, signal_1041}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_828 ( .s (rst), .b ({signal_1341, signal_1104}), .a ({Key_s1[59], Key_s0[59]}), .c ({signal_1343, signal_1040}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_829 ( .s (rst), .b ({signal_1344, signal_1103}), .a ({Key_s1[60], Key_s0[60]}), .c ({signal_1346, signal_1039}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_830 ( .s (rst), .b ({signal_1347, signal_1102}), .a ({Key_s1[61], Key_s0[61]}), .c ({signal_1349, signal_1038}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_831 ( .s (rst), .b ({signal_1350, signal_1101}), .a ({Key_s1[62], Key_s0[62]}), .c ({signal_1352, signal_1037}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_832 ( .s (rst), .b ({signal_1353, signal_1100}), .a ({Key_s1[63], Key_s0[63]}), .c ({signal_1355, signal_1036}) ) ;
    MUX2_X1 cell_961 ( .S (rst), .A (signal_1029), .B (1'b1), .Z (signal_1035) ) ;
    MUX2_X1 cell_962 ( .S (rst), .A (signal_1028), .B (1'b0), .Z (signal_1034) ) ;
    MUX2_X1 cell_963 ( .S (rst), .A (signal_1027), .B (1'b0), .Z (signal_1033) ) ;
    MUX2_X1 cell_964 ( .S (rst), .A (signal_1026), .B (1'b0), .Z (signal_1032) ) ;
    MUX2_X1 cell_965 ( .S (rst), .A (signal_1025), .B (1'b0), .Z (signal_1031) ) ;
    MUX2_X1 cell_966 ( .S (rst), .A (signal_1024), .B (1'b0), .Z (signal_1030) ) ;
    MUX2_X1 cell_979 ( .S (signal_940), .A (signal_759), .B (signal_939), .Z (signal_1029) ) ;
    NAND2_X1 cell_980 ( .A1 (signal_939), .A2 (signal_760), .ZN (signal_759) ) ;
    NAND2_X1 cell_981 ( .A1 (signal_761), .A2 (signal_762), .ZN (signal_760) ) ;
    NOR2_X1 cell_982 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_762) ) ;
    AND2_X1 cell_983 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_761) ) ;
    AND2_X1 cell_984 ( .A1 (signal_763), .A2 (signal_943), .ZN (signal_1027) ) ;
    NAND2_X1 cell_985 ( .A1 (signal_764), .A2 (signal_939), .ZN (signal_763) ) ;
    NOR2_X1 cell_986 ( .A1 (signal_940), .A2 (signal_765), .ZN (signal_764) ) ;
    NAND2_X1 cell_987 ( .A1 (signal_1028), .A2 (signal_766), .ZN (signal_765) ) ;
    NOR2_X1 cell_988 ( .A1 (signal_1026), .A2 (signal_1025), .ZN (signal_766) ) ;
    OR2_X1 cell_989 ( .A1 (signal_940), .A2 (signal_767), .ZN (signal_1024) ) ;
    NOR2_X1 cell_990 ( .A1 (signal_1025), .A2 (signal_768), .ZN (signal_767) ) ;
    NAND2_X1 cell_991 ( .A1 (signal_939), .A2 (signal_769), .ZN (signal_768) ) ;
    NOR2_X1 cell_992 ( .A1 (signal_1026), .A2 (signal_770), .ZN (signal_769) ) ;
    NAND2_X1 cell_993 ( .A1 (signal_1028), .A2 (signal_943), .ZN (signal_770) ) ;
    NOR2_X1 cell_994 ( .A1 (signal_771), .A2 (signal_772), .ZN (done) ) ;
    NAND2_X1 cell_995 ( .A1 (signal_940), .A2 (signal_939), .ZN (signal_772) ) ;
    NAND2_X1 cell_996 ( .A1 (signal_773), .A2 (signal_774), .ZN (signal_771) ) ;
    NOR2_X1 cell_997 ( .A1 (signal_1025), .A2 (signal_775), .ZN (signal_774) ) ;
    INV_X1 cell_998 ( .A (signal_1028), .ZN (signal_775) ) ;
    NOR2_X1 cell_999 ( .A1 (signal_943), .A2 (signal_1026), .ZN (signal_773) ) ;
    ClockGatingController #(3) cell_1001 ( .clk (clk), .rst (rst), .GatedClk (signal_1676), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_0 ( .s (rst), .b ({signal_1483, signal_839}), .a ({Plaintext_s1[0], Plaintext_s0[0]}), .c ({signal_1485, signal_903}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_1 ( .s (rst), .b ({signal_1482, signal_838}), .a ({Plaintext_s1[1], Plaintext_s0[1]}), .c ({signal_1487, signal_902}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_2 ( .s (rst), .b ({signal_1481, signal_837}), .a ({Plaintext_s1[2], Plaintext_s0[2]}), .c ({signal_1489, signal_901}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_3 ( .s (rst), .b ({signal_1480, signal_836}), .a ({Plaintext_s1[3], Plaintext_s0[3]}), .c ({signal_1491, signal_900}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_4 ( .s (rst), .b ({signal_1479, signal_835}), .a ({Plaintext_s1[4], Plaintext_s0[4]}), .c ({signal_1493, signal_899}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_5 ( .s (rst), .b ({signal_1478, signal_834}), .a ({Plaintext_s1[5], Plaintext_s0[5]}), .c ({signal_1495, signal_898}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_6 ( .s (rst), .b ({signal_1477, signal_833}), .a ({Plaintext_s1[6], Plaintext_s0[6]}), .c ({signal_1497, signal_897}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_7 ( .s (rst), .b ({signal_1476, signal_832}), .a ({Plaintext_s1[7], Plaintext_s0[7]}), .c ({signal_1499, signal_896}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_8 ( .s (rst), .b ({signal_1475, signal_831}), .a ({Plaintext_s1[8], Plaintext_s0[8]}), .c ({signal_1501, signal_895}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_9 ( .s (rst), .b ({signal_1474, signal_830}), .a ({Plaintext_s1[9], Plaintext_s0[9]}), .c ({signal_1503, signal_894}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_10 ( .s (rst), .b ({signal_1473, signal_829}), .a ({Plaintext_s1[10], Plaintext_s0[10]}), .c ({signal_1505, signal_893}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_11 ( .s (rst), .b ({signal_1472, signal_828}), .a ({Plaintext_s1[11], Plaintext_s0[11]}), .c ({signal_1507, signal_892}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_12 ( .s (rst), .b ({signal_1471, signal_827}), .a ({Plaintext_s1[12], Plaintext_s0[12]}), .c ({signal_1509, signal_891}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_13 ( .s (rst), .b ({signal_1470, signal_826}), .a ({Plaintext_s1[13], Plaintext_s0[13]}), .c ({signal_1511, signal_890}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_14 ( .s (rst), .b ({signal_1469, signal_825}), .a ({Plaintext_s1[14], Plaintext_s0[14]}), .c ({signal_1513, signal_889}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_15 ( .s (rst), .b ({signal_1468, signal_824}), .a ({Plaintext_s1[15], Plaintext_s0[15]}), .c ({signal_1515, signal_888}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_16 ( .s (rst), .b ({signal_1467, signal_823}), .a ({Plaintext_s1[16], Plaintext_s0[16]}), .c ({signal_1517, signal_887}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_17 ( .s (rst), .b ({signal_1466, signal_822}), .a ({Plaintext_s1[17], Plaintext_s0[17]}), .c ({signal_1519, signal_886}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_18 ( .s (rst), .b ({signal_1465, signal_821}), .a ({Plaintext_s1[18], Plaintext_s0[18]}), .c ({signal_1521, signal_885}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_19 ( .s (rst), .b ({signal_1464, signal_820}), .a ({Plaintext_s1[19], Plaintext_s0[19]}), .c ({signal_1523, signal_884}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_20 ( .s (rst), .b ({signal_1463, signal_819}), .a ({Plaintext_s1[20], Plaintext_s0[20]}), .c ({signal_1525, signal_883}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_21 ( .s (rst), .b ({signal_1462, signal_818}), .a ({Plaintext_s1[21], Plaintext_s0[21]}), .c ({signal_1527, signal_882}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_22 ( .s (rst), .b ({signal_1461, signal_817}), .a ({Plaintext_s1[22], Plaintext_s0[22]}), .c ({signal_1529, signal_881}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_23 ( .s (rst), .b ({signal_1460, signal_816}), .a ({Plaintext_s1[23], Plaintext_s0[23]}), .c ({signal_1531, signal_880}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_24 ( .s (rst), .b ({signal_1459, signal_815}), .a ({Plaintext_s1[24], Plaintext_s0[24]}), .c ({signal_1533, signal_879}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_25 ( .s (rst), .b ({signal_1458, signal_814}), .a ({Plaintext_s1[25], Plaintext_s0[25]}), .c ({signal_1535, signal_878}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_26 ( .s (rst), .b ({signal_1457, signal_813}), .a ({Plaintext_s1[26], Plaintext_s0[26]}), .c ({signal_1537, signal_877}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_27 ( .s (rst), .b ({signal_1456, signal_812}), .a ({Plaintext_s1[27], Plaintext_s0[27]}), .c ({signal_1539, signal_876}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_28 ( .s (rst), .b ({signal_1455, signal_811}), .a ({Plaintext_s1[28], Plaintext_s0[28]}), .c ({signal_1541, signal_875}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_29 ( .s (rst), .b ({signal_1454, signal_810}), .a ({Plaintext_s1[29], Plaintext_s0[29]}), .c ({signal_1543, signal_874}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_30 ( .s (rst), .b ({signal_1453, signal_809}), .a ({Plaintext_s1[30], Plaintext_s0[30]}), .c ({signal_1545, signal_873}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_31 ( .s (rst), .b ({signal_1452, signal_808}), .a ({Plaintext_s1[31], Plaintext_s0[31]}), .c ({signal_1547, signal_872}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_32 ( .s (rst), .b ({signal_1451, signal_807}), .a ({Plaintext_s1[32], Plaintext_s0[32]}), .c ({signal_1549, signal_871}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_33 ( .s (rst), .b ({signal_1450, signal_806}), .a ({Plaintext_s1[33], Plaintext_s0[33]}), .c ({signal_1551, signal_870}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_34 ( .s (rst), .b ({signal_1449, signal_805}), .a ({Plaintext_s1[34], Plaintext_s0[34]}), .c ({signal_1553, signal_869}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_35 ( .s (rst), .b ({signal_1448, signal_804}), .a ({Plaintext_s1[35], Plaintext_s0[35]}), .c ({signal_1555, signal_868}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_36 ( .s (rst), .b ({signal_1447, signal_803}), .a ({Plaintext_s1[36], Plaintext_s0[36]}), .c ({signal_1557, signal_867}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_37 ( .s (rst), .b ({signal_1446, signal_802}), .a ({Plaintext_s1[37], Plaintext_s0[37]}), .c ({signal_1559, signal_866}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_38 ( .s (rst), .b ({signal_1445, signal_801}), .a ({Plaintext_s1[38], Plaintext_s0[38]}), .c ({signal_1561, signal_865}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_39 ( .s (rst), .b ({signal_1444, signal_800}), .a ({Plaintext_s1[39], Plaintext_s0[39]}), .c ({signal_1563, signal_864}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_40 ( .s (rst), .b ({signal_1443, signal_799}), .a ({Plaintext_s1[40], Plaintext_s0[40]}), .c ({signal_1565, signal_863}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_41 ( .s (rst), .b ({signal_1442, signal_798}), .a ({Plaintext_s1[41], Plaintext_s0[41]}), .c ({signal_1567, signal_862}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_42 ( .s (rst), .b ({signal_1441, signal_797}), .a ({Plaintext_s1[42], Plaintext_s0[42]}), .c ({signal_1569, signal_861}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_43 ( .s (rst), .b ({signal_1440, signal_796}), .a ({Plaintext_s1[43], Plaintext_s0[43]}), .c ({signal_1571, signal_860}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_44 ( .s (rst), .b ({signal_1439, signal_795}), .a ({Plaintext_s1[44], Plaintext_s0[44]}), .c ({signal_1573, signal_859}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_45 ( .s (rst), .b ({signal_1438, signal_794}), .a ({Plaintext_s1[45], Plaintext_s0[45]}), .c ({signal_1575, signal_858}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_46 ( .s (rst), .b ({signal_1437, signal_793}), .a ({Plaintext_s1[46], Plaintext_s0[46]}), .c ({signal_1577, signal_857}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_47 ( .s (rst), .b ({signal_1436, signal_792}), .a ({Plaintext_s1[47], Plaintext_s0[47]}), .c ({signal_1579, signal_856}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_48 ( .s (rst), .b ({signal_1435, signal_791}), .a ({Plaintext_s1[48], Plaintext_s0[48]}), .c ({signal_1581, signal_855}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_49 ( .s (rst), .b ({signal_1434, signal_790}), .a ({Plaintext_s1[49], Plaintext_s0[49]}), .c ({signal_1583, signal_854}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_50 ( .s (rst), .b ({signal_1433, signal_789}), .a ({Plaintext_s1[50], Plaintext_s0[50]}), .c ({signal_1585, signal_853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_51 ( .s (rst), .b ({signal_1432, signal_788}), .a ({Plaintext_s1[51], Plaintext_s0[51]}), .c ({signal_1587, signal_852}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_52 ( .s (rst), .b ({signal_1431, signal_787}), .a ({Plaintext_s1[52], Plaintext_s0[52]}), .c ({signal_1589, signal_851}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_53 ( .s (rst), .b ({signal_1430, signal_786}), .a ({Plaintext_s1[53], Plaintext_s0[53]}), .c ({signal_1591, signal_850}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_54 ( .s (rst), .b ({signal_1429, signal_785}), .a ({Plaintext_s1[54], Plaintext_s0[54]}), .c ({signal_1593, signal_849}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_55 ( .s (rst), .b ({signal_1428, signal_784}), .a ({Plaintext_s1[55], Plaintext_s0[55]}), .c ({signal_1595, signal_848}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_56 ( .s (rst), .b ({signal_1427, signal_783}), .a ({Plaintext_s1[56], Plaintext_s0[56]}), .c ({signal_1597, signal_847}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_57 ( .s (rst), .b ({signal_1426, signal_782}), .a ({Plaintext_s1[57], Plaintext_s0[57]}), .c ({signal_1599, signal_846}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_58 ( .s (rst), .b ({signal_1425, signal_781}), .a ({Plaintext_s1[58], Plaintext_s0[58]}), .c ({signal_1601, signal_845}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_59 ( .s (rst), .b ({signal_1424, signal_780}), .a ({Plaintext_s1[59], Plaintext_s0[59]}), .c ({signal_1603, signal_844}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_60 ( .s (rst), .b ({signal_1423, signal_779}), .a ({Plaintext_s1[60], Plaintext_s0[60]}), .c ({signal_1605, signal_843}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_61 ( .s (rst), .b ({signal_1422, signal_778}), .a ({Plaintext_s1[61], Plaintext_s0[61]}), .c ({signal_1607, signal_842}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_62 ( .s (rst), .b ({signal_1421, signal_777}), .a ({Plaintext_s1[62], Plaintext_s0[62]}), .c ({signal_1609, signal_841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) cell_63 ( .s (rst), .b ({signal_1420, signal_776}), .a ({Plaintext_s1[63], Plaintext_s0[63]}), .c ({signal_1611, signal_840}) ) ;
    SkinnyTop_step2_ANF #(.low_latency(0), .pipeline(0)) cell_1000 ( .in0 ({signal_943, signal_940, signal_939, Ciphertext_s0[0], Ciphertext_s0[1], Ciphertext_s0[2], Ciphertext_s0[3], Ciphertext_s0[4], Ciphertext_s0[5], Ciphertext_s0[6], Ciphertext_s0[7], Ciphertext_s0[8], Ciphertext_s0[9], Ciphertext_s0[10], Ciphertext_s0[11], Ciphertext_s0[12], Ciphertext_s0[13], Ciphertext_s0[14], Ciphertext_s0[15], Ciphertext_s0[16], Ciphertext_s0[17], Ciphertext_s0[18], Ciphertext_s0[19], Ciphertext_s0[20], Ciphertext_s0[21], Ciphertext_s0[22], Ciphertext_s0[23], Ciphertext_s0[24], Ciphertext_s0[25], Ciphertext_s0[26], Ciphertext_s0[27], Ciphertext_s0[28], Ciphertext_s0[29], Ciphertext_s0[30], Ciphertext_s0[31], Ciphertext_s0[32], Ciphertext_s0[33], Ciphertext_s0[34], Ciphertext_s0[35], Ciphertext_s0[36], Ciphertext_s0[37], Ciphertext_s0[38], Ciphertext_s0[39], Ciphertext_s0[40], Ciphertext_s0[41], Ciphertext_s0[42], Ciphertext_s0[43], Ciphertext_s0[44], Ciphertext_s0[45], Ciphertext_s0[46], Ciphertext_s0[47], Ciphertext_s0[48], Ciphertext_s0[49], Ciphertext_s0[50], Ciphertext_s0[51], Ciphertext_s0[52], Ciphertext_s0[53], Ciphertext_s0[54], Ciphertext_s0[55], Ciphertext_s0[56], Ciphertext_s0[57], Ciphertext_s0[58], Ciphertext_s0[59], Ciphertext_s0[60], Ciphertext_s0[61], Ciphertext_s0[62], Ciphertext_s0[63], signal_1163, signal_1162, signal_1161, signal_1160, signal_1159, signal_1158, signal_1157, signal_1156, signal_1155, signal_1154, signal_1153, signal_1152, signal_1151, signal_1150, signal_1149, signal_1148, signal_1147, signal_1146, signal_1145, signal_1144, signal_1143, signal_1142, signal_1141, signal_1140, signal_1139, signal_1138, signal_1137, signal_1136, signal_1135, signal_1134, signal_1133, signal_1132, signal_1028, signal_1026, signal_1025, 1'b0}), .in1 ({1'b0, 1'b0, 1'b0, Ciphertext_s1[0], Ciphertext_s1[1], Ciphertext_s1[2], Ciphertext_s1[3], Ciphertext_s1[4], Ciphertext_s1[5], Ciphertext_s1[6], Ciphertext_s1[7], Ciphertext_s1[8], Ciphertext_s1[9], Ciphertext_s1[10], Ciphertext_s1[11], Ciphertext_s1[12], Ciphertext_s1[13], Ciphertext_s1[14], Ciphertext_s1[15], Ciphertext_s1[16], Ciphertext_s1[17], Ciphertext_s1[18], Ciphertext_s1[19], Ciphertext_s1[20], Ciphertext_s1[21], Ciphertext_s1[22], Ciphertext_s1[23], Ciphertext_s1[24], Ciphertext_s1[25], Ciphertext_s1[26], Ciphertext_s1[27], Ciphertext_s1[28], Ciphertext_s1[29], Ciphertext_s1[30], Ciphertext_s1[31], Ciphertext_s1[32], Ciphertext_s1[33], Ciphertext_s1[34], Ciphertext_s1[35], Ciphertext_s1[36], Ciphertext_s1[37], Ciphertext_s1[38], Ciphertext_s1[39], Ciphertext_s1[40], Ciphertext_s1[41], Ciphertext_s1[42], Ciphertext_s1[43], Ciphertext_s1[44], Ciphertext_s1[45], Ciphertext_s1[46], Ciphertext_s1[47], Ciphertext_s1[48], Ciphertext_s1[49], Ciphertext_s1[50], Ciphertext_s1[51], Ciphertext_s1[52], Ciphertext_s1[53], Ciphertext_s1[54], Ciphertext_s1[55], Ciphertext_s1[56], Ciphertext_s1[57], Ciphertext_s1[58], Ciphertext_s1[59], Ciphertext_s1[60], Ciphertext_s1[61], Ciphertext_s1[62], Ciphertext_s1[63], signal_1164, signal_1167, signal_1170, signal_1173, signal_1176, signal_1179, signal_1182, signal_1185, signal_1188, signal_1191, signal_1194, signal_1197, signal_1200, signal_1203, signal_1206, signal_1209, signal_1212, signal_1215, signal_1218, signal_1221, signal_1224, signal_1227, signal_1230, signal_1233, signal_1236, signal_1239, signal_1242, signal_1245, signal_1248, signal_1251, signal_1254, signal_1257, 1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_839, signal_838, signal_837, signal_836, signal_835, signal_834, signal_833, signal_832, signal_831, signal_830, signal_829, signal_828, signal_827, signal_826, signal_825, signal_824, signal_823, signal_822, signal_821, signal_820, signal_819, signal_818, signal_817, signal_816, signal_815, signal_814, signal_813, signal_812, signal_811, signal_810, signal_809, signal_808, signal_807, signal_806, signal_805, signal_804, signal_803, signal_802, signal_801, signal_800, signal_799, signal_798, signal_797, signal_796, signal_795, signal_794, signal_793, signal_792, signal_791, signal_790, signal_789, signal_788, signal_787, signal_786, signal_785, signal_784, signal_783, signal_782, signal_781, signal_780, signal_779, signal_778, signal_777, signal_776}), .out1 ({signal_1483, signal_1482, signal_1481, signal_1480, signal_1479, signal_1478, signal_1477, signal_1476, signal_1475, signal_1474, signal_1473, signal_1472, signal_1471, signal_1470, signal_1469, signal_1468, signal_1467, signal_1466, signal_1465, signal_1464, signal_1463, signal_1462, signal_1461, signal_1460, signal_1459, signal_1458, signal_1457, signal_1456, signal_1455, signal_1454, signal_1453, signal_1452, signal_1451, signal_1450, signal_1449, signal_1448, signal_1447, signal_1446, signal_1445, signal_1444, signal_1443, signal_1442, signal_1441, signal_1440, signal_1439, signal_1438, signal_1437, signal_1436, signal_1435, signal_1434, signal_1433, signal_1432, signal_1431, signal_1430, signal_1429, signal_1428, signal_1427, signal_1426, signal_1425, signal_1424, signal_1423, signal_1422, signal_1421, signal_1420}) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(0)) cell_65 ( .clk (signal_1676), .D ({signal_1611, signal_840}), .Q ({Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_67 ( .clk (signal_1676), .D ({signal_1609, signal_841}), .Q ({Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_69 ( .clk (signal_1676), .D ({signal_1607, signal_842}), .Q ({Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_71 ( .clk (signal_1676), .D ({signal_1605, signal_843}), .Q ({Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_73 ( .clk (signal_1676), .D ({signal_1603, signal_844}), .Q ({Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_75 ( .clk (signal_1676), .D ({signal_1601, signal_845}), .Q ({Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_77 ( .clk (signal_1676), .D ({signal_1599, signal_846}), .Q ({Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_79 ( .clk (signal_1676), .D ({signal_1597, signal_847}), .Q ({Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_81 ( .clk (signal_1676), .D ({signal_1595, signal_848}), .Q ({Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_83 ( .clk (signal_1676), .D ({signal_1593, signal_849}), .Q ({Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_85 ( .clk (signal_1676), .D ({signal_1591, signal_850}), .Q ({Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_87 ( .clk (signal_1676), .D ({signal_1589, signal_851}), .Q ({Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_89 ( .clk (signal_1676), .D ({signal_1587, signal_852}), .Q ({Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_91 ( .clk (signal_1676), .D ({signal_1585, signal_853}), .Q ({Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_93 ( .clk (signal_1676), .D ({signal_1583, signal_854}), .Q ({Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_95 ( .clk (signal_1676), .D ({signal_1581, signal_855}), .Q ({Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_97 ( .clk (signal_1676), .D ({signal_1579, signal_856}), .Q ({Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_99 ( .clk (signal_1676), .D ({signal_1577, signal_857}), .Q ({Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_101 ( .clk (signal_1676), .D ({signal_1575, signal_858}), .Q ({Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_103 ( .clk (signal_1676), .D ({signal_1573, signal_859}), .Q ({Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_105 ( .clk (signal_1676), .D ({signal_1571, signal_860}), .Q ({Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_107 ( .clk (signal_1676), .D ({signal_1569, signal_861}), .Q ({Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_109 ( .clk (signal_1676), .D ({signal_1567, signal_862}), .Q ({Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_111 ( .clk (signal_1676), .D ({signal_1565, signal_863}), .Q ({Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_113 ( .clk (signal_1676), .D ({signal_1563, signal_864}), .Q ({Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_115 ( .clk (signal_1676), .D ({signal_1561, signal_865}), .Q ({Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_117 ( .clk (signal_1676), .D ({signal_1559, signal_866}), .Q ({Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_119 ( .clk (signal_1676), .D ({signal_1557, signal_867}), .Q ({Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_121 ( .clk (signal_1676), .D ({signal_1555, signal_868}), .Q ({Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_123 ( .clk (signal_1676), .D ({signal_1553, signal_869}), .Q ({Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_125 ( .clk (signal_1676), .D ({signal_1551, signal_870}), .Q ({Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_127 ( .clk (signal_1676), .D ({signal_1549, signal_871}), .Q ({Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_129 ( .clk (signal_1676), .D ({signal_1547, signal_872}), .Q ({Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_131 ( .clk (signal_1676), .D ({signal_1545, signal_873}), .Q ({Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_133 ( .clk (signal_1676), .D ({signal_1543, signal_874}), .Q ({Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_135 ( .clk (signal_1676), .D ({signal_1541, signal_875}), .Q ({Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_137 ( .clk (signal_1676), .D ({signal_1539, signal_876}), .Q ({Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_139 ( .clk (signal_1676), .D ({signal_1537, signal_877}), .Q ({Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_141 ( .clk (signal_1676), .D ({signal_1535, signal_878}), .Q ({Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_143 ( .clk (signal_1676), .D ({signal_1533, signal_879}), .Q ({Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_145 ( .clk (signal_1676), .D ({signal_1531, signal_880}), .Q ({Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_147 ( .clk (signal_1676), .D ({signal_1529, signal_881}), .Q ({Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_149 ( .clk (signal_1676), .D ({signal_1527, signal_882}), .Q ({Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_151 ( .clk (signal_1676), .D ({signal_1525, signal_883}), .Q ({Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_153 ( .clk (signal_1676), .D ({signal_1523, signal_884}), .Q ({Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_155 ( .clk (signal_1676), .D ({signal_1521, signal_885}), .Q ({Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_157 ( .clk (signal_1676), .D ({signal_1519, signal_886}), .Q ({Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_159 ( .clk (signal_1676), .D ({signal_1517, signal_887}), .Q ({Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_161 ( .clk (signal_1676), .D ({signal_1515, signal_888}), .Q ({Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_163 ( .clk (signal_1676), .D ({signal_1513, signal_889}), .Q ({Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_165 ( .clk (signal_1676), .D ({signal_1511, signal_890}), .Q ({Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_167 ( .clk (signal_1676), .D ({signal_1509, signal_891}), .Q ({Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_169 ( .clk (signal_1676), .D ({signal_1507, signal_892}), .Q ({Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_171 ( .clk (signal_1676), .D ({signal_1505, signal_893}), .Q ({Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_173 ( .clk (signal_1676), .D ({signal_1503, signal_894}), .Q ({Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_175 ( .clk (signal_1676), .D ({signal_1501, signal_895}), .Q ({Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_177 ( .clk (signal_1676), .D ({signal_1499, signal_896}), .Q ({Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_179 ( .clk (signal_1676), .D ({signal_1497, signal_897}), .Q ({Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_181 ( .clk (signal_1676), .D ({signal_1495, signal_898}), .Q ({Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_183 ( .clk (signal_1676), .D ({signal_1493, signal_899}), .Q ({Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_185 ( .clk (signal_1676), .D ({signal_1491, signal_900}), .Q ({Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_187 ( .clk (signal_1676), .D ({signal_1489, signal_901}), .Q ({Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_189 ( .clk (signal_1676), .D ({signal_1487, signal_902}), .Q ({Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_191 ( .clk (signal_1676), .D ({signal_1485, signal_903}), .Q ({Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_834 ( .clk (signal_1676), .D ({signal_1355, signal_1036}), .Q ({signal_1257, signal_1132}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_836 ( .clk (signal_1676), .D ({signal_1352, signal_1037}), .Q ({signal_1254, signal_1133}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_838 ( .clk (signal_1676), .D ({signal_1349, signal_1038}), .Q ({signal_1251, signal_1134}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_840 ( .clk (signal_1676), .D ({signal_1346, signal_1039}), .Q ({signal_1248, signal_1135}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_842 ( .clk (signal_1676), .D ({signal_1343, signal_1040}), .Q ({signal_1245, signal_1136}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_844 ( .clk (signal_1676), .D ({signal_1340, signal_1041}), .Q ({signal_1242, signal_1137}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_846 ( .clk (signal_1676), .D ({signal_1337, signal_1042}), .Q ({signal_1239, signal_1138}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_848 ( .clk (signal_1676), .D ({signal_1334, signal_1043}), .Q ({signal_1236, signal_1139}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_850 ( .clk (signal_1676), .D ({signal_1331, signal_1044}), .Q ({signal_1233, signal_1140}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_852 ( .clk (signal_1676), .D ({signal_1328, signal_1045}), .Q ({signal_1230, signal_1141}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_854 ( .clk (signal_1676), .D ({signal_1325, signal_1046}), .Q ({signal_1227, signal_1142}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_856 ( .clk (signal_1676), .D ({signal_1322, signal_1047}), .Q ({signal_1224, signal_1143}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_858 ( .clk (signal_1676), .D ({signal_1319, signal_1048}), .Q ({signal_1221, signal_1144}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_860 ( .clk (signal_1676), .D ({signal_1316, signal_1049}), .Q ({signal_1218, signal_1145}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_862 ( .clk (signal_1676), .D ({signal_1313, signal_1050}), .Q ({signal_1215, signal_1146}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_864 ( .clk (signal_1676), .D ({signal_1310, signal_1051}), .Q ({signal_1212, signal_1147}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_866 ( .clk (signal_1676), .D ({signal_1307, signal_1052}), .Q ({signal_1209, signal_1148}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_868 ( .clk (signal_1676), .D ({signal_1304, signal_1053}), .Q ({signal_1206, signal_1149}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_870 ( .clk (signal_1676), .D ({signal_1301, signal_1054}), .Q ({signal_1203, signal_1150}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_872 ( .clk (signal_1676), .D ({signal_1298, signal_1055}), .Q ({signal_1200, signal_1151}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_874 ( .clk (signal_1676), .D ({signal_1295, signal_1056}), .Q ({signal_1197, signal_1152}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_876 ( .clk (signal_1676), .D ({signal_1292, signal_1057}), .Q ({signal_1194, signal_1153}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_878 ( .clk (signal_1676), .D ({signal_1289, signal_1058}), .Q ({signal_1191, signal_1154}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_880 ( .clk (signal_1676), .D ({signal_1286, signal_1059}), .Q ({signal_1188, signal_1155}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_882 ( .clk (signal_1676), .D ({signal_1283, signal_1060}), .Q ({signal_1185, signal_1156}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_884 ( .clk (signal_1676), .D ({signal_1280, signal_1061}), .Q ({signal_1182, signal_1157}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_886 ( .clk (signal_1676), .D ({signal_1277, signal_1062}), .Q ({signal_1179, signal_1158}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_888 ( .clk (signal_1676), .D ({signal_1274, signal_1063}), .Q ({signal_1176, signal_1159}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_890 ( .clk (signal_1676), .D ({signal_1271, signal_1064}), .Q ({signal_1173, signal_1160}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_892 ( .clk (signal_1676), .D ({signal_1268, signal_1065}), .Q ({signal_1170, signal_1161}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_894 ( .clk (signal_1676), .D ({signal_1265, signal_1066}), .Q ({signal_1167, signal_1162}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_896 ( .clk (signal_1676), .D ({signal_1262, signal_1067}), .Q ({signal_1164, signal_1163}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_898 ( .clk (signal_1676), .D ({signal_1259, signal_1068}), .Q ({signal_1329, signal_1108}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_900 ( .clk (signal_1676), .D ({signal_1256, signal_1069}), .Q ({signal_1326, signal_1109}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_902 ( .clk (signal_1676), .D ({signal_1253, signal_1070}), .Q ({signal_1323, signal_1110}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_904 ( .clk (signal_1676), .D ({signal_1250, signal_1071}), .Q ({signal_1320, signal_1111}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_906 ( .clk (signal_1676), .D ({signal_1247, signal_1072}), .Q ({signal_1353, signal_1100}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_908 ( .clk (signal_1676), .D ({signal_1244, signal_1073}), .Q ({signal_1350, signal_1101}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_910 ( .clk (signal_1676), .D ({signal_1241, signal_1074}), .Q ({signal_1347, signal_1102}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_912 ( .clk (signal_1676), .D ({signal_1238, signal_1075}), .Q ({signal_1344, signal_1103}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_914 ( .clk (signal_1676), .D ({signal_1235, signal_1076}), .Q ({signal_1305, signal_1116}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_916 ( .clk (signal_1676), .D ({signal_1232, signal_1077}), .Q ({signal_1302, signal_1117}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_918 ( .clk (signal_1676), .D ({signal_1229, signal_1078}), .Q ({signal_1299, signal_1118}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_920 ( .clk (signal_1676), .D ({signal_1226, signal_1079}), .Q ({signal_1296, signal_1119}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_922 ( .clk (signal_1676), .D ({signal_1223, signal_1080}), .Q ({signal_1269, signal_1128}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_924 ( .clk (signal_1676), .D ({signal_1220, signal_1081}), .Q ({signal_1266, signal_1129}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_926 ( .clk (signal_1676), .D ({signal_1217, signal_1082}), .Q ({signal_1263, signal_1130}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_928 ( .clk (signal_1676), .D ({signal_1214, signal_1083}), .Q ({signal_1260, signal_1131}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_930 ( .clk (signal_1676), .D ({signal_1211, signal_1084}), .Q ({signal_1281, signal_1124}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_932 ( .clk (signal_1676), .D ({signal_1208, signal_1085}), .Q ({signal_1278, signal_1125}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_934 ( .clk (signal_1676), .D ({signal_1205, signal_1086}), .Q ({signal_1275, signal_1126}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_936 ( .clk (signal_1676), .D ({signal_1202, signal_1087}), .Q ({signal_1272, signal_1127}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_938 ( .clk (signal_1676), .D ({signal_1199, signal_1088}), .Q ({signal_1317, signal_1112}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_940 ( .clk (signal_1676), .D ({signal_1196, signal_1089}), .Q ({signal_1314, signal_1113}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_942 ( .clk (signal_1676), .D ({signal_1193, signal_1090}), .Q ({signal_1311, signal_1114}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_944 ( .clk (signal_1676), .D ({signal_1190, signal_1091}), .Q ({signal_1308, signal_1115}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_946 ( .clk (signal_1676), .D ({signal_1187, signal_1092}), .Q ({signal_1293, signal_1120}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_948 ( .clk (signal_1676), .D ({signal_1184, signal_1093}), .Q ({signal_1290, signal_1121}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_950 ( .clk (signal_1676), .D ({signal_1181, signal_1094}), .Q ({signal_1287, signal_1122}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_952 ( .clk (signal_1676), .D ({signal_1178, signal_1095}), .Q ({signal_1284, signal_1123}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_954 ( .clk (signal_1676), .D ({signal_1175, signal_1096}), .Q ({signal_1341, signal_1104}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_956 ( .clk (signal_1676), .D ({signal_1172, signal_1097}), .Q ({signal_1338, signal_1105}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_958 ( .clk (signal_1676), .D ({signal_1169, signal_1098}), .Q ({signal_1335, signal_1106}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) cell_960 ( .clk (signal_1676), .D ({signal_1166, signal_1099}), .Q ({signal_1332, signal_1107}) ) ;
    DFF_X1 cell_968 ( .CK (signal_1676), .D (signal_1030), .Q (signal_939), .QN () ) ;
    DFF_X1 cell_970 ( .CK (signal_1676), .D (signal_1031), .Q (signal_940), .QN () ) ;
    DFF_X1 cell_972 ( .CK (signal_1676), .D (signal_1032), .Q (signal_1025), .QN () ) ;
    DFF_X1 cell_974 ( .CK (signal_1676), .D (signal_1033), .Q (signal_1026), .QN () ) ;
    DFF_X1 cell_976 ( .CK (signal_1676), .D (signal_1034), .Q (signal_943), .QN () ) ;
    DFF_X1 cell_978 ( .CK (signal_1676), .D (signal_1035), .Q (signal_1028), .QN () ) ;
endmodule
