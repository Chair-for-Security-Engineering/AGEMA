module Reg1(x, y);
 input [74:0] x;
 output [73:0] y;

  register_stage #(.WIDTH(74)) inst_0(.clk(x[71]), .D({x[72],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[73],x[74],x[0],x[11],x[22],x[33],x[44],x[55],x[60],x[61],x[62],x[63],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[56],x[57],x[58],x[59]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73]}));
endmodule

module Reg2(x, y);
 input [182:0] x;
 output [181:0] y;

  register_stage #(.WIDTH(182)) inst_0(.clk(x[161]), .D({x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx5(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx6(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx12(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx13(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx19(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx20(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx26(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx27(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx33(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx34(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx40(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx41(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx47(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx48(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx54(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx55(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx61(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx62(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx68(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx69(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx70(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx71(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx72(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx73(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx74(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx75(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx76(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx77(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx78(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx79(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx80(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx81(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx82(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx83(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx84(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx85(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx86(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx87(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx88(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx89(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx90(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx91(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx92(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx93(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx94(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx95(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx96(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx97(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx98(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx99(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx100(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx101(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx102(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx103(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx104(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx105(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx106(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx107(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx108(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx109(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx110(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx111(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx112(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx113(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx114(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx115(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx116(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx117(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx118(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx119(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx120(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx121(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx122(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx123(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx124(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx125(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx126(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx127(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx128(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx129(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx130(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx131(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx132(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx133(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx134(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx135(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx136(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx137(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx138(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx139(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx140(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx141(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx142(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx143(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx144(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx145(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx146(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx147(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx148(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx149(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx150(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx151(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx152(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx153(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx154(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx155(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx156(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx157(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx158(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx159(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx160(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx161(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx162(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx163(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx164(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx165(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx166(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx167(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx168(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx169(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx170(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx171(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx172(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx173(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx174(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx175(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx176(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx177(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx178(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx179(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx180(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx181(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module FX(x, y);
 input [255:0] x;
 output [181:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[3], x[0]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[4], x[0]}), .y(y[3]));
  Fx4 Fx4_inst(.x(x[5]), .y(y[4]));
  Fx5 Fx5_inst(.x(x[6]), .y(y[5]));
  Fx6 Fx6_inst(.x(x[7]), .y(y[6]));
  Fx7 Fx7_inst(.x({x[9], x[8]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[10], x[8]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[11], x[8]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[12], x[8]}), .y(y[10]));
  Fx11 Fx11_inst(.x(x[13]), .y(y[11]));
  Fx12 Fx12_inst(.x(x[14]), .y(y[12]));
  Fx13 Fx13_inst(.x(x[15]), .y(y[13]));
  Fx14 Fx14_inst(.x({x[17], x[16]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[18], x[16]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[19], x[16]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[20], x[16]}), .y(y[17]));
  Fx18 Fx18_inst(.x(x[21]), .y(y[18]));
  Fx19 Fx19_inst(.x(x[22]), .y(y[19]));
  Fx20 Fx20_inst(.x(x[23]), .y(y[20]));
  Fx21 Fx21_inst(.x({x[25], x[24]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[26], x[24]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[27], x[24]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[28], x[24]}), .y(y[24]));
  Fx25 Fx25_inst(.x(x[29]), .y(y[25]));
  Fx26 Fx26_inst(.x(x[30]), .y(y[26]));
  Fx27 Fx27_inst(.x(x[31]), .y(y[27]));
  Fx28 Fx28_inst(.x({x[33], x[32]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[34], x[32]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[35], x[32]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[36], x[32]}), .y(y[31]));
  Fx32 Fx32_inst(.x(x[37]), .y(y[32]));
  Fx33 Fx33_inst(.x(x[38]), .y(y[33]));
  Fx34 Fx34_inst(.x(x[39]), .y(y[34]));
  Fx35 Fx35_inst(.x({x[41], x[40]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[42], x[40]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[43], x[40]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[44], x[40]}), .y(y[38]));
  Fx39 Fx39_inst(.x(x[45]), .y(y[39]));
  Fx40 Fx40_inst(.x(x[46]), .y(y[40]));
  Fx41 Fx41_inst(.x(x[47]), .y(y[41]));
  Fx42 Fx42_inst(.x({x[49], x[48]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[50], x[48]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[51], x[48]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[52], x[48]}), .y(y[45]));
  Fx46 Fx46_inst(.x(x[53]), .y(y[46]));
  Fx47 Fx47_inst(.x(x[54]), .y(y[47]));
  Fx48 Fx48_inst(.x(x[55]), .y(y[48]));
  Fx49 Fx49_inst(.x({x[57], x[56]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[58], x[56]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[59], x[56]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[60], x[56]}), .y(y[52]));
  Fx53 Fx53_inst(.x(x[61]), .y(y[53]));
  Fx54 Fx54_inst(.x(x[62]), .y(y[54]));
  Fx55 Fx55_inst(.x(x[63]), .y(y[55]));
  Fx56 Fx56_inst(.x({x[65], x[64]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[66], x[64]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[67], x[64]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[68], x[64]}), .y(y[59]));
  Fx60 Fx60_inst(.x(x[69]), .y(y[60]));
  Fx61 Fx61_inst(.x(x[70]), .y(y[61]));
  Fx62 Fx62_inst(.x(x[71]), .y(y[62]));
  Fx63 Fx63_inst(.x({x[73], x[72]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[74], x[72]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[75], x[72]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[76], x[72]}), .y(y[66]));
  Fx67 Fx67_inst(.x(x[77]), .y(y[67]));
  Fx68 Fx68_inst(.x(x[78]), .y(y[68]));
  Fx69 Fx69_inst(.x(x[79]), .y(y[69]));
  Fx70 Fx70_inst(.x({x[83], x[82], x[81], x[80]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[85], x[84], x[81], x[80]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[86], x[82], x[80]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[87], x[84], x[80]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[88], x[82], x[81]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[89], x[84], x[81]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[90], x[84], x[82]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[94], x[93], x[92], x[91]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[96], x[95], x[92], x[91]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[97], x[93], x[91]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[98], x[95], x[91]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[99], x[93], x[92]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[100], x[95], x[92]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[101], x[95], x[93]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[105], x[104], x[103], x[102]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[107], x[106], x[103], x[102]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[108], x[104], x[102]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[109], x[106], x[102]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[110], x[104], x[103]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[111], x[106], x[103]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[112], x[106], x[104]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[116], x[115], x[114], x[113]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[118], x[117], x[114], x[113]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[119], x[115], x[113]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[120], x[117], x[113]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[121], x[115], x[114]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[122], x[117], x[114]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[123], x[117], x[115]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[127], x[126], x[125], x[124]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[129], x[128], x[125], x[124]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[130], x[126], x[124]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[131], x[128], x[124]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[132], x[126], x[125]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[133], x[128], x[125]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[134], x[128], x[126]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[138], x[137], x[136], x[135]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[140], x[139], x[136], x[135]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[141], x[137], x[135]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[142], x[139], x[135]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[143], x[137], x[136]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[144], x[139], x[136]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[145], x[139], x[137]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[149], x[148], x[147], x[146]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[151], x[150], x[147], x[146]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[152], x[148], x[146]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[153], x[150], x[146]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[154], x[148], x[147]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[155], x[150], x[147]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[156], x[150], x[148]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[160], x[159], x[158], x[157]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[162], x[161], x[158], x[157]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[163], x[159], x[157]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[164], x[161], x[157]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[165], x[159], x[158]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[166], x[161], x[158]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[167], x[161], x[159]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[171], x[170], x[169], x[168]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[173], x[172], x[169], x[168]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[174], x[170], x[168]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[175], x[172], x[168]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[176], x[170], x[169]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[177], x[172], x[169]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[178], x[172], x[170]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[182], x[181], x[180], x[179]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[184], x[183], x[180], x[179]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[185], x[181], x[179]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[186], x[183], x[179]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[187], x[181], x[180]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[188], x[183], x[180]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[189], x[183], x[181]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[193], x[192], x[191], x[190]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[195], x[194], x[191], x[190]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[196], x[192], x[190]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[197], x[194], x[190]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[198], x[192], x[191]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[199], x[194], x[191]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[200], x[194], x[192]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[204], x[203], x[202], x[201]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[206], x[205], x[202], x[201]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[207], x[203], x[201]}), .y(y[149]));
  Fx150 Fx150_inst(.x({x[208], x[205], x[201]}), .y(y[150]));
  Fx151 Fx151_inst(.x({x[209], x[203], x[202]}), .y(y[151]));
  Fx152 Fx152_inst(.x({x[210], x[205], x[202]}), .y(y[152]));
  Fx153 Fx153_inst(.x({x[211], x[205], x[203]}), .y(y[153]));
  Fx154 Fx154_inst(.x({x[215], x[214], x[213], x[212]}), .y(y[154]));
  Fx155 Fx155_inst(.x({x[217], x[216], x[213], x[212]}), .y(y[155]));
  Fx156 Fx156_inst(.x({x[218], x[214], x[212]}), .y(y[156]));
  Fx157 Fx157_inst(.x({x[219], x[216], x[212]}), .y(y[157]));
  Fx158 Fx158_inst(.x({x[220], x[214], x[213]}), .y(y[158]));
  Fx159 Fx159_inst(.x({x[221], x[216], x[213]}), .y(y[159]));
  Fx160 Fx160_inst(.x({x[222], x[216], x[214]}), .y(y[160]));
  Fx161 Fx161_inst(.x({x[226], x[225], x[224], x[223]}), .y(y[161]));
  Fx162 Fx162_inst(.x({x[228], x[227], x[224], x[223]}), .y(y[162]));
  Fx163 Fx163_inst(.x({x[229], x[225], x[223]}), .y(y[163]));
  Fx164 Fx164_inst(.x({x[230], x[227], x[223]}), .y(y[164]));
  Fx165 Fx165_inst(.x({x[231], x[225], x[224]}), .y(y[165]));
  Fx166 Fx166_inst(.x({x[232], x[227], x[224]}), .y(y[166]));
  Fx167 Fx167_inst(.x({x[233], x[227], x[225]}), .y(y[167]));
  Fx168 Fx168_inst(.x({x[237], x[236], x[235], x[234]}), .y(y[168]));
  Fx169 Fx169_inst(.x({x[239], x[238], x[235], x[234]}), .y(y[169]));
  Fx170 Fx170_inst(.x({x[240], x[236], x[234]}), .y(y[170]));
  Fx171 Fx171_inst(.x({x[241], x[238], x[234]}), .y(y[171]));
  Fx172 Fx172_inst(.x({x[242], x[236], x[235]}), .y(y[172]));
  Fx173 Fx173_inst(.x({x[243], x[238], x[235]}), .y(y[173]));
  Fx174 Fx174_inst(.x({x[244], x[238], x[236]}), .y(y[174]));
  Fx175 Fx175_inst(.x({x[248], x[247], x[246], x[245]}), .y(y[175]));
  Fx176 Fx176_inst(.x({x[250], x[249], x[246], x[245]}), .y(y[176]));
  Fx177 Fx177_inst(.x({x[251], x[247], x[245]}), .y(y[177]));
  Fx178 Fx178_inst(.x({x[252], x[249], x[245]}), .y(y[178]));
  Fx179 Fx179_inst(.x({x[253], x[247], x[246]}), .y(y[179]));
  Fx180 Fx180_inst(.x({x[254], x[249], x[246]}), .y(y[180]));
  Fx181 Fx181_inst(.x({x[255], x[249], x[247]}), .y(y[181]));
endmodule

module R1ind0(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [56:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~x[0] & t[12];
  assign t[10] = ~x[0] & t[17];
  assign t[11] = ~x[0] & t[18];
  assign t[12] = t[19] ^ x[8];
  assign t[13] = t[20] ^ x[16];
  assign t[14] = t[21] ^ x[24];
  assign t[15] = t[22] ^ x[32];
  assign t[16] = t[23] ^ x[40];
  assign t[17] = t[24] ^ x[48];
  assign t[18] = t[25] ^ x[56];
  assign t[19] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[20] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign t[21] = (x[17] & x[18] & x[19] & ~x[22] & ~x[23]) | (x[17] & x[18] & x[20] & ~x[21] & ~x[23]) | (x[17] & x[19] & x[20] & ~x[22] & ~x[23]) | (~x[18] & x[19] & x[20] & x[21] & ~x[23]) | (x[18] & x[19] & x[20] & ~x[22]) | (x[18] & x[20] & x[21] & ~x[22]) | (x[17] & x[19] & ~x[21] & x[22]);
  assign t[22] = (x[25] & x[26] & x[27] & ~x[30] & ~x[31]) | (x[25] & x[26] & x[28] & ~x[29] & ~x[31]) | (x[25] & x[27] & x[28] & ~x[30] & ~x[31]) | (~x[26] & x[27] & x[28] & x[29] & ~x[31]) | (x[26] & x[27] & x[28] & ~x[30]) | (x[26] & x[28] & x[29] & ~x[30]) | (x[25] & x[27] & ~x[29] & x[30]);
  assign t[23] = (x[33] & x[34] & x[35] & ~x[38] & ~x[39]) | (x[33] & x[34] & x[36] & ~x[37] & ~x[39]) | (x[33] & x[35] & x[36] & ~x[38] & ~x[39]) | (~x[34] & x[35] & x[36] & x[37] & ~x[39]) | (x[34] & x[35] & x[36] & ~x[38]) | (x[34] & x[36] & x[37] & ~x[38]) | (x[33] & x[35] & ~x[37] & x[38]);
  assign t[24] = (x[41] & x[42] & x[43] & ~x[46] & ~x[47]) | (x[41] & x[42] & x[44] & ~x[45] & ~x[47]) | (x[41] & x[43] & x[44] & ~x[46] & ~x[47]) | (~x[42] & x[43] & x[44] & x[45] & ~x[47]) | (x[42] & x[43] & x[44] & ~x[46]) | (x[42] & x[44] & x[45] & ~x[46]) | (x[41] & x[43] & ~x[45] & x[46]);
  assign t[25] = (x[49] & x[50] & x[51] & ~x[54] & ~x[55]) | (x[49] & x[50] & x[52] & ~x[53] & ~x[55]) | (x[49] & x[51] & x[52] & ~x[54] & ~x[55]) | (~x[50] & x[51] & x[52] & x[53] & ~x[55]) | (x[50] & x[51] & x[52] & ~x[54]) | (x[50] & x[52] & x[53] & ~x[54]) | (x[49] & x[51] & ~x[53] & x[54]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[7]);
  assign t[4] = ~(~x[0] & ~t[13]);
  assign t[5] = ~x[0] & t[14];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~x[0] & t[15];
  assign t[9] = ~(~x[0] & ~t[16]);
  assign y = t[0] & t[1];
endmodule

module R1ind66(x, y);
 input [8:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = t[2] ^ x[8];
  assign t[2] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~(t[0]);
endmodule

module R1ind67(x, y);
 input [16:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[2];
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = t[6] ^ x[16];
  assign t[5] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[6] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind68(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [16:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~x[0] & t[2];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = t[4] ^ x[8];
  assign t[3] = t[5] ^ x[16];
  assign t[4] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[5] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind73(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind74(x, y);
 input [16:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~(~x[0] & ~t[2]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = t[4] ^ x[8];
  assign t[3] = t[5] ^ x[16];
  assign t[4] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[5] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [22:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[19];
  assign t[14] = t[19] ^ x[20];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[22];
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[19] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[21] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[13] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] | t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind76(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind77(x, y);
 input [22:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[19];
  assign t[14] = t[19] ^ x[20];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[22];
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[19] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind78(x, y);
 input [22:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[19];
  assign t[15] = t[20] ^ x[20];
  assign t[16] = t[21] ^ x[21];
  assign t[17] = t[22] ^ x[22];
  assign t[18] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[21] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[22] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind79(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[22] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[23] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind80(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind81(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[22] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[23] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind82(x, y);
 input [22:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[19];
  assign t[15] = t[20] ^ x[20];
  assign t[16] = t[21] ^ x[21];
  assign t[17] = t[22] ^ x[22];
  assign t[18] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[21] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[22] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind83(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[22] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[23] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind84(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind85(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[22] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[23] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind86(x, y);
 input [22:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[19];
  assign t[15] = t[20] ^ x[20];
  assign t[16] = t[21] ^ x[21];
  assign t[17] = t[22] ^ x[22];
  assign t[18] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[21] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[22] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind87(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[22] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[23] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind88(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind89(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[22] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[23] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind90(x, y);
 input [22:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[19];
  assign t[15] = t[20] ^ x[20];
  assign t[16] = t[21] ^ x[21];
  assign t[17] = t[22] ^ x[22];
  assign t[18] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[21] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[22] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind91(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[22] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[23] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind92(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind93(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[22] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[23] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind94(x, y);
 input [22:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[19];
  assign t[15] = t[20] ^ x[20];
  assign t[16] = t[21] ^ x[21];
  assign t[17] = t[22] ^ x[22];
  assign t[18] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[21] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[22] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind95(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[22] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[23] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind96(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind97(x, y);
 input [22:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[19];
  assign t[14] = t[19] ^ x[20];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[22];
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[19] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind98(x, y);
 input [22:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15]);
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[19];
  assign t[13] = t[18] ^ x[20];
  assign t[14] = t[19] ^ x[21];
  assign t[15] = t[20] ^ x[22];
  assign t[16] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[17] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[18] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[11];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = t[9] | t[12];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[10] | t[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind99(x, y);
 input [22:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[19];
  assign t[14] = t[19] ^ x[20];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[22];
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[19] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[21] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[13] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] | t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind100(x, y);
 input [21:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~t[2];
  assign t[10] = t[14] ^ x[11];
  assign t[11] = t[15] ^ x[19];
  assign t[12] = t[16] ^ x[20];
  assign t[13] = t[17] ^ x[21];
  assign t[14] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[15] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[16] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[17] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[10];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[11] & t[7]);
  assign t[6] = ~(t[12] & t[8]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[13] & t[9]);
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind101(x, y);
 input [22:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[19];
  assign t[14] = t[19] ^ x[20];
  assign t[15] = t[20] ^ x[21];
  assign t[16] = t[21] ^ x[22];
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[19] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind102(x, y);
 input [22:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15]);
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[19];
  assign t[13] = t[18] ^ x[20];
  assign t[14] = t[19] ^ x[21];
  assign t[15] = t[20] ^ x[22];
  assign t[16] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[17] = (x[12] & x[13] & ~x[15] & x[16] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[12] & x[13] & ~x[14] & x[17] & ~x[18]) | (x[12] & ~x[15] & x[16] & x[17] & ~x[18]) | (x[12] & ~x[14] & x[15] & x[16]) | (x[13] & x[14] & ~x[15] & x[17]) | (x[13] & ~x[15] & x[16] & x[17]);
  assign t[18] = (x[13] & ~x[14] & x[15] & ~x[16] & x[17]) | (x[13] & ~x[14] & x[15] & ~x[16] & x[18]) | (x[13] & ~x[14] & ~x[16] & x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[12] & ~x[14] & x[15] & x[18]) | (x[12] & ~x[16] & x[17] & x[18]) | (x[15] & x[17] & x[18]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[14] & ~x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[15] & ~x[17] & x[18]) | (x[12] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[12] & x[14] & x[15] & x[16] & x[17]) | (x[13] & x[14] & ~x[15] & x[18]) | (x[13] & x[16] & ~x[17] & x[18]) | (x[14] & x[16] & x[18]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[11];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = t[9] | t[12];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[10] | t[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind103(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[22] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[23] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind104(x, y);
 input [21:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = t[18] ^ x[20];
  assign t[15] = t[19] ^ x[21];
  assign t[16] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[17] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[18] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[19] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind105(x, y);
 input [22:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = t[22] ^ x[21];
  assign t[18] = t[23] ^ x[22];
  assign t[19] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[21] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[22] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[23] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind106(x, y);
 input [22:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[19];
  assign t[15] = t[20] ^ x[20];
  assign t[16] = t[21] ^ x[21];
  assign t[17] = t[22] ^ x[22];
  assign t[18] = (x[4] & x[5] & ~x[7] & x[8] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[4] & x[5] & ~x[6] & x[9] & ~x[10]) | (x[4] & ~x[7] & x[8] & x[9] & ~x[10]) | (x[4] & ~x[6] & x[7] & x[8]) | (x[5] & x[6] & ~x[7] & x[9]) | (x[5] & ~x[7] & x[8] & x[9]);
  assign t[19] = (x[12] & x[13] & x[14] & ~x[17] & ~x[18]) | (x[12] & x[13] & x[15] & ~x[16] & ~x[18]) | (x[12] & x[14] & x[15] & ~x[17] & ~x[18]) | (~x[13] & x[14] & x[15] & x[16] & ~x[18]) | (x[13] & x[14] & x[15] & ~x[17]) | (x[13] & x[15] & x[16] & ~x[17]) | (x[12] & x[14] & ~x[16] & x[17]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[5] & ~x[6] & x[7] & ~x[8] & x[9]) | (x[5] & ~x[6] & x[7] & ~x[8] & x[10]) | (x[5] & ~x[6] & ~x[8] & x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[4] & ~x[6] & x[7] & x[10]) | (x[4] & ~x[8] & x[9] & x[10]) | (x[7] & x[9] & x[10]);
  assign t[21] = (x[4] & x[5] & x[6] & ~x[9] & ~x[10]) | (x[4] & x[5] & x[7] & ~x[8] & ~x[10]) | (x[4] & x[6] & x[7] & ~x[9] & ~x[10]) | (~x[5] & x[6] & x[7] & x[8] & ~x[10]) | (x[5] & x[6] & x[7] & ~x[9]) | (x[5] & x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[8] & x[9]);
  assign t[22] = (x[4] & x[6] & ~x[7] & x[8] & ~x[9]) | (x[4] & x[6] & ~x[7] & ~x[9] & x[10]) | (x[4] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[4] & x[6] & x[7] & x[8] & x[9]) | (x[5] & x[6] & ~x[7] & x[10]) | (x[5] & x[8] & ~x[9] & x[10]) | (x[6] & x[8] & x[10]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind107(x, y);
 input [34:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[26] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[27] | t[20]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[20];
  assign t[27] = t[36] ^ x[28];
  assign t[28] = t[37] ^ x[29];
  assign t[29] = t[38] ^ x[30];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[31];
  assign t[31] = t[40] ^ x[32];
  assign t[32] = t[41] ^ x[33];
  assign t[33] = t[42] ^ x[34];
  assign t[34] = (x[5] & x[6] & x[7] & ~x[10] & ~x[11]) | (x[5] & x[6] & x[8] & ~x[9] & ~x[11]) | (x[5] & x[7] & x[8] & ~x[10] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[6] & x[7] & x[8] & ~x[10]) | (x[6] & x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[9] & x[10]);
  assign t[35] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[36] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[37] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[38] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[41] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[42] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind108(x, y);
 input [32:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[21] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[24] & t[17]);
  assign t[15] = ~(t[25]);
  assign t[16] = ~(t[25] & t[18]);
  assign t[17] = ~(t[20]);
  assign t[18] = ~(t[22]);
  assign t[19] = t[26] ^ x[10];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = t[27] ^ x[20];
  assign t[21] = t[28] ^ x[21];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = t[30] ^ x[30];
  assign t[24] = t[31] ^ x[31];
  assign t[25] = t[32] ^ x[32];
  assign t[26] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[27] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[28] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[29] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[31] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[32] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[3] = ~x[2] & t[19];
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[11] : t[7];
  assign t[6] = x[2] ? x[12] : t[8];
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[20] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind109(x, y);
 input [34:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[26]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[29] & t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[31] & t[30]);
  assign t[24] = ~(t[33]);
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[20];
  assign t[27] = t[36] ^ x[28];
  assign t[28] = t[37] ^ x[29];
  assign t[29] = t[38] ^ x[30];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[31];
  assign t[31] = t[40] ^ x[32];
  assign t[32] = t[41] ^ x[33];
  assign t[33] = t[42] ^ x[34];
  assign t[34] = (x[5] & x[6] & x[7] & ~x[10] & ~x[11]) | (x[5] & x[6] & x[8] & ~x[9] & ~x[11]) | (x[5] & x[7] & x[8] & ~x[10] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[6] & x[7] & x[8] & ~x[10]) | (x[6] & x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[9] & x[10]);
  assign t[35] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[36] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[37] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[38] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[39] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[41] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[42] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind110(x, y);
 input [34:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = t[17] | t[24];
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = t[20] | t[25];
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[21] | t[15]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[29]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[22] | t[18]);
  assign t[21] = ~(t[30]);
  assign t[22] = ~(t[31]);
  assign t[23] = t[32] ^ x[12];
  assign t[24] = t[33] ^ x[20];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[29];
  assign t[27] = t[36] ^ x[30];
  assign t[28] = t[37] ^ x[31];
  assign t[29] = t[38] ^ x[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[33];
  assign t[31] = t[40] ^ x[34];
  assign t[32] = (x[5] & x[6] & x[7] & ~x[10] & ~x[11]) | (x[5] & x[6] & x[8] & ~x[9] & ~x[11]) | (x[5] & x[7] & x[8] & ~x[10] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[6] & x[7] & x[8] & ~x[10]) | (x[6] & x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[9] & x[10]);
  assign t[33] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[34] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[35] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[36] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[37] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind111(x, y);
 input [34:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[24] | t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[25] | t[18]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[27]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[30]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = t[32] ^ x[10];
  assign t[24] = t[33] ^ x[20];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[29];
  assign t[27] = t[36] ^ x[30];
  assign t[28] = t[37] ^ x[31];
  assign t[29] = t[38] ^ x[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[33];
  assign t[31] = t[40] ^ x[34];
  assign t[32] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[33] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[34] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[35] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[36] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[37] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[38] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[39] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[3] = ~x[2] & t[23];
  assign t[40] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[11] : t[7];
  assign t[6] = x[2] ? x[12] : t[8];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13] | t[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind112(x, y);
 input [32:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25] & t[18]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[26] & t[19]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[27] & t[20]);
  assign t[19] = ~(t[22]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[24]);
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[20];
  assign t[23] = t[30] ^ x[21];
  assign t[24] = t[31] ^ x[29];
  assign t[25] = t[32] ^ x[30];
  assign t[26] = t[33] ^ x[31];
  assign t[27] = t[34] ^ x[32];
  assign t[28] = (x[5] & x[6] & x[7] & ~x[10] & ~x[11]) | (x[5] & x[6] & x[8] & ~x[9] & ~x[11]) | (x[5] & x[7] & x[8] & ~x[10] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[6] & x[7] & x[8] & ~x[10]) | (x[6] & x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[9] & x[10]);
  assign t[29] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[31] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[32] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[33] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[34] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[21];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind113(x, y);
 input [34:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[26]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[29] & t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[31] & t[30]);
  assign t[24] = ~(t[33]);
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[20];
  assign t[27] = t[36] ^ x[28];
  assign t[28] = t[37] ^ x[29];
  assign t[29] = t[38] ^ x[30];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[31];
  assign t[31] = t[40] ^ x[32];
  assign t[32] = t[41] ^ x[33];
  assign t[33] = t[42] ^ x[34];
  assign t[34] = (x[5] & x[6] & x[7] & ~x[10] & ~x[11]) | (x[5] & x[6] & x[8] & ~x[9] & ~x[11]) | (x[5] & x[7] & x[8] & ~x[10] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[6] & x[7] & x[8] & ~x[10]) | (x[6] & x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[9] & x[10]);
  assign t[35] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[36] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[37] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[38] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[39] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[41] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[42] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind114(x, y);
 input [34:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~t[2];
  assign t[10] = t[15] | t[22];
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = t[18] | t[23];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[19] | t[13]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[20] | t[16]);
  assign t[19] = ~(t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[29]);
  assign t[21] = t[30] ^ x[10];
  assign t[22] = t[31] ^ x[20];
  assign t[23] = t[32] ^ x[28];
  assign t[24] = t[33] ^ x[29];
  assign t[25] = t[34] ^ x[30];
  assign t[26] = t[35] ^ x[31];
  assign t[27] = t[36] ^ x[32];
  assign t[28] = t[37] ^ x[33];
  assign t[29] = t[38] ^ x[34];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[31] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[32] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[33] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[34] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[35] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[36] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[37] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[38] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~x[2] & t[21];
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[11] : t[7];
  assign t[6] = x[2] ? x[12] : t[8];
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind115(x, y);
 input [42:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[28] | t[19]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[30] | t[22]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[37] ^ x[10];
  assign t[28] = t[38] ^ x[20];
  assign t[29] = t[39] ^ x[28];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[36];
  assign t[31] = t[41] ^ x[37];
  assign t[32] = t[42] ^ x[38];
  assign t[33] = t[43] ^ x[39];
  assign t[34] = t[44] ^ x[40];
  assign t[35] = t[45] ^ x[41];
  assign t[36] = t[46] ^ x[42];
  assign t[37] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[38] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[39] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[41] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[42] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[43] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[44] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[45] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[46] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[4] = ~(~x[2] & ~t[27]);
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind116(x, y);
 input [40:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[24] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[27] & t[19]);
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[29] & t[21]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[30] & t[22]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[27]);
  assign t[23] = t[31] ^ x[10];
  assign t[24] = t[32] ^ x[20];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[29];
  assign t[27] = t[35] ^ x[37];
  assign t[28] = t[36] ^ x[38];
  assign t[29] = t[37] ^ x[39];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[38] ^ x[40];
  assign t[31] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[32] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[33] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[34] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[35] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[36] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[37] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[38] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[4] = ~x[2] & t[23];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind117(x, y);
 input [42:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[28]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[30]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[32] & t[31]);
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[34] & t[33]);
  assign t[26] = ~(t[36]);
  assign t[27] = t[37] ^ x[10];
  assign t[28] = t[38] ^ x[20];
  assign t[29] = t[39] ^ x[28];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[36];
  assign t[31] = t[41] ^ x[37];
  assign t[32] = t[42] ^ x[38];
  assign t[33] = t[43] ^ x[39];
  assign t[34] = t[44] ^ x[40];
  assign t[35] = t[45] ^ x[41];
  assign t[36] = t[46] ^ x[42];
  assign t[37] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[38] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[39] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[41] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[42] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[43] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[44] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[45] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[46] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[4] = ~x[2] & t[27];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind118(x, y);
 input [34:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = t[18] | t[24];
  assign t[13] = ~x[2] & t[25];
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = t[21] | t[26];
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[22] | t[16]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[23] | t[19]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[32]);
  assign t[24] = t[33] ^ x[12];
  assign t[25] = t[34] ^ x[20];
  assign t[26] = t[35] ^ x[28];
  assign t[27] = t[36] ^ x[29];
  assign t[28] = t[37] ^ x[30];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[32];
  assign t[31] = t[40] ^ x[33];
  assign t[32] = t[41] ^ x[34];
  assign t[33] = (x[5] & x[6] & ~x[8] & x[9] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[5] & x[6] & ~x[7] & x[10] & ~x[11]) | (x[5] & ~x[8] & x[9] & x[10] & ~x[11]) | (x[5] & ~x[7] & x[8] & x[9]) | (x[6] & x[7] & ~x[8] & x[10]) | (x[6] & ~x[8] & x[9] & x[10]);
  assign t[34] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[35] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[36] = (x[6] & ~x[7] & x[8] & ~x[9] & x[10]) | (x[6] & ~x[7] & x[8] & ~x[9] & x[11]) | (x[6] & ~x[7] & ~x[9] & x[10] & x[11]) | (x[5] & x[7] & x[8] & x[9] & x[10]) | (x[5] & ~x[7] & x[8] & x[11]) | (x[5] & ~x[9] & x[10] & x[11]) | (x[8] & x[10] & x[11]);
  assign t[37] = (x[5] & x[6] & x[7] & ~x[10] & ~x[11]) | (x[5] & x[6] & x[8] & ~x[9] & ~x[11]) | (x[5] & x[7] & x[8] & ~x[10] & ~x[11]) | (~x[6] & x[7] & x[8] & x[9] & ~x[11]) | (x[6] & x[7] & x[8] & ~x[10]) | (x[6] & x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[9] & x[10]);
  assign t[38] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[39] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[3] = t[6] ? x[1] : x[0];
  assign t[40] = (x[5] & x[7] & ~x[8] & x[9] & ~x[10]) | (x[5] & x[7] & ~x[8] & ~x[10] & x[11]) | (x[5] & ~x[8] & x[9] & ~x[10] & x[11]) | (x[5] & x[7] & x[8] & x[9] & x[10]) | (x[6] & x[7] & ~x[8] & x[11]) | (x[6] & x[9] & ~x[10] & x[11]) | (x[7] & x[9] & x[11]);
  assign t[41] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind119(x, y);
 input [42:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[28] | t[19]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[30] | t[22]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[37] ^ x[10];
  assign t[28] = t[38] ^ x[20];
  assign t[29] = t[39] ^ x[28];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[36];
  assign t[31] = t[41] ^ x[37];
  assign t[32] = t[42] ^ x[38];
  assign t[33] = t[43] ^ x[39];
  assign t[34] = t[44] ^ x[40];
  assign t[35] = t[45] ^ x[41];
  assign t[36] = t[46] ^ x[42];
  assign t[37] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[38] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[39] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[41] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[42] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[43] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[44] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[45] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[46] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[4] = ~(~x[2] & ~t[27]);
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind120(x, y);
 input [40:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[24] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[27] & t[19]);
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[29] & t[21]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[30] & t[22]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[27]);
  assign t[23] = t[31] ^ x[10];
  assign t[24] = t[32] ^ x[20];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[29];
  assign t[27] = t[35] ^ x[37];
  assign t[28] = t[36] ^ x[38];
  assign t[29] = t[37] ^ x[39];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[38] ^ x[40];
  assign t[31] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[32] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[33] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[34] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[35] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[36] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[37] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[38] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[4] = ~x[2] & t[23];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind121(x, y);
 input [42:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[28]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[30]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[32] & t[31]);
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[34] & t[33]);
  assign t[26] = ~(t[36]);
  assign t[27] = t[37] ^ x[10];
  assign t[28] = t[38] ^ x[20];
  assign t[29] = t[39] ^ x[28];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[36];
  assign t[31] = t[41] ^ x[37];
  assign t[32] = t[42] ^ x[38];
  assign t[33] = t[43] ^ x[39];
  assign t[34] = t[44] ^ x[40];
  assign t[35] = t[45] ^ x[41];
  assign t[36] = t[46] ^ x[42];
  assign t[37] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[38] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[39] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[41] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[42] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[43] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[44] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[45] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[46] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[4] = ~x[2] & t[27];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind122(x, y);
 input [42:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[26];
  assign t[14] = ~x[2] & t[27];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = t[22] | t[28];
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[23] | t[17]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[24] | t[20]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34]);
  assign t[25] = t[35] ^ x[10];
  assign t[26] = t[36] ^ x[20];
  assign t[27] = t[37] ^ x[28];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[37];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[38];
  assign t[31] = t[41] ^ x[39];
  assign t[32] = t[42] ^ x[40];
  assign t[33] = t[43] ^ x[41];
  assign t[34] = t[44] ^ x[42];
  assign t[35] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[36] = (x[13] & x[14] & ~x[16] & x[17] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[13] & x[14] & ~x[15] & x[18] & ~x[19]) | (x[13] & ~x[16] & x[17] & x[18] & ~x[19]) | (x[13] & ~x[15] & x[16] & x[17]) | (x[14] & x[15] & ~x[16] & x[18]) | (x[14] & ~x[16] & x[17] & x[18]);
  assign t[37] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[38] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[39] = (x[14] & ~x[15] & x[16] & ~x[17] & x[18]) | (x[14] & ~x[15] & x[16] & ~x[17] & x[19]) | (x[14] & ~x[15] & ~x[17] & x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[13] & ~x[15] & x[16] & x[19]) | (x[13] & ~x[17] & x[18] & x[19]) | (x[16] & x[18] & x[19]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[13] & x[14] & x[15] & ~x[18] & ~x[19]) | (x[13] & x[14] & x[16] & ~x[17] & ~x[19]) | (x[13] & x[15] & x[16] & ~x[18] & ~x[19]) | (~x[14] & x[15] & x[16] & x[17] & ~x[19]) | (x[14] & x[15] & x[16] & ~x[18]) | (x[14] & x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[17] & x[18]);
  assign t[41] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[42] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[43] = (x[13] & x[15] & ~x[16] & x[17] & ~x[18]) | (x[13] & x[15] & ~x[16] & ~x[18] & x[19]) | (x[13] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[13] & x[15] & x[16] & x[17] & x[18]) | (x[14] & x[15] & ~x[16] & x[19]) | (x[14] & x[17] & ~x[18] & x[19]) | (x[15] & x[17] & x[19]);
  assign t[44] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[4] = ~x[2] & t[25];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind123(x, y);
 input [46:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[13];
  assign t[36] = t[49] ^ x[21];
  assign t[37] = t[50] ^ x[29];
  assign t[38] = t[51] ^ x[37];
  assign t[39] = t[52] ^ x[38];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[39];
  assign t[41] = t[54] ^ x[40];
  assign t[42] = t[55] ^ x[41];
  assign t[43] = t[56] ^ x[42];
  assign t[44] = t[57] ^ x[43];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = t[59] ^ x[45];
  assign t[47] = t[60] ^ x[46];
  assign t[48] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[49] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[51] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[52] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[53] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[54] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[55] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[56] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[57] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[58] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[59] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind124(x, y);
 input [43:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[22];
  assign t[32] = t[42] ^ x[30];
  assign t[33] = t[43] ^ x[31];
  assign t[34] = t[44] ^ x[39];
  assign t[35] = t[45] ^ x[40];
  assign t[36] = t[46] ^ x[41];
  assign t[37] = t[47] ^ x[42];
  assign t[38] = t[48] ^ x[43];
  assign t[39] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[41] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[42] = (x[23] & x[25] & ~x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[26] & ~x[28] & x[29]) | (x[23] & ~x[26] & x[27] & ~x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[24] & x[25] & ~x[26] & x[29]) | (x[24] & x[27] & ~x[28] & x[29]) | (x[25] & x[27] & x[29]);
  assign t[43] = (x[23] & x[24] & x[25] & ~x[28] & ~x[29]) | (x[23] & x[24] & x[26] & ~x[27] & ~x[29]) | (x[23] & x[25] & x[26] & ~x[28] & ~x[29]) | (~x[24] & x[25] & x[26] & x[27] & ~x[29]) | (x[24] & x[25] & x[26] & ~x[28]) | (x[24] & x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[27] & x[28]);
  assign t[44] = (x[32] & x[34] & ~x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[35] & ~x[37] & x[38]) | (x[32] & ~x[35] & x[36] & ~x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[33] & x[34] & ~x[35] & x[38]) | (x[33] & x[36] & ~x[37] & x[38]) | (x[34] & x[36] & x[38]);
  assign t[45] = (x[32] & x[33] & x[34] & ~x[37] & ~x[38]) | (x[32] & x[33] & x[35] & ~x[36] & ~x[38]) | (x[32] & x[34] & x[35] & ~x[37] & ~x[38]) | (~x[33] & x[34] & x[35] & x[36] & ~x[38]) | (x[33] & x[34] & x[35] & ~x[37]) | (x[33] & x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[36] & x[37]);
  assign t[46] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[47] = (x[24] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[24] & ~x[25] & x[26] & ~x[27] & x[29]) | (x[24] & ~x[25] & ~x[27] & x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[23] & ~x[25] & x[26] & x[29]) | (x[23] & ~x[27] & x[28] & x[29]) | (x[26] & x[28] & x[29]);
  assign t[48] = (x[33] & ~x[34] & x[35] & ~x[36] & x[37]) | (x[33] & ~x[34] & x[35] & ~x[36] & x[38]) | (x[33] & ~x[34] & ~x[36] & x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[32] & ~x[34] & x[35] & x[38]) | (x[32] & ~x[36] & x[37] & x[38]) | (x[35] & x[37] & x[38]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind125(x, y);
 input [46:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = ~(t[22] & t[36]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[37]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] & t[34]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[44] & t[43]);
  assign t[34] = ~(t[47]);
  assign t[35] = t[48] ^ x[13];
  assign t[36] = t[49] ^ x[21];
  assign t[37] = t[50] ^ x[29];
  assign t[38] = t[51] ^ x[37];
  assign t[39] = t[52] ^ x[38];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[39];
  assign t[41] = t[54] ^ x[40];
  assign t[42] = t[55] ^ x[41];
  assign t[43] = t[56] ^ x[42];
  assign t[44] = t[57] ^ x[43];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = t[59] ^ x[45];
  assign t[47] = t[60] ^ x[46];
  assign t[48] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[49] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[51] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[52] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[53] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[54] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[55] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[56] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[57] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[58] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[59] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind126(x, y);
 input [46:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[13];
  assign t[33] = t[46] ^ x[21];
  assign t[34] = t[47] ^ x[29];
  assign t[35] = t[48] ^ x[37];
  assign t[36] = t[49] ^ x[38];
  assign t[37] = t[50] ^ x[39];
  assign t[38] = t[51] ^ x[40];
  assign t[39] = t[52] ^ x[41];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[42];
  assign t[41] = t[54] ^ x[43];
  assign t[42] = t[55] ^ x[44];
  assign t[43] = t[56] ^ x[45];
  assign t[44] = t[57] ^ x[46];
  assign t[45] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[46] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[47] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[48] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[49] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[4] = t[7];
  assign t[50] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[51] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[52] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[53] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[54] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[55] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[56] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[57] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind127(x, y);
 input [46:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[13];
  assign t[36] = t[49] ^ x[21];
  assign t[37] = t[50] ^ x[29];
  assign t[38] = t[51] ^ x[37];
  assign t[39] = t[52] ^ x[38];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[39];
  assign t[41] = t[54] ^ x[40];
  assign t[42] = t[55] ^ x[41];
  assign t[43] = t[56] ^ x[42];
  assign t[44] = t[57] ^ x[43];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = t[59] ^ x[45];
  assign t[47] = t[60] ^ x[46];
  assign t[48] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[49] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[51] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[52] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[53] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[54] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[55] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[56] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[57] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[58] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[59] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind128(x, y);
 input [43:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[28] & t[18]);
  assign t[13] = ~(t[29] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[34] & t[24]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[35] & t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = ~(t[36] & t[26]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[30]);
  assign t[26] = ~(t[32]);
  assign t[27] = t[37] ^ x[10];
  assign t[28] = t[38] ^ x[21];
  assign t[29] = t[39] ^ x[22];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[30];
  assign t[31] = t[41] ^ x[31];
  assign t[32] = t[42] ^ x[39];
  assign t[33] = t[43] ^ x[40];
  assign t[34] = t[44] ^ x[41];
  assign t[35] = t[45] ^ x[42];
  assign t[36] = t[46] ^ x[43];
  assign t[37] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[38] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[39] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[3] = ~x[2] & t[27];
  assign t[40] = (x[23] & x[25] & ~x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[26] & ~x[28] & x[29]) | (x[23] & ~x[26] & x[27] & ~x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[24] & x[25] & ~x[26] & x[29]) | (x[24] & x[27] & ~x[28] & x[29]) | (x[25] & x[27] & x[29]);
  assign t[41] = (x[23] & x[24] & x[25] & ~x[28] & ~x[29]) | (x[23] & x[24] & x[26] & ~x[27] & ~x[29]) | (x[23] & x[25] & x[26] & ~x[28] & ~x[29]) | (~x[24] & x[25] & x[26] & x[27] & ~x[29]) | (x[24] & x[25] & x[26] & ~x[28]) | (x[24] & x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[27] & x[28]);
  assign t[42] = (x[32] & x[34] & ~x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[35] & ~x[37] & x[38]) | (x[32] & ~x[35] & x[36] & ~x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[33] & x[34] & ~x[35] & x[38]) | (x[33] & x[36] & ~x[37] & x[38]) | (x[34] & x[36] & x[38]);
  assign t[43] = (x[32] & x[33] & x[34] & ~x[37] & ~x[38]) | (x[32] & x[33] & x[35] & ~x[36] & ~x[38]) | (x[32] & x[34] & x[35] & ~x[37] & ~x[38]) | (~x[33] & x[34] & x[35] & x[36] & ~x[38]) | (x[33] & x[34] & x[35] & ~x[37]) | (x[33] & x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[36] & x[37]);
  assign t[44] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[45] = (x[24] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[24] & ~x[25] & x[26] & ~x[27] & x[29]) | (x[24] & ~x[25] & ~x[27] & x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[23] & ~x[25] & x[26] & x[29]) | (x[23] & ~x[27] & x[28] & x[29]) | (x[26] & x[28] & x[29]);
  assign t[46] = (x[33] & ~x[34] & x[35] & ~x[36] & x[37]) | (x[33] & ~x[34] & x[35] & ~x[36] & x[38]) | (x[33] & ~x[34] & ~x[36] & x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[32] & ~x[34] & x[35] & x[38]) | (x[32] & ~x[36] & x[37] & x[38]) | (x[35] & x[37] & x[38]);
  assign t[4] = t[6];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = x[2] ? x[12] : t[10];
  assign t[8] = x[2] ? x[13] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind129(x, y);
 input [46:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = ~(t[20] & t[34]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = ~(t[23] & t[35]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26] & t[36]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] & t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] & t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[38] & t[37]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[45]);
  assign t[33] = t[46] ^ x[10];
  assign t[34] = t[47] ^ x[21];
  assign t[35] = t[48] ^ x[29];
  assign t[36] = t[49] ^ x[37];
  assign t[37] = t[50] ^ x[38];
  assign t[38] = t[51] ^ x[39];
  assign t[39] = t[52] ^ x[40];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[41];
  assign t[41] = t[54] ^ x[42];
  assign t[42] = t[55] ^ x[43];
  assign t[43] = t[56] ^ x[44];
  assign t[44] = t[57] ^ x[45];
  assign t[45] = t[58] ^ x[46];
  assign t[46] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[47] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[48] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[49] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[4] = t[6];
  assign t[50] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[51] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[52] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[53] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[54] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[55] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[56] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[57] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[58] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = x[2] ? x[12] : t[10];
  assign t[8] = x[2] ? x[13] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind130(x, y);
 input [46:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[13];
  assign t[33] = t[46] ^ x[21];
  assign t[34] = t[47] ^ x[29];
  assign t[35] = t[48] ^ x[37];
  assign t[36] = t[49] ^ x[38];
  assign t[37] = t[50] ^ x[39];
  assign t[38] = t[51] ^ x[40];
  assign t[39] = t[52] ^ x[41];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[42];
  assign t[41] = t[54] ^ x[43];
  assign t[42] = t[55] ^ x[44];
  assign t[43] = t[56] ^ x[45];
  assign t[44] = t[57] ^ x[46];
  assign t[45] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[46] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[47] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[48] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[49] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[4] = t[7];
  assign t[50] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[51] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[52] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[53] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[54] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[55] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[56] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[57] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind131(x, y);
 input [46:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[18] | t[19]);
  assign t[13] = ~(t[34] | t[20]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[15] = ~(t[35] | t[23]);
  assign t[16] = ~(t[24] | t[25]);
  assign t[17] = ~(t[36] | t[26]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] | t[32]);
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[37] | t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = t[46] ^ x[10];
  assign t[34] = t[47] ^ x[21];
  assign t[35] = t[48] ^ x[29];
  assign t[36] = t[49] ^ x[37];
  assign t[37] = t[50] ^ x[38];
  assign t[38] = t[51] ^ x[39];
  assign t[39] = t[52] ^ x[40];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[41];
  assign t[41] = t[54] ^ x[42];
  assign t[42] = t[55] ^ x[43];
  assign t[43] = t[56] ^ x[44];
  assign t[44] = t[57] ^ x[45];
  assign t[45] = t[58] ^ x[46];
  assign t[46] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[47] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[48] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[49] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[4] = t[6];
  assign t[50] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[51] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[52] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[53] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[54] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[55] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[56] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[57] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[58] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = x[2] ? x[12] : t[10];
  assign t[8] = x[2] ? x[13] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind132(x, y);
 input [43:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[22];
  assign t[32] = t[42] ^ x[30];
  assign t[33] = t[43] ^ x[31];
  assign t[34] = t[44] ^ x[39];
  assign t[35] = t[45] ^ x[40];
  assign t[36] = t[46] ^ x[41];
  assign t[37] = t[47] ^ x[42];
  assign t[38] = t[48] ^ x[43];
  assign t[39] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[41] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[42] = (x[23] & x[25] & ~x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[26] & ~x[28] & x[29]) | (x[23] & ~x[26] & x[27] & ~x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[24] & x[25] & ~x[26] & x[29]) | (x[24] & x[27] & ~x[28] & x[29]) | (x[25] & x[27] & x[29]);
  assign t[43] = (x[23] & x[24] & x[25] & ~x[28] & ~x[29]) | (x[23] & x[24] & x[26] & ~x[27] & ~x[29]) | (x[23] & x[25] & x[26] & ~x[28] & ~x[29]) | (~x[24] & x[25] & x[26] & x[27] & ~x[29]) | (x[24] & x[25] & x[26] & ~x[28]) | (x[24] & x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[27] & x[28]);
  assign t[44] = (x[32] & x[34] & ~x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[35] & ~x[37] & x[38]) | (x[32] & ~x[35] & x[36] & ~x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[33] & x[34] & ~x[35] & x[38]) | (x[33] & x[36] & ~x[37] & x[38]) | (x[34] & x[36] & x[38]);
  assign t[45] = (x[32] & x[33] & x[34] & ~x[37] & ~x[38]) | (x[32] & x[33] & x[35] & ~x[36] & ~x[38]) | (x[32] & x[34] & x[35] & ~x[37] & ~x[38]) | (~x[33] & x[34] & x[35] & x[36] & ~x[38]) | (x[33] & x[34] & x[35] & ~x[37]) | (x[33] & x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[36] & x[37]);
  assign t[46] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[47] = (x[24] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[24] & ~x[25] & x[26] & ~x[27] & x[29]) | (x[24] & ~x[25] & ~x[27] & x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[23] & ~x[25] & x[26] & x[29]) | (x[23] & ~x[27] & x[28] & x[29]) | (x[26] & x[28] & x[29]);
  assign t[48] = (x[33] & ~x[34] & x[35] & ~x[36] & x[37]) | (x[33] & ~x[34] & x[35] & ~x[36] & x[38]) | (x[33] & ~x[34] & ~x[36] & x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[32] & ~x[34] & x[35] & x[38]) | (x[32] & ~x[36] & x[37] & x[38]) | (x[35] & x[37] & x[38]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind133(x, y);
 input [46:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = ~(t[22] & t[36]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[37]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] & t[34]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[44] & t[43]);
  assign t[34] = ~(t[47]);
  assign t[35] = t[48] ^ x[13];
  assign t[36] = t[49] ^ x[21];
  assign t[37] = t[50] ^ x[29];
  assign t[38] = t[51] ^ x[37];
  assign t[39] = t[52] ^ x[38];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[39];
  assign t[41] = t[54] ^ x[40];
  assign t[42] = t[55] ^ x[41];
  assign t[43] = t[56] ^ x[42];
  assign t[44] = t[57] ^ x[43];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = t[59] ^ x[45];
  assign t[47] = t[60] ^ x[46];
  assign t[48] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[49] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[51] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[52] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[53] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[54] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[55] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[56] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[57] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[58] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[59] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind134(x, y);
 input [46:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = t[20] | t[31];
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = t[23] | t[32];
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = t[26] | t[33];
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[35]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] | t[18]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[28] | t[21]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[29] | t[24]);
  assign t[27] = ~(t[40]);
  assign t[28] = ~(t[41]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ x[10];
  assign t[31] = t[44] ^ x[21];
  assign t[32] = t[45] ^ x[29];
  assign t[33] = t[46] ^ x[37];
  assign t[34] = t[47] ^ x[38];
  assign t[35] = t[48] ^ x[39];
  assign t[36] = t[49] ^ x[40];
  assign t[37] = t[50] ^ x[41];
  assign t[38] = t[51] ^ x[42];
  assign t[39] = t[52] ^ x[43];
  assign t[3] = ~x[2] & t[30];
  assign t[40] = t[53] ^ x[44];
  assign t[41] = t[54] ^ x[45];
  assign t[42] = t[55] ^ x[46];
  assign t[43] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[44] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[45] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[46] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[47] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[48] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[49] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[4] = t[6];
  assign t[50] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[51] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[52] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[53] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[54] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[55] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = x[2] ? x[12] : t[10];
  assign t[8] = x[2] ? x[13] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind135(x, y);
 input [46:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[13];
  assign t[36] = t[49] ^ x[21];
  assign t[37] = t[50] ^ x[29];
  assign t[38] = t[51] ^ x[37];
  assign t[39] = t[52] ^ x[38];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[39];
  assign t[41] = t[54] ^ x[40];
  assign t[42] = t[55] ^ x[41];
  assign t[43] = t[56] ^ x[42];
  assign t[44] = t[57] ^ x[43];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = t[59] ^ x[45];
  assign t[47] = t[60] ^ x[46];
  assign t[48] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[49] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[51] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[52] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[53] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[54] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[55] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[56] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[57] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[58] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[59] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind136(x, y);
 input [43:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[22];
  assign t[32] = t[42] ^ x[30];
  assign t[33] = t[43] ^ x[31];
  assign t[34] = t[44] ^ x[39];
  assign t[35] = t[45] ^ x[40];
  assign t[36] = t[46] ^ x[41];
  assign t[37] = t[47] ^ x[42];
  assign t[38] = t[48] ^ x[43];
  assign t[39] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[41] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[42] = (x[23] & x[25] & ~x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[26] & ~x[28] & x[29]) | (x[23] & ~x[26] & x[27] & ~x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[24] & x[25] & ~x[26] & x[29]) | (x[24] & x[27] & ~x[28] & x[29]) | (x[25] & x[27] & x[29]);
  assign t[43] = (x[23] & x[24] & x[25] & ~x[28] & ~x[29]) | (x[23] & x[24] & x[26] & ~x[27] & ~x[29]) | (x[23] & x[25] & x[26] & ~x[28] & ~x[29]) | (~x[24] & x[25] & x[26] & x[27] & ~x[29]) | (x[24] & x[25] & x[26] & ~x[28]) | (x[24] & x[26] & x[27] & ~x[28]) | (x[23] & x[25] & ~x[27] & x[28]);
  assign t[44] = (x[32] & x[34] & ~x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[35] & ~x[37] & x[38]) | (x[32] & ~x[35] & x[36] & ~x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[33] & x[34] & ~x[35] & x[38]) | (x[33] & x[36] & ~x[37] & x[38]) | (x[34] & x[36] & x[38]);
  assign t[45] = (x[32] & x[33] & x[34] & ~x[37] & ~x[38]) | (x[32] & x[33] & x[35] & ~x[36] & ~x[38]) | (x[32] & x[34] & x[35] & ~x[37] & ~x[38]) | (~x[33] & x[34] & x[35] & x[36] & ~x[38]) | (x[33] & x[34] & x[35] & ~x[37]) | (x[33] & x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[36] & x[37]);
  assign t[46] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[47] = (x[24] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[24] & ~x[25] & x[26] & ~x[27] & x[29]) | (x[24] & ~x[25] & ~x[27] & x[28] & x[29]) | (x[23] & x[25] & x[26] & x[27] & x[28]) | (x[23] & ~x[25] & x[26] & x[29]) | (x[23] & ~x[27] & x[28] & x[29]) | (x[26] & x[28] & x[29]);
  assign t[48] = (x[33] & ~x[34] & x[35] & ~x[36] & x[37]) | (x[33] & ~x[34] & x[35] & ~x[36] & x[38]) | (x[33] & ~x[34] & ~x[36] & x[37] & x[38]) | (x[32] & x[34] & x[35] & x[36] & x[37]) | (x[32] & ~x[34] & x[35] & x[38]) | (x[32] & ~x[36] & x[37] & x[38]) | (x[35] & x[37] & x[38]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind137(x, y);
 input [46:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = ~(t[20] & t[34]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = ~(t[23] & t[35]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26] & t[36]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] & t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] & t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[38] & t[37]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[45]);
  assign t[33] = t[46] ^ x[10];
  assign t[34] = t[47] ^ x[21];
  assign t[35] = t[48] ^ x[29];
  assign t[36] = t[49] ^ x[37];
  assign t[37] = t[50] ^ x[38];
  assign t[38] = t[51] ^ x[39];
  assign t[39] = t[52] ^ x[40];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[41];
  assign t[41] = t[54] ^ x[42];
  assign t[42] = t[55] ^ x[43];
  assign t[43] = t[56] ^ x[44];
  assign t[44] = t[57] ^ x[45];
  assign t[45] = t[58] ^ x[46];
  assign t[46] = (x[3] & x[4] & x[5] & ~x[8] & ~x[9]) | (x[3] & x[4] & x[6] & ~x[7] & ~x[9]) | (x[3] & x[5] & x[6] & ~x[8] & ~x[9]) | (~x[4] & x[5] & x[6] & x[7] & ~x[9]) | (x[4] & x[5] & x[6] & ~x[8]) | (x[4] & x[6] & x[7] & ~x[8]) | (x[3] & x[5] & ~x[7] & x[8]);
  assign t[47] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[48] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[49] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[4] = t[6];
  assign t[50] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[51] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[52] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[53] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[54] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[55] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[56] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[57] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[58] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[11] : t[9];
  assign t[7] = x[2] ? x[12] : t[10];
  assign t[8] = x[2] ? x[13] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind138(x, y);
 input [46:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[13];
  assign t[33] = t[46] ^ x[21];
  assign t[34] = t[47] ^ x[29];
  assign t[35] = t[48] ^ x[37];
  assign t[36] = t[49] ^ x[38];
  assign t[37] = t[50] ^ x[39];
  assign t[38] = t[51] ^ x[40];
  assign t[39] = t[52] ^ x[41];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[42];
  assign t[41] = t[54] ^ x[43];
  assign t[42] = t[55] ^ x[44];
  assign t[43] = t[56] ^ x[45];
  assign t[44] = t[57] ^ x[46];
  assign t[45] = (x[6] & x[7] & x[8] & ~x[11] & ~x[12]) | (x[6] & x[7] & x[9] & ~x[10] & ~x[12]) | (x[6] & x[8] & x[9] & ~x[11] & ~x[12]) | (~x[7] & x[8] & x[9] & x[10] & ~x[12]) | (x[7] & x[8] & x[9] & ~x[11]) | (x[7] & x[9] & x[10] & ~x[11]) | (x[6] & x[8] & ~x[10] & x[11]);
  assign t[46] = (x[14] & x[15] & ~x[17] & x[18] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[14] & x[15] & ~x[16] & x[19] & ~x[20]) | (x[14] & ~x[17] & x[18] & x[19] & ~x[20]) | (x[14] & ~x[16] & x[17] & x[18]) | (x[15] & x[16] & ~x[17] & x[19]) | (x[15] & ~x[17] & x[18] & x[19]);
  assign t[47] = (x[22] & x[23] & ~x[25] & x[26] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[22] & x[23] & ~x[24] & x[27] & ~x[28]) | (x[22] & ~x[25] & x[26] & x[27] & ~x[28]) | (x[22] & ~x[24] & x[25] & x[26]) | (x[23] & x[24] & ~x[25] & x[27]) | (x[23] & ~x[25] & x[26] & x[27]);
  assign t[48] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[49] = (x[15] & ~x[16] & x[17] & ~x[18] & x[19]) | (x[15] & ~x[16] & x[17] & ~x[18] & x[20]) | (x[15] & ~x[16] & ~x[18] & x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[14] & ~x[16] & x[17] & x[20]) | (x[14] & ~x[18] & x[19] & x[20]) | (x[17] & x[19] & x[20]);
  assign t[4] = t[7];
  assign t[50] = (x[14] & x[15] & x[16] & ~x[19] & ~x[20]) | (x[14] & x[15] & x[17] & ~x[18] & ~x[20]) | (x[14] & x[16] & x[17] & ~x[19] & ~x[20]) | (~x[15] & x[16] & x[17] & x[18] & ~x[20]) | (x[15] & x[16] & x[17] & ~x[19]) | (x[15] & x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[18] & x[19]);
  assign t[51] = (x[23] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[23] & ~x[24] & x[25] & ~x[26] & x[28]) | (x[23] & ~x[24] & ~x[26] & x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[22] & ~x[24] & x[25] & x[28]) | (x[22] & ~x[26] & x[27] & x[28]) | (x[25] & x[27] & x[28]);
  assign t[52] = (x[22] & x[23] & x[24] & ~x[27] & ~x[28]) | (x[22] & x[23] & x[25] & ~x[26] & ~x[28]) | (x[22] & x[24] & x[25] & ~x[27] & ~x[28]) | (~x[23] & x[24] & x[25] & x[26] & ~x[28]) | (x[23] & x[24] & x[25] & ~x[27]) | (x[23] & x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[26] & x[27]);
  assign t[53] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[54] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[55] = (x[14] & x[16] & ~x[17] & x[18] & ~x[19]) | (x[14] & x[16] & ~x[17] & ~x[19] & x[20]) | (x[14] & ~x[17] & x[18] & ~x[19] & x[20]) | (x[14] & x[16] & x[17] & x[18] & x[19]) | (x[15] & x[16] & ~x[17] & x[20]) | (x[15] & x[18] & ~x[19] & x[20]) | (x[16] & x[18] & x[20]);
  assign t[56] = (x[22] & x[24] & ~x[25] & x[26] & ~x[27]) | (x[22] & x[24] & ~x[25] & ~x[27] & x[28]) | (x[22] & ~x[25] & x[26] & ~x[27] & x[28]) | (x[22] & x[24] & x[25] & x[26] & x[27]) | (x[23] & x[24] & ~x[25] & x[28]) | (x[23] & x[26] & ~x[27] & x[28]) | (x[24] & x[26] & x[28]);
  assign t[57] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1_ind(x, y);
 input [448:0] x;
 output [138:0] y;

  R1ind0 R1ind0_inst(.x({x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[17], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[28], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[29], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[39], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[40], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[50], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[51], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[61], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[72], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[73], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[84], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[94], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[95], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[105], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[106], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[116], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[117], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[127], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[128], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[138], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[139], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[150], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[161], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[172], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[183], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[184]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[184]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[184]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[184]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[184]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[184]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[184]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[180], x[183], x[182], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[259], x[184], x[258], x[257]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[183], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[180], x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[262], x[184], x[261], x[260]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[182], x[180], x[183], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[265], x[184], x[264], x[263]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[182], x[180], x[183], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[268], x[184], x[267], x[266]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[147], x[150], x[149], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[271], x[184], x[270], x[269]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[150], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[147], x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[274], x[184], x[273], x[272]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[149], x[147], x[150], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[277], x[184], x[276], x[275]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[149], x[147], x[150], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[280], x[184], x[279], x[278]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[158], x[161], x[160], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[283], x[184], x[282], x[281]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[161], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[158], x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[286], x[184], x[285], x[284]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[160], x[158], x[161], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[289], x[184], x[288], x[287]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[160], x[158], x[161], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[292], x[184], x[291], x[290]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[169], x[172], x[171], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[295], x[184], x[294], x[293]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[172], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[169], x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[298], x[184], x[297], x[296]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[171], x[169], x[172], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[301], x[184], x[300], x[299]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[171], x[169], x[172], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[304], x[184], x[303], x[302]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[103], x[106], x[105], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[307], x[184], x[306], x[305]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[106], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[103], x[105], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[310], x[184], x[309], x[308]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[105], x[103], x[106], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[313], x[184], x[312], x[311]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[105], x[103], x[106], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[316], x[184], x[315], x[314]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[136], x[139], x[138], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[319], x[184], x[318], x[317]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[139], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[136], x[138], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[322], x[184], x[321], x[320]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[138], x[136], x[139], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[325], x[184], x[324], x[323]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[138], x[136], x[139], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[328], x[184], x[327], x[326]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[125], x[128], x[127], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[331], x[184], x[330], x[329]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[128], x[125], x[127], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[334], x[184], x[333], x[332]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[127], x[125], x[128], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[337], x[184], x[336], x[335]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[127], x[125], x[128], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[340], x[184], x[339], x[338]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[114], x[117], x[116], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[343], x[184], x[342], x[341]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[117], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[114], x[116], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[346], x[184], x[345], x[344]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[116], x[114], x[117], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[349], x[184], x[348], x[347]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[116], x[114], x[117], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[352], x[184], x[351], x[350]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[59], x[180], x[62], x[61], x[183], x[182], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[355], x[259], x[184], x[354], x[353]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[62], x[183], x[59], x[61], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[180], x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[358], x[262], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[357], x[356]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[61], x[182], x[59], x[62], x[180], x[183], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[361], x[265], x[184], x[360], x[359]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[61], x[182], x[59], x[62], x[180], x[183], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[364], x[268], x[184], x[363], x[362]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[92], x[147], x[95], x[94], x[150], x[149], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[367], x[271], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[366], x[365]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[95], x[150], x[92], x[94], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[147], x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[370], x[274], x[184], x[369], x[368]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[94], x[149], x[92], x[95], x[147], x[150], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[373], x[277], x[184], x[372], x[371]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[94], x[149], x[92], x[95], x[147], x[150], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[376], x[280], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[375], x[374]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[81], x[158], x[84], x[83], x[161], x[160], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[379], x[283], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[184], x[378], x[377]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[84], x[161], x[81], x[83], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[158], x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[382], x[286], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[184], x[381], x[380]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[83], x[160], x[81], x[84], x[158], x[161], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[385], x[289], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[184], x[384], x[383]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[83], x[160], x[81], x[84], x[158], x[161], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[388], x[292], x[184], x[387], x[386]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[70], x[169], x[73], x[72], x[172], x[171], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[391], x[295], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[184], x[390], x[389]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[73], x[172], x[70], x[72], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[169], x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[394], x[298], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[184], x[393], x[392]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[72], x[171], x[70], x[73], x[169], x[172], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[397], x[301], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[184], x[396], x[395]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[72], x[171], x[70], x[73], x[169], x[172], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[400], x[304], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[399], x[398]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[180], x[103], x[26], x[183], x[182], x[106], x[105], x[29], x[28], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[259], x[307], x[403], x[184], x[402], x[401]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[183], x[106], x[29], x[180], x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[103], x[105], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[26], x[28], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[262], x[310], x[406], x[184], x[405], x[404]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[182], x[105], x[28], x[180], x[183], x[103], x[106], x[26], x[29], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[265], x[313], x[409], x[184], x[408], x[407]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[182], x[105], x[28], x[180], x[183], x[103], x[106], x[26], x[29], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[268], x[316], x[412], x[184], x[411], x[410]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[147], x[136], x[37], x[150], x[149], x[139], x[138], x[40], x[39], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[271], x[319], x[415], x[184], x[414], x[413]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[150], x[139], x[40], x[147], x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[136], x[138], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[37], x[39], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[274], x[322], x[418], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[417], x[416]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[149], x[138], x[39], x[147], x[150], x[136], x[139], x[37], x[40], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[277], x[325], x[421], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[420], x[419]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[149], x[138], x[39], x[147], x[150], x[136], x[139], x[37], x[40], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[280], x[328], x[424], x[184], x[423], x[422]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[158], x[125], x[48], x[161], x[160], x[128], x[127], x[51], x[50], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[283], x[331], x[427], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[426], x[425]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[161], x[128], x[51], x[158], x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[125], x[127], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[48], x[50], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[286], x[334], x[430], x[184], x[429], x[428]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[160], x[127], x[50], x[158], x[161], x[125], x[128], x[48], x[51], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[289], x[337], x[433], x[184], x[432], x[431]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[160], x[127], x[50], x[158], x[161], x[125], x[128], x[48], x[51], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[292], x[340], x[436], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[435], x[434]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[169], x[114], x[15], x[172], x[171], x[117], x[116], x[18], x[17], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[295], x[343], x[439], x[184], x[438], x[437]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[172], x[117], x[18], x[169], x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[114], x[116], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[15], x[17], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[298], x[346], x[442], x[184], x[441], x[440]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[171], x[116], x[17], x[169], x[172], x[114], x[117], x[15], x[18], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[301], x[349], x[445], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[184], x[444], x[443]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[171], x[116], x[17], x[169], x[172], x[114], x[117], x[15], x[18], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[304], x[352], x[448], x[184], x[447], x[446]}), .y(y[138]));
endmodule

module R2ind0(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[4] & ~t[5] & ~t[6] & ~t[7]) | (t[2] & ~t[3] & ~t[5] & ~t[6] & ~t[8]) | (t[2] & ~t[3] & ~t[4] & ~t[7] & ~t[8]) | (~t[2] & t[3] & t[4] & t[5] & ~t[8]) | (~t[2] & t[3] & t[6] & t[7] & ~t[8]) | (t[2] & ~t[4] & ~t[6] & t[8]) | (~t[2] & t[4] & t[6] & t[8]);
  assign t[2] = t[9] ^ x[7];
  assign t[3] = t[10] ^ x[1];
  assign t[4] = t[11] ^ x[2];
  assign t[5] = t[12] ^ x[3];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[3] & ~t[4] & ~t[5] & ~t[6] & ~t[7]) | (~t[2] & t[3] & ~t[5] & ~t[6] & ~t[8]) | (~t[2] & t[3] & ~t[4] & ~t[7] & ~t[8]) | (t[2] & ~t[3] & t[4] & t[5] & ~t[8]) | (t[2] & ~t[3] & t[6] & t[7] & ~t[8]) | (t[3] & ~t[5] & ~t[7] & t[8]) | (~t[3] & t[5] & t[7] & t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[7];
  assign t[4] = t[11] ^ x[2];
  assign t[5] = t[12] ^ x[3];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & ~t[4] & t[5] & ~t[6] & ~t[8]) | (t[2] & ~t[4] & ~t[5] & t[6] & ~t[7] & t[8]) | (~t[3] & t[4] & ~t[5] & ~t[6] & ~t[8]) | (~t[2] & t[4] & ~t[5] & ~t[6] & ~t[7]) | (~t[2] & ~t[3] & t[4] & ~t[7] & ~t[8]) | (~t[2] & t[4] & t[5] & ~t[6] & t[7]) | (t[4] & ~t[5] & t[7] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[7];
  assign t[5] = t[12] ^ x[3];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & t[4] & ~t[5] & ~t[7] & ~t[8]) | (t[3] & ~t[4] & ~t[5] & ~t[6] & t[7] & t[8]) | (~t[3] & ~t[4] & t[5] & ~t[6] & ~t[7]) | (~t[2] & ~t[4] & t[5] & ~t[7] & ~t[8]) | (~t[2] & ~t[3] & t[5] & ~t[6] & ~t[8]) | (~t[3] & t[4] & t[5] & t[6] & ~t[7]) | (~t[4] & t[5] & t[6] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[7];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & ~t[4] & ~t[6] & t[7] & ~t[8]) | (t[2] & t[4] & ~t[5] & ~t[6] & ~t[7] & t[8]) | (~t[3] & ~t[4] & t[6] & ~t[7] & ~t[8]) | (~t[2] & ~t[4] & ~t[5] & t[6] & ~t[7]) | (~t[2] & ~t[3] & ~t[5] & t[6] & ~t[8]) | (~t[2] & ~t[4] & t[5] & t[6] & t[7]) | (t[5] & t[6] & ~t[7] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[4];
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & ~t[5] & t[6] & ~t[7] & ~t[8]) | (t[3] & ~t[4] & t[5] & ~t[6] & ~t[7] & t[8]) | (~t[3] & ~t[4] & ~t[5] & ~t[6] & t[7]) | (~t[2] & ~t[5] & ~t[6] & t[7] & ~t[8]) | (~t[2] & ~t[3] & ~t[4] & t[7] & ~t[8]) | (~t[3] & t[4] & ~t[5] & t[6] & t[7]) | (t[4] & ~t[6] & t[7] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[4];
  assign t[6] = t[13] ^ x[5];
  assign t[7] = t[14] ^ x[7];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind6(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[4] & ~t[5] & t[6] & ~t[7] & ~t[8]) | (t[3] & ~t[4] & t[5] & ~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[5] & ~t[6] & ~t[7] & t[8]) | (~t[2] & ~t[3] & ~t[6] & ~t[7] & t[8]) | (~t[2] & ~t[3] & ~t[4] & ~t[5] & t[8]) | (t[2] & t[3] & ~t[6] & ~t[7] & t[8]) | (t[2] & t[3] & ~t[4] & ~t[5] & t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[4];
  assign t[6] = t[13] ^ x[5];
  assign t[7] = t[14] ^ x[6];
  assign t[8] = t[15] ^ x[7];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind7(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = t[1] & t[2];
  assign t[100] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[105] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[106] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[107] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[112] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[113] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[114] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[115] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[119] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[11] = ~x[0] & t[18];
  assign t[120] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[121] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[124] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[125] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[126] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[127] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[128] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~x[0] & t[19];
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[133] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[134] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[135] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[136] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[137] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[138] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[139] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[13] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[140] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[141] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[142] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[15] = (t[24] & ~t[25]) | (~t[24] & t[25]);
  assign t[16] = (t[26] & ~t[27]) | (~t[26] & t[27]);
  assign t[17] = (t[28] & ~t[29]) | (~t[28] & t[29]);
  assign t[18] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[19] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[34] ^ x[7];
  assign t[21] = t[35] ^ x[8];
  assign t[22] = t[36] ^ x[15];
  assign t[23] = t[37] ^ x[16];
  assign t[24] = t[38] ^ x[23];
  assign t[25] = t[39] ^ x[24];
  assign t[26] = t[40] ^ x[31];
  assign t[27] = t[41] ^ x[32];
  assign t[28] = t[42] ^ x[39];
  assign t[29] = t[43] ^ x[40];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = t[44] ^ x[47];
  assign t[31] = t[45] ^ x[48];
  assign t[32] = t[46] ^ x[55];
  assign t[33] = t[47] ^ x[56];
  assign t[34] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[35] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[36] = (t[55] & ~t[57] & ~t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[58] & ~t[59] & ~t[61]) | (t[55] & ~t[56] & ~t[57] & ~t[60] & ~t[61]) | (~t[55] & t[56] & t[57] & t[58] & ~t[61]) | (~t[55] & t[56] & t[59] & t[60] & ~t[61]) | (t[55] & ~t[57] & ~t[59] & t[61]) | (~t[55] & t[57] & t[59] & t[61]);
  assign t[37] = (t[55] & t[56] & ~t[57] & ~t[59] & t[60] & ~t[61]) | (t[55] & t[57] & ~t[58] & ~t[59] & ~t[60] & t[61]) | (~t[56] & ~t[57] & t[59] & ~t[60] & ~t[61]) | (~t[55] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[55] & ~t[56] & ~t[58] & t[59] & ~t[61]) | (~t[55] & ~t[57] & t[58] & t[59] & t[60]) | (t[58] & t[59] & ~t[60] & ~t[61]);
  assign t[38] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[39] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[41] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[42] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[43] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[44] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[45] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[46] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[47] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[48] = t[97] ^ x[7];
  assign t[49] = t[98] ^ x[2];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[99] ^ x[3];
  assign t[51] = t[100] ^ x[4];
  assign t[52] = t[101] ^ x[8];
  assign t[53] = t[102] ^ x[5];
  assign t[54] = t[103] ^ x[6];
  assign t[55] = t[104] ^ x[15];
  assign t[56] = t[105] ^ x[10];
  assign t[57] = t[106] ^ x[11];
  assign t[58] = t[107] ^ x[12];
  assign t[59] = t[108] ^ x[16];
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = t[109] ^ x[13];
  assign t[61] = t[110] ^ x[14];
  assign t[62] = t[111] ^ x[23];
  assign t[63] = t[112] ^ x[18];
  assign t[64] = t[113] ^ x[19];
  assign t[65] = t[114] ^ x[20];
  assign t[66] = t[115] ^ x[24];
  assign t[67] = t[116] ^ x[21];
  assign t[68] = t[117] ^ x[22];
  assign t[69] = t[118] ^ x[31];
  assign t[6] = ~x[0] & t[15];
  assign t[70] = t[119] ^ x[26];
  assign t[71] = t[120] ^ x[27];
  assign t[72] = t[121] ^ x[28];
  assign t[73] = t[122] ^ x[32];
  assign t[74] = t[123] ^ x[29];
  assign t[75] = t[124] ^ x[30];
  assign t[76] = t[125] ^ x[39];
  assign t[77] = t[126] ^ x[34];
  assign t[78] = t[127] ^ x[35];
  assign t[79] = t[128] ^ x[36];
  assign t[7] = ~(t[9] | t[10]);
  assign t[80] = t[129] ^ x[40];
  assign t[81] = t[130] ^ x[37];
  assign t[82] = t[131] ^ x[38];
  assign t[83] = t[132] ^ x[47];
  assign t[84] = t[133] ^ x[42];
  assign t[85] = t[134] ^ x[43];
  assign t[86] = t[135] ^ x[44];
  assign t[87] = t[136] ^ x[48];
  assign t[88] = t[137] ^ x[45];
  assign t[89] = t[138] ^ x[46];
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = t[139] ^ x[55];
  assign t[91] = t[140] ^ x[50];
  assign t[92] = t[141] ^ x[51];
  assign t[93] = t[142] ^ x[52];
  assign t[94] = t[143] ^ x[56];
  assign t[95] = t[144] ^ x[53];
  assign t[96] = t[145] ^ x[54];
  assign t[97] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[98] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[99] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind8(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = t[1] & t[2];
  assign t[100] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[105] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[106] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[107] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[112] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[113] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[114] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[115] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[119] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[11] = ~x[0] & t[18];
  assign t[120] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[121] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[124] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[125] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[126] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[127] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[128] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~x[0] & t[19];
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[133] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[134] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[135] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[136] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[137] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[138] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[139] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[13] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[140] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[141] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[142] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[15] = (t[24] & ~t[25]) | (~t[24] & t[25]);
  assign t[16] = (t[26] & ~t[27]) | (~t[26] & t[27]);
  assign t[17] = (t[28] & ~t[29]) | (~t[28] & t[29]);
  assign t[18] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[19] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[34] ^ x[7];
  assign t[21] = t[35] ^ x[8];
  assign t[22] = t[36] ^ x[15];
  assign t[23] = t[37] ^ x[16];
  assign t[24] = t[38] ^ x[23];
  assign t[25] = t[39] ^ x[24];
  assign t[26] = t[40] ^ x[31];
  assign t[27] = t[41] ^ x[32];
  assign t[28] = t[42] ^ x[39];
  assign t[29] = t[43] ^ x[40];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = t[44] ^ x[47];
  assign t[31] = t[45] ^ x[48];
  assign t[32] = t[46] ^ x[55];
  assign t[33] = t[47] ^ x[56];
  assign t[34] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[35] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[36] = (t[55] & ~t[57] & ~t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[58] & ~t[59] & ~t[61]) | (t[55] & ~t[56] & ~t[57] & ~t[60] & ~t[61]) | (~t[55] & t[56] & t[57] & t[58] & ~t[61]) | (~t[55] & t[56] & t[59] & t[60] & ~t[61]) | (t[55] & ~t[57] & ~t[59] & t[61]) | (~t[55] & t[57] & t[59] & t[61]);
  assign t[37] = (t[55] & t[56] & ~t[57] & ~t[59] & t[60] & ~t[61]) | (t[55] & t[57] & ~t[58] & ~t[59] & ~t[60] & t[61]) | (~t[56] & ~t[57] & t[59] & ~t[60] & ~t[61]) | (~t[55] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[55] & ~t[56] & ~t[58] & t[59] & ~t[61]) | (~t[55] & ~t[57] & t[58] & t[59] & t[60]) | (t[58] & t[59] & ~t[60] & ~t[61]);
  assign t[38] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[39] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[41] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[42] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[43] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[44] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[45] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[46] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[47] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[48] = t[97] ^ x[7];
  assign t[49] = t[98] ^ x[2];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[99] ^ x[3];
  assign t[51] = t[100] ^ x[4];
  assign t[52] = t[101] ^ x[8];
  assign t[53] = t[102] ^ x[5];
  assign t[54] = t[103] ^ x[6];
  assign t[55] = t[104] ^ x[15];
  assign t[56] = t[105] ^ x[10];
  assign t[57] = t[106] ^ x[11];
  assign t[58] = t[107] ^ x[12];
  assign t[59] = t[108] ^ x[16];
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = t[109] ^ x[13];
  assign t[61] = t[110] ^ x[14];
  assign t[62] = t[111] ^ x[23];
  assign t[63] = t[112] ^ x[18];
  assign t[64] = t[113] ^ x[19];
  assign t[65] = t[114] ^ x[20];
  assign t[66] = t[115] ^ x[24];
  assign t[67] = t[116] ^ x[21];
  assign t[68] = t[117] ^ x[22];
  assign t[69] = t[118] ^ x[31];
  assign t[6] = ~x[0] & t[15];
  assign t[70] = t[119] ^ x[26];
  assign t[71] = t[120] ^ x[27];
  assign t[72] = t[121] ^ x[28];
  assign t[73] = t[122] ^ x[32];
  assign t[74] = t[123] ^ x[29];
  assign t[75] = t[124] ^ x[30];
  assign t[76] = t[125] ^ x[39];
  assign t[77] = t[126] ^ x[34];
  assign t[78] = t[127] ^ x[35];
  assign t[79] = t[128] ^ x[36];
  assign t[7] = ~(t[9] | t[10]);
  assign t[80] = t[129] ^ x[40];
  assign t[81] = t[130] ^ x[37];
  assign t[82] = t[131] ^ x[38];
  assign t[83] = t[132] ^ x[47];
  assign t[84] = t[133] ^ x[42];
  assign t[85] = t[134] ^ x[43];
  assign t[86] = t[135] ^ x[44];
  assign t[87] = t[136] ^ x[48];
  assign t[88] = t[137] ^ x[45];
  assign t[89] = t[138] ^ x[46];
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = t[139] ^ x[55];
  assign t[91] = t[140] ^ x[50];
  assign t[92] = t[141] ^ x[51];
  assign t[93] = t[142] ^ x[52];
  assign t[94] = t[143] ^ x[56];
  assign t[95] = t[144] ^ x[53];
  assign t[96] = t[145] ^ x[54];
  assign t[97] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[98] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[99] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind9(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = t[1] & t[2];
  assign t[100] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[105] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[106] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[107] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[112] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[113] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[114] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[115] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[119] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[11] = ~x[0] & t[18];
  assign t[120] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[121] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[124] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[125] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[126] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[127] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[128] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~x[0] & t[19];
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[133] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[134] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[135] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[136] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[137] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[138] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[139] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[13] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[140] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[141] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[142] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[15] = (t[24] & ~t[25]) | (~t[24] & t[25]);
  assign t[16] = (t[26] & ~t[27]) | (~t[26] & t[27]);
  assign t[17] = (t[28] & ~t[29]) | (~t[28] & t[29]);
  assign t[18] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[19] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[34] ^ x[7];
  assign t[21] = t[35] ^ x[8];
  assign t[22] = t[36] ^ x[15];
  assign t[23] = t[37] ^ x[16];
  assign t[24] = t[38] ^ x[23];
  assign t[25] = t[39] ^ x[24];
  assign t[26] = t[40] ^ x[31];
  assign t[27] = t[41] ^ x[32];
  assign t[28] = t[42] ^ x[39];
  assign t[29] = t[43] ^ x[40];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = t[44] ^ x[47];
  assign t[31] = t[45] ^ x[48];
  assign t[32] = t[46] ^ x[55];
  assign t[33] = t[47] ^ x[56];
  assign t[34] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[35] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[36] = (t[55] & ~t[57] & ~t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[58] & ~t[59] & ~t[61]) | (t[55] & ~t[56] & ~t[57] & ~t[60] & ~t[61]) | (~t[55] & t[56] & t[57] & t[58] & ~t[61]) | (~t[55] & t[56] & t[59] & t[60] & ~t[61]) | (t[55] & ~t[57] & ~t[59] & t[61]) | (~t[55] & t[57] & t[59] & t[61]);
  assign t[37] = (t[55] & t[56] & ~t[57] & ~t[59] & t[60] & ~t[61]) | (t[55] & t[57] & ~t[58] & ~t[59] & ~t[60] & t[61]) | (~t[56] & ~t[57] & t[59] & ~t[60] & ~t[61]) | (~t[55] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[55] & ~t[56] & ~t[58] & t[59] & ~t[61]) | (~t[55] & ~t[57] & t[58] & t[59] & t[60]) | (t[58] & t[59] & ~t[60] & ~t[61]);
  assign t[38] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[39] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[41] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[42] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[43] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[44] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[45] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[46] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[47] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[48] = t[97] ^ x[7];
  assign t[49] = t[98] ^ x[2];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[99] ^ x[3];
  assign t[51] = t[100] ^ x[4];
  assign t[52] = t[101] ^ x[8];
  assign t[53] = t[102] ^ x[5];
  assign t[54] = t[103] ^ x[6];
  assign t[55] = t[104] ^ x[15];
  assign t[56] = t[105] ^ x[10];
  assign t[57] = t[106] ^ x[11];
  assign t[58] = t[107] ^ x[12];
  assign t[59] = t[108] ^ x[16];
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = t[109] ^ x[13];
  assign t[61] = t[110] ^ x[14];
  assign t[62] = t[111] ^ x[23];
  assign t[63] = t[112] ^ x[18];
  assign t[64] = t[113] ^ x[19];
  assign t[65] = t[114] ^ x[20];
  assign t[66] = t[115] ^ x[24];
  assign t[67] = t[116] ^ x[21];
  assign t[68] = t[117] ^ x[22];
  assign t[69] = t[118] ^ x[31];
  assign t[6] = ~x[0] & t[15];
  assign t[70] = t[119] ^ x[26];
  assign t[71] = t[120] ^ x[27];
  assign t[72] = t[121] ^ x[28];
  assign t[73] = t[122] ^ x[32];
  assign t[74] = t[123] ^ x[29];
  assign t[75] = t[124] ^ x[30];
  assign t[76] = t[125] ^ x[39];
  assign t[77] = t[126] ^ x[34];
  assign t[78] = t[127] ^ x[35];
  assign t[79] = t[128] ^ x[36];
  assign t[7] = ~(t[9] | t[10]);
  assign t[80] = t[129] ^ x[40];
  assign t[81] = t[130] ^ x[37];
  assign t[82] = t[131] ^ x[38];
  assign t[83] = t[132] ^ x[47];
  assign t[84] = t[133] ^ x[42];
  assign t[85] = t[134] ^ x[43];
  assign t[86] = t[135] ^ x[44];
  assign t[87] = t[136] ^ x[48];
  assign t[88] = t[137] ^ x[45];
  assign t[89] = t[138] ^ x[46];
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = t[139] ^ x[55];
  assign t[91] = t[140] ^ x[50];
  assign t[92] = t[141] ^ x[51];
  assign t[93] = t[142] ^ x[52];
  assign t[94] = t[143] ^ x[56];
  assign t[95] = t[144] ^ x[53];
  assign t[96] = t[145] ^ x[54];
  assign t[97] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[98] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[99] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind10(x, y);
 input [56:0] x;
 output y;

 wire [145:0] t;
  assign t[0] = t[1] & t[2];
  assign t[100] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[105] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[106] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[107] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[112] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[113] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[114] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[115] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[119] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[11] = ~x[0] & t[18];
  assign t[120] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[121] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[124] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[125] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[126] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[127] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[128] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~x[0] & t[19];
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[133] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[134] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[135] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[136] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[137] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[138] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[139] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[13] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[140] = (x[49] & ~1'b0 & ~1'b0) | (~x[49] & 1'b0 & ~1'b0) | (~x[49] & ~1'b0 & 1'b0) | (x[49] & 1'b0 & 1'b0);
  assign t[141] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[142] = (x[49] & ~1'b0) | (~x[49] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[15] = (t[24] & ~t[25]) | (~t[24] & t[25]);
  assign t[16] = (t[26] & ~t[27]) | (~t[26] & t[27]);
  assign t[17] = (t[28] & ~t[29]) | (~t[28] & t[29]);
  assign t[18] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[19] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[34] ^ x[7];
  assign t[21] = t[35] ^ x[8];
  assign t[22] = t[36] ^ x[15];
  assign t[23] = t[37] ^ x[16];
  assign t[24] = t[38] ^ x[23];
  assign t[25] = t[39] ^ x[24];
  assign t[26] = t[40] ^ x[31];
  assign t[27] = t[41] ^ x[32];
  assign t[28] = t[42] ^ x[39];
  assign t[29] = t[43] ^ x[40];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = t[44] ^ x[47];
  assign t[31] = t[45] ^ x[48];
  assign t[32] = t[46] ^ x[55];
  assign t[33] = t[47] ^ x[56];
  assign t[34] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[35] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[36] = (t[55] & ~t[57] & ~t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[58] & ~t[59] & ~t[61]) | (t[55] & ~t[56] & ~t[57] & ~t[60] & ~t[61]) | (~t[55] & t[56] & t[57] & t[58] & ~t[61]) | (~t[55] & t[56] & t[59] & t[60] & ~t[61]) | (t[55] & ~t[57] & ~t[59] & t[61]) | (~t[55] & t[57] & t[59] & t[61]);
  assign t[37] = (t[55] & t[56] & ~t[57] & ~t[59] & t[60] & ~t[61]) | (t[55] & t[57] & ~t[58] & ~t[59] & ~t[60] & t[61]) | (~t[56] & ~t[57] & t[59] & ~t[60] & ~t[61]) | (~t[55] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[55] & ~t[56] & ~t[58] & t[59] & ~t[61]) | (~t[55] & ~t[57] & t[58] & t[59] & t[60]) | (t[58] & t[59] & ~t[60] & ~t[61]);
  assign t[38] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[39] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[41] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[42] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[43] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[44] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[45] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[46] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[47] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[48] = t[97] ^ x[7];
  assign t[49] = t[98] ^ x[2];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[99] ^ x[3];
  assign t[51] = t[100] ^ x[4];
  assign t[52] = t[101] ^ x[8];
  assign t[53] = t[102] ^ x[5];
  assign t[54] = t[103] ^ x[6];
  assign t[55] = t[104] ^ x[15];
  assign t[56] = t[105] ^ x[10];
  assign t[57] = t[106] ^ x[11];
  assign t[58] = t[107] ^ x[12];
  assign t[59] = t[108] ^ x[16];
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = t[109] ^ x[13];
  assign t[61] = t[110] ^ x[14];
  assign t[62] = t[111] ^ x[23];
  assign t[63] = t[112] ^ x[18];
  assign t[64] = t[113] ^ x[19];
  assign t[65] = t[114] ^ x[20];
  assign t[66] = t[115] ^ x[24];
  assign t[67] = t[116] ^ x[21];
  assign t[68] = t[117] ^ x[22];
  assign t[69] = t[118] ^ x[31];
  assign t[6] = ~x[0] & t[15];
  assign t[70] = t[119] ^ x[26];
  assign t[71] = t[120] ^ x[27];
  assign t[72] = t[121] ^ x[28];
  assign t[73] = t[122] ^ x[32];
  assign t[74] = t[123] ^ x[29];
  assign t[75] = t[124] ^ x[30];
  assign t[76] = t[125] ^ x[39];
  assign t[77] = t[126] ^ x[34];
  assign t[78] = t[127] ^ x[35];
  assign t[79] = t[128] ^ x[36];
  assign t[7] = ~(t[9] | t[10]);
  assign t[80] = t[129] ^ x[40];
  assign t[81] = t[130] ^ x[37];
  assign t[82] = t[131] ^ x[38];
  assign t[83] = t[132] ^ x[47];
  assign t[84] = t[133] ^ x[42];
  assign t[85] = t[134] ^ x[43];
  assign t[86] = t[135] ^ x[44];
  assign t[87] = t[136] ^ x[48];
  assign t[88] = t[137] ^ x[45];
  assign t[89] = t[138] ^ x[46];
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = t[139] ^ x[55];
  assign t[91] = t[140] ^ x[50];
  assign t[92] = t[141] ^ x[51];
  assign t[93] = t[142] ^ x[52];
  assign t[94] = t[143] ^ x[56];
  assign t[95] = t[144] ^ x[53];
  assign t[96] = t[145] ^ x[54];
  assign t[97] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[98] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[99] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind14(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind15(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind16(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind17(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind19(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind20(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind21(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind22(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind23(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind24(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind25(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind28(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~x[0] & t[3];
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind29(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~x[0] & t[3];
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind30(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~x[0] & t[3];
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind31(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~x[0] & t[3];
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind34(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind35(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind36(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind37(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind38(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind39(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind40(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind41(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind42(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind43(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind44(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind45(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind46(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind47(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind48(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind49(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind50(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind51(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind52(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind53(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind54(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind55(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind56(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind57(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind58(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind59(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13] & t[14] & ~t[15] & ~t[17] & t[18] & ~t[19]) | (t[13] & t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[19]) | (~t[13] & ~t[15] & ~t[16] & t[17] & ~t[18]) | (~t[13] & ~t[14] & ~t[16] & t[17] & ~t[19]) | (~t[13] & ~t[15] & t[16] & t[17] & t[18]) | (t[16] & t[17] & ~t[18] & ~t[19]);
  assign t[11] = (t[20] & ~t[22] & ~t[23] & ~t[24] & ~t[25]) | (t[20] & ~t[21] & ~t[23] & ~t[24] & ~t[26]) | (t[20] & ~t[21] & ~t[22] & ~t[25] & ~t[26]) | (~t[20] & t[21] & t[22] & t[23] & ~t[26]) | (~t[20] & t[21] & t[24] & t[25] & ~t[26]) | (t[20] & ~t[22] & ~t[24] & t[26]) | (~t[20] & t[22] & t[24] & t[26]);
  assign t[12] = (t[20] & t[21] & ~t[22] & ~t[24] & t[25] & ~t[26]) | (t[20] & t[22] & ~t[23] & ~t[24] & ~t[25] & t[26]) | (~t[21] & ~t[22] & t[24] & ~t[25] & ~t[26]) | (~t[20] & ~t[22] & ~t[23] & t[24] & ~t[25]) | (~t[20] & ~t[21] & ~t[23] & t[24] & ~t[26]) | (~t[20] & ~t[22] & t[23] & t[24] & t[25]) | (t[23] & t[24] & ~t[25] & ~t[26]);
  assign t[13] = t[27] ^ x[7];
  assign t[14] = t[28] ^ x[2];
  assign t[15] = t[29] ^ x[3];
  assign t[16] = t[30] ^ x[4];
  assign t[17] = t[31] ^ x[8];
  assign t[18] = t[32] ^ x[5];
  assign t[19] = t[33] ^ x[6];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[20] = t[34] ^ x[15];
  assign t[21] = t[35] ^ x[10];
  assign t[22] = t[36] ^ x[11];
  assign t[23] = t[37] ^ x[12];
  assign t[24] = t[38] ^ x[16];
  assign t[25] = t[39] ^ x[13];
  assign t[26] = t[40] ^ x[14];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = (t[5] & ~t[6]) | (~t[5] & t[6]);
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[7] & ~t[8]) | (~t[7] & t[8]);
  assign t[5] = t[9] ^ x[7];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[15];
  assign t[8] = t[12] ^ x[16];
  assign t[9] = (t[13] & ~t[15] & ~t[16] & ~t[17] & ~t[18]) | (t[13] & ~t[14] & ~t[16] & ~t[17] & ~t[19]) | (t[13] & ~t[14] & ~t[15] & ~t[18] & ~t[19]) | (~t[13] & t[14] & t[15] & t[16] & ~t[19]) | (~t[13] & t[14] & t[17] & t[18] & ~t[19]) | (t[13] & ~t[15] & ~t[17] & t[19]) | (~t[13] & t[15] & t[17] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind60(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind61(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind62(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind63(x, y);
 input [8:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[17] ^ x[4];
  assign t[11] = t[18] ^ x[8];
  assign t[12] = t[19] ^ x[5];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = ~x[0] & t[2];
  assign t[20] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[2] = (t[3] & ~t[4]) | (~t[3] & t[4]);
  assign t[3] = t[5] ^ x[7];
  assign t[4] = t[6] ^ x[8];
  assign t[5] = (t[7] & ~t[9] & ~t[10] & ~t[11] & ~t[12]) | (t[7] & ~t[8] & ~t[10] & ~t[11] & ~t[13]) | (t[7] & ~t[8] & ~t[9] & ~t[12] & ~t[13]) | (~t[7] & t[8] & t[9] & t[10] & ~t[13]) | (~t[7] & t[8] & t[11] & t[12] & ~t[13]) | (t[7] & ~t[9] & ~t[11] & t[13]) | (~t[7] & t[9] & t[11] & t[13]);
  assign t[6] = (t[7] & t[8] & ~t[9] & ~t[11] & t[12] & ~t[13]) | (t[7] & t[9] & ~t[10] & ~t[11] & ~t[12] & t[13]) | (~t[8] & ~t[9] & t[11] & ~t[12] & ~t[13]) | (~t[7] & ~t[9] & ~t[10] & t[11] & ~t[12]) | (~t[7] & ~t[8] & ~t[10] & t[11] & ~t[13]) | (~t[7] & ~t[9] & t[10] & t[11] & t[12]) | (t[10] & t[11] & ~t[12] & ~t[13]);
  assign t[7] = t[14] ^ x[7];
  assign t[8] = t[15] ^ x[2];
  assign t[9] = t[16] ^ x[3];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind64(x, y);
 input [8:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[17] ^ x[4];
  assign t[11] = t[18] ^ x[8];
  assign t[12] = t[19] ^ x[5];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = ~x[0] & t[2];
  assign t[20] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[2] = (t[3] & ~t[4]) | (~t[3] & t[4]);
  assign t[3] = t[5] ^ x[7];
  assign t[4] = t[6] ^ x[8];
  assign t[5] = (t[7] & ~t[9] & ~t[10] & ~t[11] & ~t[12]) | (t[7] & ~t[8] & ~t[10] & ~t[11] & ~t[13]) | (t[7] & ~t[8] & ~t[9] & ~t[12] & ~t[13]) | (~t[7] & t[8] & t[9] & t[10] & ~t[13]) | (~t[7] & t[8] & t[11] & t[12] & ~t[13]) | (t[7] & ~t[9] & ~t[11] & t[13]) | (~t[7] & t[9] & t[11] & t[13]);
  assign t[6] = (t[7] & t[8] & ~t[9] & ~t[11] & t[12] & ~t[13]) | (t[7] & t[9] & ~t[10] & ~t[11] & ~t[12] & t[13]) | (~t[8] & ~t[9] & t[11] & ~t[12] & ~t[13]) | (~t[7] & ~t[9] & ~t[10] & t[11] & ~t[12]) | (~t[7] & ~t[8] & ~t[10] & t[11] & ~t[13]) | (~t[7] & ~t[9] & t[10] & t[11] & t[12]) | (t[10] & t[11] & ~t[12] & ~t[13]);
  assign t[7] = t[14] ^ x[7];
  assign t[8] = t[15] ^ x[2];
  assign t[9] = t[16] ^ x[3];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind65(x, y);
 input [8:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[17] ^ x[4];
  assign t[11] = t[18] ^ x[8];
  assign t[12] = t[19] ^ x[5];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = ~x[0] & t[2];
  assign t[20] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[2] = (t[3] & ~t[4]) | (~t[3] & t[4]);
  assign t[3] = t[5] ^ x[7];
  assign t[4] = t[6] ^ x[8];
  assign t[5] = (t[7] & ~t[9] & ~t[10] & ~t[11] & ~t[12]) | (t[7] & ~t[8] & ~t[10] & ~t[11] & ~t[13]) | (t[7] & ~t[8] & ~t[9] & ~t[12] & ~t[13]) | (~t[7] & t[8] & t[9] & t[10] & ~t[13]) | (~t[7] & t[8] & t[11] & t[12] & ~t[13]) | (t[7] & ~t[9] & ~t[11] & t[13]) | (~t[7] & t[9] & t[11] & t[13]);
  assign t[6] = (t[7] & t[8] & ~t[9] & ~t[11] & t[12] & ~t[13]) | (t[7] & t[9] & ~t[10] & ~t[11] & ~t[12] & t[13]) | (~t[8] & ~t[9] & t[11] & ~t[12] & ~t[13]) | (~t[7] & ~t[9] & ~t[10] & t[11] & ~t[12]) | (~t[7] & ~t[8] & ~t[10] & t[11] & ~t[13]) | (~t[7] & ~t[9] & t[10] & t[11] & t[12]) | (t[10] & t[11] & ~t[12] & ~t[13]);
  assign t[7] = t[14] ^ x[7];
  assign t[8] = t[15] ^ x[2];
  assign t[9] = t[16] ^ x[3];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind66(x, y);
 input [8:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[17] ^ x[4];
  assign t[11] = t[18] ^ x[8];
  assign t[12] = t[19] ^ x[5];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = ~x[0] & t[2];
  assign t[20] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[2] = (t[3] & ~t[4]) | (~t[3] & t[4]);
  assign t[3] = t[5] ^ x[7];
  assign t[4] = t[6] ^ x[8];
  assign t[5] = (t[7] & ~t[9] & ~t[10] & ~t[11] & ~t[12]) | (t[7] & ~t[8] & ~t[10] & ~t[11] & ~t[13]) | (t[7] & ~t[8] & ~t[9] & ~t[12] & ~t[13]) | (~t[7] & t[8] & t[9] & t[10] & ~t[13]) | (~t[7] & t[8] & t[11] & t[12] & ~t[13]) | (t[7] & ~t[9] & ~t[11] & t[13]) | (~t[7] & t[9] & t[11] & t[13]);
  assign t[6] = (t[7] & t[8] & ~t[9] & ~t[11] & t[12] & ~t[13]) | (t[7] & t[9] & ~t[10] & ~t[11] & ~t[12] & t[13]) | (~t[8] & ~t[9] & t[11] & ~t[12] & ~t[13]) | (~t[7] & ~t[9] & ~t[10] & t[11] & ~t[12]) | (~t[7] & ~t[8] & ~t[10] & t[11] & ~t[13]) | (~t[7] & ~t[9] & t[10] & t[11] & t[12]) | (t[10] & t[11] & ~t[12] & ~t[13]);
  assign t[7] = t[14] ^ x[7];
  assign t[8] = t[15] ^ x[2];
  assign t[9] = t[16] ^ x[3];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind67(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind68(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind69(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind70(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign t[11] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[12] = (t[21] & ~t[23] & ~t[24] & ~t[25] & ~t[26]) | (t[21] & ~t[22] & ~t[24] & ~t[25] & ~t[27]) | (t[21] & ~t[22] & ~t[23] & ~t[26] & ~t[27]) | (~t[21] & t[22] & t[23] & t[24] & ~t[27]) | (~t[21] & t[22] & t[25] & t[26] & ~t[27]) | (t[21] & ~t[23] & ~t[25] & t[27]) | (~t[21] & t[23] & t[25] & t[27]);
  assign t[13] = (t[21] & t[22] & ~t[23] & ~t[25] & t[26] & ~t[27]) | (t[21] & t[23] & ~t[24] & ~t[25] & ~t[26] & t[27]) | (~t[22] & ~t[23] & t[25] & ~t[26] & ~t[27]) | (~t[21] & ~t[23] & ~t[24] & t[25] & ~t[26]) | (~t[21] & ~t[22] & ~t[24] & t[25] & ~t[27]) | (~t[21] & ~t[23] & t[24] & t[25] & t[26]) | (t[24] & t[25] & ~t[26] & ~t[27]);
  assign t[14] = t[28] ^ x[7];
  assign t[15] = t[29] ^ x[2];
  assign t[16] = t[30] ^ x[3];
  assign t[17] = t[31] ^ x[4];
  assign t[18] = t[32] ^ x[8];
  assign t[19] = t[33] ^ x[5];
  assign t[1] = ~t[3];
  assign t[20] = t[34] ^ x[6];
  assign t[21] = t[35] ^ x[15];
  assign t[22] = t[36] ^ x[10];
  assign t[23] = t[37] ^ x[11];
  assign t[24] = t[38] ^ x[12];
  assign t[25] = t[39] ^ x[16];
  assign t[26] = t[40] ^ x[13];
  assign t[27] = t[41] ^ x[14];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = ~x[0] & t[5];
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[41] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[5] = (t[8] & ~t[9]) | (~t[8] & t[9]);
  assign t[6] = t[10] ^ x[7];
  assign t[7] = t[11] ^ x[8];
  assign t[8] = t[12] ^ x[15];
  assign t[9] = t[13] ^ x[16];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind71(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign t[11] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[12] = (t[21] & ~t[23] & ~t[24] & ~t[25] & ~t[26]) | (t[21] & ~t[22] & ~t[24] & ~t[25] & ~t[27]) | (t[21] & ~t[22] & ~t[23] & ~t[26] & ~t[27]) | (~t[21] & t[22] & t[23] & t[24] & ~t[27]) | (~t[21] & t[22] & t[25] & t[26] & ~t[27]) | (t[21] & ~t[23] & ~t[25] & t[27]) | (~t[21] & t[23] & t[25] & t[27]);
  assign t[13] = (t[21] & t[22] & ~t[23] & ~t[25] & t[26] & ~t[27]) | (t[21] & t[23] & ~t[24] & ~t[25] & ~t[26] & t[27]) | (~t[22] & ~t[23] & t[25] & ~t[26] & ~t[27]) | (~t[21] & ~t[23] & ~t[24] & t[25] & ~t[26]) | (~t[21] & ~t[22] & ~t[24] & t[25] & ~t[27]) | (~t[21] & ~t[23] & t[24] & t[25] & t[26]) | (t[24] & t[25] & ~t[26] & ~t[27]);
  assign t[14] = t[28] ^ x[7];
  assign t[15] = t[29] ^ x[2];
  assign t[16] = t[30] ^ x[3];
  assign t[17] = t[31] ^ x[4];
  assign t[18] = t[32] ^ x[8];
  assign t[19] = t[33] ^ x[5];
  assign t[1] = ~t[3];
  assign t[20] = t[34] ^ x[6];
  assign t[21] = t[35] ^ x[15];
  assign t[22] = t[36] ^ x[10];
  assign t[23] = t[37] ^ x[11];
  assign t[24] = t[38] ^ x[12];
  assign t[25] = t[39] ^ x[16];
  assign t[26] = t[40] ^ x[13];
  assign t[27] = t[41] ^ x[14];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = ~x[0] & t[5];
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[41] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[5] = (t[8] & ~t[9]) | (~t[8] & t[9]);
  assign t[6] = t[10] ^ x[7];
  assign t[7] = t[11] ^ x[8];
  assign t[8] = t[12] ^ x[15];
  assign t[9] = t[13] ^ x[16];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind72(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign t[11] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[12] = (t[21] & ~t[23] & ~t[24] & ~t[25] & ~t[26]) | (t[21] & ~t[22] & ~t[24] & ~t[25] & ~t[27]) | (t[21] & ~t[22] & ~t[23] & ~t[26] & ~t[27]) | (~t[21] & t[22] & t[23] & t[24] & ~t[27]) | (~t[21] & t[22] & t[25] & t[26] & ~t[27]) | (t[21] & ~t[23] & ~t[25] & t[27]) | (~t[21] & t[23] & t[25] & t[27]);
  assign t[13] = (t[21] & t[22] & ~t[23] & ~t[25] & t[26] & ~t[27]) | (t[21] & t[23] & ~t[24] & ~t[25] & ~t[26] & t[27]) | (~t[22] & ~t[23] & t[25] & ~t[26] & ~t[27]) | (~t[21] & ~t[23] & ~t[24] & t[25] & ~t[26]) | (~t[21] & ~t[22] & ~t[24] & t[25] & ~t[27]) | (~t[21] & ~t[23] & t[24] & t[25] & t[26]) | (t[24] & t[25] & ~t[26] & ~t[27]);
  assign t[14] = t[28] ^ x[7];
  assign t[15] = t[29] ^ x[2];
  assign t[16] = t[30] ^ x[3];
  assign t[17] = t[31] ^ x[4];
  assign t[18] = t[32] ^ x[8];
  assign t[19] = t[33] ^ x[5];
  assign t[1] = ~t[3];
  assign t[20] = t[34] ^ x[6];
  assign t[21] = t[35] ^ x[15];
  assign t[22] = t[36] ^ x[10];
  assign t[23] = t[37] ^ x[11];
  assign t[24] = t[38] ^ x[12];
  assign t[25] = t[39] ^ x[16];
  assign t[26] = t[40] ^ x[13];
  assign t[27] = t[41] ^ x[14];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = ~x[0] & t[5];
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[41] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[5] = (t[8] & ~t[9]) | (~t[8] & t[9]);
  assign t[6] = t[10] ^ x[7];
  assign t[7] = t[11] ^ x[8];
  assign t[8] = t[12] ^ x[15];
  assign t[9] = t[13] ^ x[16];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind73(x, y);
 input [16:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign t[11] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[12] = (t[21] & ~t[23] & ~t[24] & ~t[25] & ~t[26]) | (t[21] & ~t[22] & ~t[24] & ~t[25] & ~t[27]) | (t[21] & ~t[22] & ~t[23] & ~t[26] & ~t[27]) | (~t[21] & t[22] & t[23] & t[24] & ~t[27]) | (~t[21] & t[22] & t[25] & t[26] & ~t[27]) | (t[21] & ~t[23] & ~t[25] & t[27]) | (~t[21] & t[23] & t[25] & t[27]);
  assign t[13] = (t[21] & t[22] & ~t[23] & ~t[25] & t[26] & ~t[27]) | (t[21] & t[23] & ~t[24] & ~t[25] & ~t[26] & t[27]) | (~t[22] & ~t[23] & t[25] & ~t[26] & ~t[27]) | (~t[21] & ~t[23] & ~t[24] & t[25] & ~t[26]) | (~t[21] & ~t[22] & ~t[24] & t[25] & ~t[27]) | (~t[21] & ~t[23] & t[24] & t[25] & t[26]) | (t[24] & t[25] & ~t[26] & ~t[27]);
  assign t[14] = t[28] ^ x[7];
  assign t[15] = t[29] ^ x[2];
  assign t[16] = t[30] ^ x[3];
  assign t[17] = t[31] ^ x[4];
  assign t[18] = t[32] ^ x[8];
  assign t[19] = t[33] ^ x[5];
  assign t[1] = ~t[3];
  assign t[20] = t[34] ^ x[6];
  assign t[21] = t[35] ^ x[15];
  assign t[22] = t[36] ^ x[10];
  assign t[23] = t[37] ^ x[11];
  assign t[24] = t[38] ^ x[12];
  assign t[25] = t[39] ^ x[16];
  assign t[26] = t[40] ^ x[13];
  assign t[27] = t[41] ^ x[14];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[29] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[2] = ~x[0] & t[4];
  assign t[30] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[31] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[32] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[33] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[34] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[35] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[36] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[37] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[38] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[39] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[3] = ~x[0] & t[5];
  assign t[40] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[41] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[4] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[5] = (t[8] & ~t[9]) | (~t[8] & t[9]);
  assign t[6] = t[10] ^ x[7];
  assign t[7] = t[11] ^ x[8];
  assign t[8] = t[12] ^ x[15];
  assign t[9] = t[13] ^ x[16];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind74(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind75(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind76(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind77(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[36]);
  assign t[12] = ~(t[34] | t[35]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[17] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[18];
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[4]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[9]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[8]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[9] & t[11]);
  assign t[29] = ~(t[30] & t[33]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[8]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[39] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[39] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[39] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[39] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[39] & ~t[43]) | (~t[39] & t[43]);
  assign t[37] = t[45] ^ x[10];
  assign t[38] = t[46] ^ x[11];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[49] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[4] = ~x[2] & t[32];
  assign t[50] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[51] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[52] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[6];
  assign t[56] = t[70] ^ x[7];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[8];
  assign t[59] = t[73] ^ x[9];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[19];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[20];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[22];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[68] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[69] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[73] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[74] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[75] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[76] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[77] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[78] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[79] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[7] = ~(t[33] | t[10]);
  assign t[80] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[8] = ~(t[34]);
  assign t[9] = ~(t[35]);
  assign y = (t[0] & ~t[13] & ~t[23]) | (~t[0] & t[13] & ~t[23]) | (~t[0] & ~t[13] & t[23]) | (t[0] & t[13] & t[23]);
endmodule

module R2ind78(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[34]);
  assign t[12] = ~(t[32] | t[33]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[17] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[18];
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[4]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[9]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[8]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[17] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[9] & t[11]);
  assign t[29] = t[6] | t[31];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[37] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[37] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[37] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[37] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[37] & ~t[41]) | (~t[37] & t[41]);
  assign t[35] = t[43] ^ x[10];
  assign t[36] = t[44] ^ x[11];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[60] & ~t[61] & t[62] & ~t[63] & t[64]) | (~t[59] & t[60] & ~t[61] & ~t[62] & ~t[64]) | (~t[58] & t[60] & ~t[61] & ~t[62] & ~t[63]) | (~t[58] & ~t[59] & t[60] & ~t[63] & ~t[64]) | (~t[58] & t[60] & t[61] & ~t[62] & t[63]) | (t[60] & ~t[61] & t[63] & ~t[64]);
  assign t[47] = (t[59] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (~t[58] & t[59] & ~t[61] & ~t[62] & ~t[64]) | (~t[58] & t[59] & ~t[60] & ~t[63] & ~t[64]) | (t[58] & ~t[59] & t[60] & t[61] & ~t[64]) | (t[58] & ~t[59] & t[62] & t[63] & ~t[64]) | (t[59] & ~t[61] & ~t[63] & t[64]) | (~t[59] & t[61] & t[63] & t[64]);
  assign t[48] = (t[58] & t[59] & t[60] & ~t[61] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & ~t[61] & ~t[62] & t[63] & t[64]) | (~t[59] & ~t[60] & t[61] & ~t[62] & ~t[63]) | (~t[58] & ~t[60] & t[61] & ~t[63] & ~t[64]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[64]) | (~t[59] & t[60] & t[61] & t[62] & ~t[63]) | (~t[60] & t[61] & t[62] & ~t[64]);
  assign t[49] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[4] = ~x[2] & t[30];
  assign t[50] = (t[58] & t[59] & ~t[61] & t[62] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[61] & ~t[62] & t[63] & ~t[64]) | (~t[58] & ~t[59] & ~t[60] & t[63] & ~t[64]) | (~t[59] & t[60] & ~t[61] & t[62] & t[63]) | (t[60] & ~t[62] & t[63] & ~t[64]);
  assign t[51] = t[65] ^ x[10];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[6];
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[8];
  assign t[57] = t[71] ^ x[9];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[19];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[74] ^ x[18];
  assign t[61] = t[75] ^ x[20];
  assign t[62] = t[76] ^ x[21];
  assign t[63] = t[77] ^ x[22];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[66] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[67] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[68] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[73] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[74] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[75] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[76] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[77] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[78] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[31] | t[10]);
  assign t[8] = ~(t[32]);
  assign t[9] = ~(t[33]);
  assign y = (t[0] & ~t[13] & ~t[23]) | (~t[0] & t[13] & ~t[23]) | (~t[0] & ~t[13] & t[23]) | (t[0] & t[13] & t[23]);
endmodule

module R2ind79(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[24] | t[25]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[9] & t[11]);
  assign t[19] = ~(t[20] & t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[21] & t[8]);
  assign t[21] = ~(t[26] & t[25]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[29] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[29] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[29] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[29] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[29] & ~t[33]) | (~t[29] & t[33]);
  assign t[27] = t[35] ^ x[10];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[52] & ~t[53] & t[54] & ~t[55] & t[56]) | (~t[51] & t[52] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[51] & t[52] & ~t[55] & ~t[56]) | (~t[50] & t[52] & t[53] & ~t[54] & t[55]) | (t[52] & ~t[53] & t[55] & ~t[56]);
  assign t[39] = (t[51] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & t[51] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[51] & ~t[52] & ~t[55] & ~t[56]) | (t[50] & ~t[51] & t[52] & t[53] & ~t[56]) | (t[50] & ~t[51] & t[54] & t[55] & ~t[56]) | (t[51] & ~t[53] & ~t[55] & t[56]) | (~t[51] & t[53] & t[55] & t[56]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & t[51] & t[52] & ~t[53] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[53] & ~t[54] & t[55] & t[56]) | (~t[51] & ~t[52] & t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[52] & t[53] & ~t[55] & ~t[56]) | (~t[50] & ~t[51] & t[53] & ~t[54] & ~t[56]) | (~t[51] & t[52] & t[53] & t[54] & ~t[55]) | (~t[52] & t[53] & t[54] & ~t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[50] & t[51] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[51] & ~t[52] & t[55] & ~t[56]) | (~t[51] & t[52] & ~t[53] & t[54] & t[55]) | (t[52] & ~t[54] & t[55] & ~t[56]);
  assign t[43] = t[57] ^ x[10];
  assign t[44] = t[58] ^ x[5];
  assign t[45] = t[59] ^ x[6];
  assign t[46] = t[60] ^ x[7];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[8];
  assign t[49] = t[63] ^ x[9];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[20];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[22];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[59] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[63] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[64] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[65] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[66] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[67] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[68] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[23] | t[10]);
  assign t[8] = ~(t[24]);
  assign t[9] = ~(t[25]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind80(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[24] | t[25]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[17] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[18];
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[4]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[9] & t[11]);
  assign t[21] = t[6] | t[23];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[29] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[29] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[29] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[29] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[29] & ~t[33]) | (~t[29] & t[33]);
  assign t[27] = t[35] ^ x[10];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[52] & ~t[53] & t[54] & ~t[55] & t[56]) | (~t[51] & t[52] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[51] & t[52] & ~t[55] & ~t[56]) | (~t[50] & t[52] & t[53] & ~t[54] & t[55]) | (t[52] & ~t[53] & t[55] & ~t[56]);
  assign t[39] = (t[51] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & t[51] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[51] & ~t[52] & ~t[55] & ~t[56]) | (t[50] & ~t[51] & t[52] & t[53] & ~t[56]) | (t[50] & ~t[51] & t[54] & t[55] & ~t[56]) | (t[51] & ~t[53] & ~t[55] & t[56]) | (~t[51] & t[53] & t[55] & t[56]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & t[51] & t[52] & ~t[53] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[53] & ~t[54] & t[55] & t[56]) | (~t[51] & ~t[52] & t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[52] & t[53] & ~t[55] & ~t[56]) | (~t[50] & ~t[51] & t[53] & ~t[54] & ~t[56]) | (~t[51] & t[52] & t[53] & t[54] & ~t[55]) | (~t[52] & t[53] & t[54] & ~t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[50] & t[51] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[51] & ~t[52] & t[55] & ~t[56]) | (~t[51] & t[52] & ~t[53] & t[54] & t[55]) | (t[52] & ~t[54] & t[55] & ~t[56]);
  assign t[43] = t[57] ^ x[10];
  assign t[44] = t[58] ^ x[5];
  assign t[45] = t[59] ^ x[6];
  assign t[46] = t[60] ^ x[7];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[8];
  assign t[49] = t[63] ^ x[9];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[20];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[22];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[59] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[63] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[64] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[65] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[66] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[67] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[68] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[23] | t[10]);
  assign t[8] = ~(t[24]);
  assign t[9] = ~(t[25]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind81(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[9] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind82(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind83(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[25] & t[24]);
  assign t[12] = ~(t[26]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[17] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[18];
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[6] & t[20]);
  assign t[19] = ~(t[4]);
  assign t[1] = ~t[3];
  assign t[20] = t[21] | t[23];
  assign t[21] = ~(t[12] | t[8]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[29] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[29] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[25] = (t[29] & ~t[33]) | (~t[29] & t[33]);
  assign t[26] = (t[29] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[29] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[27] = t[35] ^ x[10];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[52] & ~t[53] & t[54] & ~t[55] & t[56]) | (~t[51] & t[52] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[51] & t[52] & ~t[55] & ~t[56]) | (~t[50] & t[52] & t[53] & ~t[54] & t[55]) | (t[52] & ~t[53] & t[55] & ~t[56]);
  assign t[39] = (t[51] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & t[51] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[51] & ~t[52] & ~t[55] & ~t[56]) | (t[50] & ~t[51] & t[52] & t[53] & ~t[56]) | (t[50] & ~t[51] & t[54] & t[55] & ~t[56]) | (t[51] & ~t[53] & ~t[55] & t[56]) | (~t[51] & t[53] & t[55] & t[56]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & t[51] & t[52] & ~t[53] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[53] & ~t[54] & t[55] & t[56]) | (~t[51] & ~t[52] & t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[52] & t[53] & ~t[55] & ~t[56]) | (~t[50] & ~t[51] & t[53] & ~t[54] & ~t[56]) | (~t[51] & t[52] & t[53] & t[54] & ~t[55]) | (~t[52] & t[53] & t[54] & ~t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[50] & t[51] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[51] & ~t[52] & t[55] & ~t[56]) | (~t[51] & t[52] & ~t[53] & t[54] & t[55]) | (t[52] & ~t[54] & t[55] & ~t[56]);
  assign t[43] = t[57] ^ x[10];
  assign t[44] = t[58] ^ x[5];
  assign t[45] = t[59] ^ x[6];
  assign t[46] = t[60] ^ x[7];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[8];
  assign t[49] = t[63] ^ x[9];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[20];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[22];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[59] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[5] = ~(t[6] & t[7]);
  assign t[60] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[63] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[64] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[65] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[66] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[67] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[68] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[10] & t[23]);
  assign t[8] = ~(t[24]);
  assign t[9] = ~(t[25]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind84(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[36]);
  assign t[14] = ~(t[34] | t[35]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[11]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[37] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[37] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[37] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[37] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[37] & ~t[43]) | (~t[37] & t[43]);
  assign t[37] = t[45] ^ x[9];
  assign t[38] = t[46] ^ x[10];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[8];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[12];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[15];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[68] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[69] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[71] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[72] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[73] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[75] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[76] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[77] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[79] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = ~(t[32] | t[12]);
  assign t[9] = ~x[2] & t[33];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind85(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[32] | t[33]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[11]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = t[7] | t[30];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[35] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[35] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[35] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[35] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[35] & ~t[41]) | (~t[35] & t[41]);
  assign t[35] = t[43] ^ x[9];
  assign t[36] = t[44] ^ x[10];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[53] & ~t[54] & t[55] & ~t[56] & t[57]) | (~t[52] & t[53] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[52] & t[53] & ~t[56] & ~t[57]) | (~t[51] & t[53] & t[54] & ~t[55] & t[56]) | (t[53] & ~t[54] & t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[47] = (t[52] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & t[52] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[52] & ~t[53] & ~t[56] & ~t[57]) | (t[51] & ~t[52] & t[53] & t[54] & ~t[57]) | (t[51] & ~t[52] & t[55] & t[56] & ~t[57]) | (t[52] & ~t[54] & ~t[56] & t[57]) | (~t[52] & t[54] & t[56] & t[57]);
  assign t[48] = (t[51] & t[52] & t[53] & ~t[54] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[54] & ~t[55] & t[56] & t[57]) | (~t[52] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[53] & t[54] & ~t[56] & ~t[57]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[57]) | (~t[52] & t[53] & t[54] & t[55] & ~t[56]) | (~t[53] & t[54] & t[55] & ~t[57]);
  assign t[49] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[51] & t[52] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[51] & ~t[52] & ~t[53] & t[56] & ~t[57]) | (~t[52] & t[53] & ~t[54] & t[55] & t[56]) | (t[53] & ~t[55] & t[56] & ~t[57]);
  assign t[51] = t[65] ^ x[9];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[8];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[12];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[66] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[67] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[68] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[69] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[71] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[74] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[75] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[76] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[77] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[30] | t[12]);
  assign t[9] = ~x[2] & t[31];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind86(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[28]);
  assign t[14] = ~(t[26] | t[27]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = ~(t[22] & t[24]);
  assign t[22] = ~(t[23] & t[10]);
  assign t[23] = ~(t[28] & t[27]);
  assign t[24] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[29] & ~t[34] & ~t[36]) | (~t[33] & t[34] & ~t[35]) | (~t[29] & ~t[34] & t[36]) | (t[33] & t[34] & t[35]);
  assign t[27] = (t[29] & ~t[34] & ~t[35]) | (~t[33] & t[34] & ~t[36]) | (~t[29] & ~t[34] & t[35]) | (t[33] & t[34] & t[36]);
  assign t[28] = (t[29] & ~t[35]) | (~t[29] & t[35]);
  assign t[29] = t[37] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[10];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[18];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[20];
  assign t[35] = t[43] ^ x[21];
  assign t[36] = t[44] ^ x[22];
  assign t[37] = (t[45] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[46] & ~t[47] & ~t[50] & ~t[51]) | (~t[45] & t[46] & t[47] & t[48] & ~t[51]) | (~t[45] & t[46] & t[49] & t[50] & ~t[51]) | (t[45] & ~t[47] & ~t[49] & t[51]) | (~t[45] & t[47] & t[49] & t[51]);
  assign t[38] = (t[45] & t[46] & ~t[47] & t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[47] & ~t[48] & t[49] & ~t[50] & t[51]) | (~t[46] & t[47] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[46] & t[47] & ~t[50] & ~t[51]) | (~t[45] & t[47] & t[48] & ~t[49] & t[50]) | (t[47] & ~t[48] & t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[41] = (t[46] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & t[46] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[46] & ~t[47] & ~t[50] & ~t[51]) | (t[45] & ~t[46] & t[47] & t[48] & ~t[51]) | (t[45] & ~t[46] & t[49] & t[50] & ~t[51]) | (t[46] & ~t[48] & ~t[50] & t[51]) | (~t[46] & t[48] & t[50] & t[51]);
  assign t[42] = (t[45] & t[46] & t[47] & ~t[48] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[48] & ~t[49] & t[50] & t[51]) | (~t[46] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[47] & t[48] & ~t[50] & ~t[51]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[51]) | (~t[46] & t[47] & t[48] & t[49] & ~t[50]) | (~t[47] & t[48] & t[49] & ~t[51]);
  assign t[43] = (t[45] & t[46] & ~t[47] & ~t[49] & t[50] & ~t[51]) | (t[45] & t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[51]) | (~t[45] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[45] & ~t[46] & ~t[48] & t[49] & ~t[51]) | (~t[45] & ~t[47] & t[48] & t[49] & t[50]) | (t[48] & t[49] & ~t[50] & ~t[51]);
  assign t[44] = (t[45] & t[46] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[45] & ~t[46] & ~t[47] & t[50] & ~t[51]) | (~t[46] & t[47] & ~t[48] & t[49] & t[50]) | (t[47] & ~t[49] & t[50] & ~t[51]);
  assign t[45] = t[59] ^ x[9];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[20];
  assign t[49] = t[63] ^ x[21];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[22];
  assign t[51] = t[65] ^ x[8];
  assign t[52] = t[66] ^ x[17];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[13];
  assign t[55] = t[69] ^ x[14];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[61] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[62] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[63] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[64] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[65] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[68] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[69] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[24] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind87(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[24] | t[25]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = t[7] | t[22];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[22] | t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind88(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind89(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind90(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] & t[24]);
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[7] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = t[21] | t[22];
  assign t[21] = ~(t[14] | t[10]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[25] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[26] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[22]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind91(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[36]);
  assign t[14] = ~(t[34] | t[35]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[11]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[37] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[37] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[37] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[37] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[37] & ~t[43]) | (~t[37] & t[43]);
  assign t[37] = t[45] ^ x[9];
  assign t[38] = t[46] ^ x[10];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[8];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[12];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[15];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[68] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[69] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[71] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[72] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[73] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[75] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[76] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[77] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[79] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = ~(t[32] | t[12]);
  assign t[9] = ~x[2] & t[33];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind92(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[32] | t[33]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[11]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = t[7] | t[30];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[35] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[35] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[35] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[35] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[35] & ~t[41]) | (~t[35] & t[41]);
  assign t[35] = t[43] ^ x[9];
  assign t[36] = t[44] ^ x[10];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[53] & ~t[54] & t[55] & ~t[56] & t[57]) | (~t[52] & t[53] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[52] & t[53] & ~t[56] & ~t[57]) | (~t[51] & t[53] & t[54] & ~t[55] & t[56]) | (t[53] & ~t[54] & t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[47] = (t[52] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & t[52] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[52] & ~t[53] & ~t[56] & ~t[57]) | (t[51] & ~t[52] & t[53] & t[54] & ~t[57]) | (t[51] & ~t[52] & t[55] & t[56] & ~t[57]) | (t[52] & ~t[54] & ~t[56] & t[57]) | (~t[52] & t[54] & t[56] & t[57]);
  assign t[48] = (t[51] & t[52] & t[53] & ~t[54] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[54] & ~t[55] & t[56] & t[57]) | (~t[52] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[53] & t[54] & ~t[56] & ~t[57]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[57]) | (~t[52] & t[53] & t[54] & t[55] & ~t[56]) | (~t[53] & t[54] & t[55] & ~t[57]);
  assign t[49] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[51] & t[52] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[51] & ~t[52] & ~t[53] & t[56] & ~t[57]) | (~t[52] & t[53] & ~t[54] & t[55] & t[56]) | (t[53] & ~t[55] & t[56] & ~t[57]);
  assign t[51] = t[65] ^ x[9];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[8];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[12];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[66] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[67] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[68] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[69] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[71] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[74] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[75] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[76] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[77] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[30] | t[12]);
  assign t[9] = ~x[2] & t[31];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind93(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[28]);
  assign t[14] = ~(t[26] | t[27]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = ~(t[22] & t[24]);
  assign t[22] = ~(t[23] & t[10]);
  assign t[23] = ~(t[28] & t[27]);
  assign t[24] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[29] & ~t[34] & ~t[36]) | (~t[33] & t[34] & ~t[35]) | (~t[29] & ~t[34] & t[36]) | (t[33] & t[34] & t[35]);
  assign t[27] = (t[29] & ~t[34] & ~t[35]) | (~t[33] & t[34] & ~t[36]) | (~t[29] & ~t[34] & t[35]) | (t[33] & t[34] & t[36]);
  assign t[28] = (t[29] & ~t[35]) | (~t[29] & t[35]);
  assign t[29] = t[37] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[10];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[18];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[20];
  assign t[35] = t[43] ^ x[21];
  assign t[36] = t[44] ^ x[22];
  assign t[37] = (t[45] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[46] & ~t[47] & ~t[50] & ~t[51]) | (~t[45] & t[46] & t[47] & t[48] & ~t[51]) | (~t[45] & t[46] & t[49] & t[50] & ~t[51]) | (t[45] & ~t[47] & ~t[49] & t[51]) | (~t[45] & t[47] & t[49] & t[51]);
  assign t[38] = (t[45] & t[46] & ~t[47] & t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[47] & ~t[48] & t[49] & ~t[50] & t[51]) | (~t[46] & t[47] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[46] & t[47] & ~t[50] & ~t[51]) | (~t[45] & t[47] & t[48] & ~t[49] & t[50]) | (t[47] & ~t[48] & t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[41] = (t[46] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & t[46] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[46] & ~t[47] & ~t[50] & ~t[51]) | (t[45] & ~t[46] & t[47] & t[48] & ~t[51]) | (t[45] & ~t[46] & t[49] & t[50] & ~t[51]) | (t[46] & ~t[48] & ~t[50] & t[51]) | (~t[46] & t[48] & t[50] & t[51]);
  assign t[42] = (t[45] & t[46] & t[47] & ~t[48] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[48] & ~t[49] & t[50] & t[51]) | (~t[46] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[47] & t[48] & ~t[50] & ~t[51]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[51]) | (~t[46] & t[47] & t[48] & t[49] & ~t[50]) | (~t[47] & t[48] & t[49] & ~t[51]);
  assign t[43] = (t[45] & t[46] & ~t[47] & ~t[49] & t[50] & ~t[51]) | (t[45] & t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[51]) | (~t[45] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[45] & ~t[46] & ~t[48] & t[49] & ~t[51]) | (~t[45] & ~t[47] & t[48] & t[49] & t[50]) | (t[48] & t[49] & ~t[50] & ~t[51]);
  assign t[44] = (t[45] & t[46] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[45] & ~t[46] & ~t[47] & t[50] & ~t[51]) | (~t[46] & t[47] & ~t[48] & t[49] & t[50]) | (t[47] & ~t[49] & t[50] & ~t[51]);
  assign t[45] = t[59] ^ x[9];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[20];
  assign t[49] = t[63] ^ x[21];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[22];
  assign t[51] = t[65] ^ x[8];
  assign t[52] = t[66] ^ x[17];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[13];
  assign t[55] = t[69] ^ x[14];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[61] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[62] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[63] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[64] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[65] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[68] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[69] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[24] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind94(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[24] | t[25]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = t[7] | t[22];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[22] | t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind95(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind96(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind97(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] & t[24]);
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[7] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = t[21] | t[22];
  assign t[21] = ~(t[14] | t[10]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[25] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[26] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[22]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind98(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[36]);
  assign t[14] = ~(t[34] | t[35]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[11]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[37] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[37] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[37] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[37] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[37] & ~t[43]) | (~t[37] & t[43]);
  assign t[37] = t[45] ^ x[9];
  assign t[38] = t[46] ^ x[10];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[8];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[12];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[15];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[68] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[69] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[71] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[72] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[73] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[75] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[76] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[77] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[79] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = ~(t[32] | t[12]);
  assign t[9] = ~x[2] & t[33];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind99(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[32] | t[33]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[11]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = t[7] | t[30];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[35] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[35] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[35] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[35] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[35] & ~t[41]) | (~t[35] & t[41]);
  assign t[35] = t[43] ^ x[9];
  assign t[36] = t[44] ^ x[10];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[53] & ~t[54] & t[55] & ~t[56] & t[57]) | (~t[52] & t[53] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[52] & t[53] & ~t[56] & ~t[57]) | (~t[51] & t[53] & t[54] & ~t[55] & t[56]) | (t[53] & ~t[54] & t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[47] = (t[52] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & t[52] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[52] & ~t[53] & ~t[56] & ~t[57]) | (t[51] & ~t[52] & t[53] & t[54] & ~t[57]) | (t[51] & ~t[52] & t[55] & t[56] & ~t[57]) | (t[52] & ~t[54] & ~t[56] & t[57]) | (~t[52] & t[54] & t[56] & t[57]);
  assign t[48] = (t[51] & t[52] & t[53] & ~t[54] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[54] & ~t[55] & t[56] & t[57]) | (~t[52] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[53] & t[54] & ~t[56] & ~t[57]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[57]) | (~t[52] & t[53] & t[54] & t[55] & ~t[56]) | (~t[53] & t[54] & t[55] & ~t[57]);
  assign t[49] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[51] & t[52] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[51] & ~t[52] & ~t[53] & t[56] & ~t[57]) | (~t[52] & t[53] & ~t[54] & t[55] & t[56]) | (t[53] & ~t[55] & t[56] & ~t[57]);
  assign t[51] = t[65] ^ x[9];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[8];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[12];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[66] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[67] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[68] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[69] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[71] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[74] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[75] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[76] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[77] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[30] | t[12]);
  assign t[9] = ~x[2] & t[31];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind100(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[28]);
  assign t[14] = ~(t[26] | t[27]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = ~(t[22] & t[24]);
  assign t[22] = ~(t[23] & t[10]);
  assign t[23] = ~(t[28] & t[27]);
  assign t[24] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[29] & ~t[34] & ~t[36]) | (~t[33] & t[34] & ~t[35]) | (~t[29] & ~t[34] & t[36]) | (t[33] & t[34] & t[35]);
  assign t[27] = (t[29] & ~t[34] & ~t[35]) | (~t[33] & t[34] & ~t[36]) | (~t[29] & ~t[34] & t[35]) | (t[33] & t[34] & t[36]);
  assign t[28] = (t[29] & ~t[35]) | (~t[29] & t[35]);
  assign t[29] = t[37] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[10];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[18];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[20];
  assign t[35] = t[43] ^ x[21];
  assign t[36] = t[44] ^ x[22];
  assign t[37] = (t[45] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[46] & ~t[47] & ~t[50] & ~t[51]) | (~t[45] & t[46] & t[47] & t[48] & ~t[51]) | (~t[45] & t[46] & t[49] & t[50] & ~t[51]) | (t[45] & ~t[47] & ~t[49] & t[51]) | (~t[45] & t[47] & t[49] & t[51]);
  assign t[38] = (t[45] & t[46] & ~t[47] & t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[47] & ~t[48] & t[49] & ~t[50] & t[51]) | (~t[46] & t[47] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[46] & t[47] & ~t[50] & ~t[51]) | (~t[45] & t[47] & t[48] & ~t[49] & t[50]) | (t[47] & ~t[48] & t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[41] = (t[46] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & t[46] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[46] & ~t[47] & ~t[50] & ~t[51]) | (t[45] & ~t[46] & t[47] & t[48] & ~t[51]) | (t[45] & ~t[46] & t[49] & t[50] & ~t[51]) | (t[46] & ~t[48] & ~t[50] & t[51]) | (~t[46] & t[48] & t[50] & t[51]);
  assign t[42] = (t[45] & t[46] & t[47] & ~t[48] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[48] & ~t[49] & t[50] & t[51]) | (~t[46] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[47] & t[48] & ~t[50] & ~t[51]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[51]) | (~t[46] & t[47] & t[48] & t[49] & ~t[50]) | (~t[47] & t[48] & t[49] & ~t[51]);
  assign t[43] = (t[45] & t[46] & ~t[47] & ~t[49] & t[50] & ~t[51]) | (t[45] & t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[51]) | (~t[45] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[45] & ~t[46] & ~t[48] & t[49] & ~t[51]) | (~t[45] & ~t[47] & t[48] & t[49] & t[50]) | (t[48] & t[49] & ~t[50] & ~t[51]);
  assign t[44] = (t[45] & t[46] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[45] & ~t[46] & ~t[47] & t[50] & ~t[51]) | (~t[46] & t[47] & ~t[48] & t[49] & t[50]) | (t[47] & ~t[49] & t[50] & ~t[51]);
  assign t[45] = t[59] ^ x[9];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[20];
  assign t[49] = t[63] ^ x[21];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[22];
  assign t[51] = t[65] ^ x[8];
  assign t[52] = t[66] ^ x[17];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[13];
  assign t[55] = t[69] ^ x[14];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[61] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[62] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[63] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[64] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[65] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[68] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[69] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[24] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind101(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[24] | t[25]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = t[7] | t[22];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[22] | t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind102(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind103(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind104(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] & t[24]);
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[7] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = t[21] | t[22];
  assign t[21] = ~(t[14] | t[10]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[25] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[26] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[22]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind105(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[36]);
  assign t[14] = ~(t[34] | t[35]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[11]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[37] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[37] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[37] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[37] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[37] & ~t[43]) | (~t[37] & t[43]);
  assign t[37] = t[45] ^ x[9];
  assign t[38] = t[46] ^ x[10];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[8];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[12];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[15];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[68] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[69] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[71] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[72] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[73] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[75] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[76] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[77] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[79] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = ~(t[32] | t[12]);
  assign t[9] = ~x[2] & t[33];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind106(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[32] | t[33]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[11]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = t[7] | t[30];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[35] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[35] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[35] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[35] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[35] & ~t[41]) | (~t[35] & t[41]);
  assign t[35] = t[43] ^ x[9];
  assign t[36] = t[44] ^ x[10];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[53] & ~t[54] & t[55] & ~t[56] & t[57]) | (~t[52] & t[53] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[52] & t[53] & ~t[56] & ~t[57]) | (~t[51] & t[53] & t[54] & ~t[55] & t[56]) | (t[53] & ~t[54] & t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[47] = (t[52] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & t[52] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[52] & ~t[53] & ~t[56] & ~t[57]) | (t[51] & ~t[52] & t[53] & t[54] & ~t[57]) | (t[51] & ~t[52] & t[55] & t[56] & ~t[57]) | (t[52] & ~t[54] & ~t[56] & t[57]) | (~t[52] & t[54] & t[56] & t[57]);
  assign t[48] = (t[51] & t[52] & t[53] & ~t[54] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[54] & ~t[55] & t[56] & t[57]) | (~t[52] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[53] & t[54] & ~t[56] & ~t[57]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[57]) | (~t[52] & t[53] & t[54] & t[55] & ~t[56]) | (~t[53] & t[54] & t[55] & ~t[57]);
  assign t[49] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[51] & t[52] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[51] & ~t[52] & ~t[53] & t[56] & ~t[57]) | (~t[52] & t[53] & ~t[54] & t[55] & t[56]) | (t[53] & ~t[55] & t[56] & ~t[57]);
  assign t[51] = t[65] ^ x[9];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[8];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[12];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[66] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[67] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[68] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[69] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[71] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[74] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[75] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[76] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[77] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[30] | t[12]);
  assign t[9] = ~x[2] & t[31];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind107(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[28]);
  assign t[14] = ~(t[26] | t[27]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = ~(t[22] & t[24]);
  assign t[22] = ~(t[23] & t[10]);
  assign t[23] = ~(t[28] & t[27]);
  assign t[24] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[29] & ~t[34] & ~t[36]) | (~t[33] & t[34] & ~t[35]) | (~t[29] & ~t[34] & t[36]) | (t[33] & t[34] & t[35]);
  assign t[27] = (t[29] & ~t[34] & ~t[35]) | (~t[33] & t[34] & ~t[36]) | (~t[29] & ~t[34] & t[35]) | (t[33] & t[34] & t[36]);
  assign t[28] = (t[29] & ~t[35]) | (~t[29] & t[35]);
  assign t[29] = t[37] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[10];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[18];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[20];
  assign t[35] = t[43] ^ x[21];
  assign t[36] = t[44] ^ x[22];
  assign t[37] = (t[45] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[46] & ~t[47] & ~t[50] & ~t[51]) | (~t[45] & t[46] & t[47] & t[48] & ~t[51]) | (~t[45] & t[46] & t[49] & t[50] & ~t[51]) | (t[45] & ~t[47] & ~t[49] & t[51]) | (~t[45] & t[47] & t[49] & t[51]);
  assign t[38] = (t[45] & t[46] & ~t[47] & t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[47] & ~t[48] & t[49] & ~t[50] & t[51]) | (~t[46] & t[47] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[46] & t[47] & ~t[50] & ~t[51]) | (~t[45] & t[47] & t[48] & ~t[49] & t[50]) | (t[47] & ~t[48] & t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[41] = (t[46] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & t[46] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[46] & ~t[47] & ~t[50] & ~t[51]) | (t[45] & ~t[46] & t[47] & t[48] & ~t[51]) | (t[45] & ~t[46] & t[49] & t[50] & ~t[51]) | (t[46] & ~t[48] & ~t[50] & t[51]) | (~t[46] & t[48] & t[50] & t[51]);
  assign t[42] = (t[45] & t[46] & t[47] & ~t[48] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[48] & ~t[49] & t[50] & t[51]) | (~t[46] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[47] & t[48] & ~t[50] & ~t[51]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[51]) | (~t[46] & t[47] & t[48] & t[49] & ~t[50]) | (~t[47] & t[48] & t[49] & ~t[51]);
  assign t[43] = (t[45] & t[46] & ~t[47] & ~t[49] & t[50] & ~t[51]) | (t[45] & t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[51]) | (~t[45] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[45] & ~t[46] & ~t[48] & t[49] & ~t[51]) | (~t[45] & ~t[47] & t[48] & t[49] & t[50]) | (t[48] & t[49] & ~t[50] & ~t[51]);
  assign t[44] = (t[45] & t[46] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[45] & ~t[46] & ~t[47] & t[50] & ~t[51]) | (~t[46] & t[47] & ~t[48] & t[49] & t[50]) | (t[47] & ~t[49] & t[50] & ~t[51]);
  assign t[45] = t[59] ^ x[9];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[20];
  assign t[49] = t[63] ^ x[21];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[22];
  assign t[51] = t[65] ^ x[8];
  assign t[52] = t[66] ^ x[17];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[13];
  assign t[55] = t[69] ^ x[14];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[61] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[62] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[63] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[64] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[65] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[68] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[69] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[24] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind108(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[24] | t[25]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = t[7] | t[22];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[22] | t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind109(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind110(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind111(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] & t[24]);
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[7] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = t[21] | t[22];
  assign t[21] = ~(t[14] | t[10]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[25] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[26] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[22]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind112(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[36]);
  assign t[14] = ~(t[34] | t[35]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[11]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[9] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[37] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[37] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[37] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[37] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[37] & ~t[43]) | (~t[37] & t[43]);
  assign t[37] = t[45] ^ x[9];
  assign t[38] = t[46] ^ x[10];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[8];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[12];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[15];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[68] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[69] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[71] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[72] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[73] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[75] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[76] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[77] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[79] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = ~(t[32] | t[12]);
  assign t[9] = ~x[2] & t[33];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind113(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[32] | t[33]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[11]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[9] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = t[7] | t[30];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[35] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[35] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[35] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[35] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[35] & ~t[41]) | (~t[35] & t[41]);
  assign t[35] = t[43] ^ x[9];
  assign t[36] = t[44] ^ x[10];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[53] & ~t[54] & t[55] & ~t[56] & t[57]) | (~t[52] & t[53] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[52] & t[53] & ~t[56] & ~t[57]) | (~t[51] & t[53] & t[54] & ~t[55] & t[56]) | (t[53] & ~t[54] & t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[47] = (t[52] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & t[52] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[52] & ~t[53] & ~t[56] & ~t[57]) | (t[51] & ~t[52] & t[53] & t[54] & ~t[57]) | (t[51] & ~t[52] & t[55] & t[56] & ~t[57]) | (t[52] & ~t[54] & ~t[56] & t[57]) | (~t[52] & t[54] & t[56] & t[57]);
  assign t[48] = (t[51] & t[52] & t[53] & ~t[54] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[54] & ~t[55] & t[56] & t[57]) | (~t[52] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[53] & t[54] & ~t[56] & ~t[57]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[57]) | (~t[52] & t[53] & t[54] & t[55] & ~t[56]) | (~t[53] & t[54] & t[55] & ~t[57]);
  assign t[49] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[51] & t[52] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[51] & ~t[52] & ~t[53] & t[56] & ~t[57]) | (~t[52] & t[53] & ~t[54] & t[55] & t[56]) | (t[53] & ~t[55] & t[56] & ~t[57]);
  assign t[51] = t[65] ^ x[9];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[8];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[12];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[66] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[67] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[68] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[69] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[71] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[74] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[75] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[76] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[77] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[30] | t[12]);
  assign t[9] = ~x[2] & t[31];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind114(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[28]);
  assign t[14] = ~(t[26] | t[27]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[9] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = ~(t[22] & t[24]);
  assign t[22] = ~(t[23] & t[10]);
  assign t[23] = ~(t[28] & t[27]);
  assign t[24] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[29] & ~t[34] & ~t[36]) | (~t[33] & t[34] & ~t[35]) | (~t[29] & ~t[34] & t[36]) | (t[33] & t[34] & t[35]);
  assign t[27] = (t[29] & ~t[34] & ~t[35]) | (~t[33] & t[34] & ~t[36]) | (~t[29] & ~t[34] & t[35]) | (t[33] & t[34] & t[36]);
  assign t[28] = (t[29] & ~t[35]) | (~t[29] & t[35]);
  assign t[29] = t[37] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[10];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[18];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[20];
  assign t[35] = t[43] ^ x[21];
  assign t[36] = t[44] ^ x[22];
  assign t[37] = (t[45] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[46] & ~t[47] & ~t[50] & ~t[51]) | (~t[45] & t[46] & t[47] & t[48] & ~t[51]) | (~t[45] & t[46] & t[49] & t[50] & ~t[51]) | (t[45] & ~t[47] & ~t[49] & t[51]) | (~t[45] & t[47] & t[49] & t[51]);
  assign t[38] = (t[45] & t[46] & ~t[47] & t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[47] & ~t[48] & t[49] & ~t[50] & t[51]) | (~t[46] & t[47] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[46] & t[47] & ~t[50] & ~t[51]) | (~t[45] & t[47] & t[48] & ~t[49] & t[50]) | (t[47] & ~t[48] & t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[41] = (t[46] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & t[46] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[46] & ~t[47] & ~t[50] & ~t[51]) | (t[45] & ~t[46] & t[47] & t[48] & ~t[51]) | (t[45] & ~t[46] & t[49] & t[50] & ~t[51]) | (t[46] & ~t[48] & ~t[50] & t[51]) | (~t[46] & t[48] & t[50] & t[51]);
  assign t[42] = (t[45] & t[46] & t[47] & ~t[48] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[48] & ~t[49] & t[50] & t[51]) | (~t[46] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[47] & t[48] & ~t[50] & ~t[51]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[51]) | (~t[46] & t[47] & t[48] & t[49] & ~t[50]) | (~t[47] & t[48] & t[49] & ~t[51]);
  assign t[43] = (t[45] & t[46] & ~t[47] & ~t[49] & t[50] & ~t[51]) | (t[45] & t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[51]) | (~t[45] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[45] & ~t[46] & ~t[48] & t[49] & ~t[51]) | (~t[45] & ~t[47] & t[48] & t[49] & t[50]) | (t[48] & t[49] & ~t[50] & ~t[51]);
  assign t[44] = (t[45] & t[46] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[45] & ~t[46] & ~t[47] & t[50] & ~t[51]) | (~t[46] & t[47] & ~t[48] & t[49] & t[50]) | (t[47] & ~t[49] & t[50] & ~t[51]);
  assign t[45] = t[59] ^ x[9];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[20];
  assign t[49] = t[63] ^ x[21];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[22];
  assign t[51] = t[65] ^ x[8];
  assign t[52] = t[66] ^ x[17];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[13];
  assign t[55] = t[69] ^ x[14];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[61] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[62] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[63] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[64] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[65] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[68] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[69] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[24] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind115(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[24] | t[25]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[9] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = t[7] | t[22];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[22] | t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind116(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[9] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind117(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[9] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind118(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[23] & t[22]);
  assign t[12] = ~(t[24]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[6] & t[18]);
  assign t[18] = t[19] | t[21];
  assign t[19] = ~(t[12] | t[8]);
  assign t[1] = ~t[3];
  assign t[20] = (t[25] & ~t[26]) | (~t[25] & t[26]);
  assign t[21] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[22] = (t[27] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[27] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[23] = (t[27] & ~t[31]) | (~t[27] & t[31]);
  assign t[24] = (t[27] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[27] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[18];
  assign t[29] = t[37] ^ x[19];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[20];
  assign t[31] = t[39] ^ x[21];
  assign t[32] = t[40] ^ x[22];
  assign t[33] = (t[41] & ~t[43] & ~t[44] & ~t[45] & ~t[46]) | (t[41] & ~t[42] & ~t[44] & ~t[45] & ~t[47]) | (t[41] & ~t[42] & ~t[43] & ~t[46] & ~t[47]) | (~t[41] & t[42] & t[43] & t[44] & ~t[47]) | (~t[41] & t[42] & t[45] & t[46] & ~t[47]) | (t[41] & ~t[43] & ~t[45] & t[47]) | (~t[41] & t[43] & t[45] & t[47]);
  assign t[34] = (t[41] & t[42] & ~t[43] & ~t[45] & t[46] & ~t[47]) | (t[41] & t[43] & ~t[44] & ~t[45] & ~t[46] & t[47]) | (~t[42] & ~t[43] & t[45] & ~t[46] & ~t[47]) | (~t[41] & ~t[43] & ~t[44] & t[45] & ~t[46]) | (~t[41] & ~t[42] & ~t[44] & t[45] & ~t[47]) | (~t[41] & ~t[43] & t[44] & t[45] & t[46]) | (t[44] & t[45] & ~t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[36] = (t[48] & t[49] & ~t[50] & t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[50] & ~t[51] & t[52] & ~t[53] & t[54]) | (~t[49] & t[50] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[49] & t[50] & ~t[53] & ~t[54]) | (~t[48] & t[50] & t[51] & ~t[52] & t[53]) | (t[50] & ~t[51] & t[53] & ~t[54]);
  assign t[37] = (t[49] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & t[49] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[49] & ~t[50] & ~t[53] & ~t[54]) | (t[48] & ~t[49] & t[50] & t[51] & ~t[54]) | (t[48] & ~t[49] & t[52] & t[53] & ~t[54]) | (t[49] & ~t[51] & ~t[53] & t[54]) | (~t[49] & t[51] & t[53] & t[54]);
  assign t[38] = (t[48] & t[49] & t[50] & ~t[51] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & ~t[51] & ~t[52] & t[53] & t[54]) | (~t[49] & ~t[50] & t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[50] & t[51] & ~t[53] & ~t[54]) | (~t[48] & ~t[49] & t[51] & ~t[52] & ~t[54]) | (~t[49] & t[50] & t[51] & t[52] & ~t[53]) | (~t[50] & t[51] & t[52] & ~t[54]);
  assign t[39] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[48] & t[49] & ~t[51] & t[52] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & ~t[51] & ~t[52] & t[53]) | (~t[48] & ~t[51] & ~t[52] & t[53] & ~t[54]) | (~t[48] & ~t[49] & ~t[50] & t[53] & ~t[54]) | (~t[49] & t[50] & ~t[51] & t[52] & t[53]) | (t[50] & ~t[52] & t[53] & ~t[54]);
  assign t[41] = t[55] ^ x[10];
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[7];
  assign t[45] = t[59] ^ x[11];
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[17];
  assign t[49] = t[63] ^ x[19];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[21];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[16];
  assign t[55] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[56] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[57] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[58] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[59] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[5] = ~(t[6] & t[7]);
  assign t[60] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[63] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[64] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[65] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[66] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[67] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[68] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[21]);
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[23]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind119(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[34]);
  assign t[12] = ~(t[32] | t[33]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[32] & t[9]);
  assign t[19] = ~(t[34] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[33] & t[8]);
  assign t[21] = ~(t[22] ^ t[23]);
  assign t[22] = ~t[24];
  assign t[23] = t[4] ? x[27] : x[26];
  assign t[24] = x[2] ? x[28] : t[25];
  assign t[25] = ~(t[26] & t[27]);
  assign t[26] = ~(t[9] & t[11]);
  assign t[27] = ~(t[28] & t[31]);
  assign t[28] = ~(t[29] & t[8]);
  assign t[29] = ~(t[34] & t[33]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[37] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[37] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[37] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[37] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[37] & ~t[41]) | (~t[37] & t[41]);
  assign t[35] = t[43] ^ x[10];
  assign t[36] = t[44] ^ x[11];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[60] & ~t[61] & t[62] & ~t[63] & t[64]) | (~t[59] & t[60] & ~t[61] & ~t[62] & ~t[64]) | (~t[58] & t[60] & ~t[61] & ~t[62] & ~t[63]) | (~t[58] & ~t[59] & t[60] & ~t[63] & ~t[64]) | (~t[58] & t[60] & t[61] & ~t[62] & t[63]) | (t[60] & ~t[61] & t[63] & ~t[64]);
  assign t[47] = (t[59] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (~t[58] & t[59] & ~t[61] & ~t[62] & ~t[64]) | (~t[58] & t[59] & ~t[60] & ~t[63] & ~t[64]) | (t[58] & ~t[59] & t[60] & t[61] & ~t[64]) | (t[58] & ~t[59] & t[62] & t[63] & ~t[64]) | (t[59] & ~t[61] & ~t[63] & t[64]) | (~t[59] & t[61] & t[63] & t[64]);
  assign t[48] = (t[58] & t[59] & t[60] & ~t[61] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & ~t[61] & ~t[62] & t[63] & t[64]) | (~t[59] & ~t[60] & t[61] & ~t[62] & ~t[63]) | (~t[58] & ~t[60] & t[61] & ~t[63] & ~t[64]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[64]) | (~t[59] & t[60] & t[61] & t[62] & ~t[63]) | (~t[60] & t[61] & t[62] & ~t[64]);
  assign t[49] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[4] = ~x[2] & t[30];
  assign t[50] = (t[58] & t[59] & ~t[61] & t[62] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[61] & ~t[62] & t[63] & ~t[64]) | (~t[58] & ~t[59] & ~t[60] & t[63] & ~t[64]) | (~t[59] & t[60] & ~t[61] & t[62] & t[63]) | (t[60] & ~t[62] & t[63] & ~t[64]);
  assign t[51] = t[65] ^ x[10];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[6];
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[8];
  assign t[57] = t[71] ^ x[9];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[19];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[74] ^ x[18];
  assign t[61] = t[75] ^ x[20];
  assign t[62] = t[76] ^ x[21];
  assign t[63] = t[77] ^ x[22];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[66] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[67] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[68] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[73] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[74] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[75] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[76] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[77] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[78] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[31] | t[10]);
  assign t[8] = ~(t[32]);
  assign t[9] = ~(t[33]);
  assign y = (t[0] & ~t[13] & ~t[21]) | (~t[0] & t[13] & ~t[21]) | (~t[0] & ~t[13] & t[21]) | (t[0] & t[13] & t[21]);
endmodule

module R2ind120(x, y);
 input [28:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[30] | t[31]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[30] & t[9]);
  assign t[19] = ~(t[32] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[31] & t[8]);
  assign t[21] = ~(t[22] ^ t[23]);
  assign t[22] = ~t[24];
  assign t[23] = t[4] ? x[27] : x[26];
  assign t[24] = x[2] ? x[28] : t[25];
  assign t[25] = ~(t[26] & t[27]);
  assign t[26] = ~(t[9] & t[11]);
  assign t[27] = t[6] | t[29];
  assign t[28] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[29] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[38] & ~t[40]) | (~t[37] & t[38] & ~t[39]) | (~t[35] & ~t[38] & t[40]) | (t[37] & t[38] & t[39]);
  assign t[31] = (t[35] & ~t[38] & ~t[39]) | (~t[37] & t[38] & ~t[40]) | (~t[35] & ~t[38] & t[39]) | (t[37] & t[38] & t[40]);
  assign t[32] = (t[35] & ~t[39]) | (~t[35] & t[39]);
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[11];
  assign t[35] = t[43] ^ x[17];
  assign t[36] = t[44] ^ x[18];
  assign t[37] = t[45] ^ x[19];
  assign t[38] = t[46] ^ x[20];
  assign t[39] = t[47] ^ x[21];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[22];
  assign t[41] = (t[49] & ~t[51] & ~t[52] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & ~t[52] & ~t[53] & ~t[55]) | (t[49] & ~t[50] & ~t[51] & ~t[54] & ~t[55]) | (~t[49] & t[50] & t[51] & t[52] & ~t[55]) | (~t[49] & t[50] & t[53] & t[54] & ~t[55]) | (t[49] & ~t[51] & ~t[53] & t[55]) | (~t[49] & t[51] & t[53] & t[55]);
  assign t[42] = (t[49] & t[50] & ~t[51] & ~t[53] & t[54] & ~t[55]) | (t[49] & t[51] & ~t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[51] & t[53] & ~t[54] & ~t[55]) | (~t[49] & ~t[51] & ~t[52] & t[53] & ~t[54]) | (~t[49] & ~t[50] & ~t[52] & t[53] & ~t[55]) | (~t[49] & ~t[51] & t[52] & t[53] & t[54]) | (t[52] & t[53] & ~t[54] & ~t[55]);
  assign t[43] = (t[56] & ~t[58] & ~t[59] & ~t[60] & ~t[61]) | (t[56] & ~t[57] & ~t[59] & ~t[60] & ~t[62]) | (t[56] & ~t[57] & ~t[58] & ~t[61] & ~t[62]) | (~t[56] & t[57] & t[58] & t[59] & ~t[62]) | (~t[56] & t[57] & t[60] & t[61] & ~t[62]) | (t[56] & ~t[58] & ~t[60] & t[62]) | (~t[56] & t[58] & t[60] & t[62]);
  assign t[44] = (t[56] & t[57] & ~t[58] & t[59] & ~t[60] & ~t[62]) | (t[56] & ~t[58] & ~t[59] & t[60] & ~t[61] & t[62]) | (~t[57] & t[58] & ~t[59] & ~t[60] & ~t[62]) | (~t[56] & t[58] & ~t[59] & ~t[60] & ~t[61]) | (~t[56] & ~t[57] & t[58] & ~t[61] & ~t[62]) | (~t[56] & t[58] & t[59] & ~t[60] & t[61]) | (t[58] & ~t[59] & t[61] & ~t[62]);
  assign t[45] = (t[57] & ~t[58] & ~t[59] & ~t[60] & ~t[61]) | (~t[56] & t[57] & ~t[59] & ~t[60] & ~t[62]) | (~t[56] & t[57] & ~t[58] & ~t[61] & ~t[62]) | (t[56] & ~t[57] & t[58] & t[59] & ~t[62]) | (t[56] & ~t[57] & t[60] & t[61] & ~t[62]) | (t[57] & ~t[59] & ~t[61] & t[62]) | (~t[57] & t[59] & t[61] & t[62]);
  assign t[46] = (t[56] & t[57] & t[58] & ~t[59] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[59] & ~t[60] & t[61] & t[62]) | (~t[57] & ~t[58] & t[59] & ~t[60] & ~t[61]) | (~t[56] & ~t[58] & t[59] & ~t[61] & ~t[62]) | (~t[56] & ~t[57] & t[59] & ~t[60] & ~t[62]) | (~t[57] & t[58] & t[59] & t[60] & ~t[61]) | (~t[58] & t[59] & t[60] & ~t[62]);
  assign t[47] = (t[56] & t[57] & ~t[58] & ~t[60] & t[61] & ~t[62]) | (t[56] & t[58] & ~t[59] & ~t[60] & ~t[61] & t[62]) | (~t[57] & ~t[58] & t[60] & ~t[61] & ~t[62]) | (~t[56] & ~t[58] & ~t[59] & t[60] & ~t[61]) | (~t[56] & ~t[57] & ~t[59] & t[60] & ~t[62]) | (~t[56] & ~t[58] & t[59] & t[60] & t[61]) | (t[59] & t[60] & ~t[61] & ~t[62]);
  assign t[48] = (t[56] & t[57] & ~t[59] & t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & t[59] & ~t[60] & ~t[61] & t[62]) | (~t[57] & ~t[58] & ~t[59] & ~t[60] & t[61]) | (~t[56] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[56] & ~t[57] & ~t[58] & t[61] & ~t[62]) | (~t[57] & t[58] & ~t[59] & t[60] & t[61]) | (t[58] & ~t[60] & t[61] & ~t[62]);
  assign t[49] = t[63] ^ x[10];
  assign t[4] = ~x[2] & t[28];
  assign t[50] = t[64] ^ x[5];
  assign t[51] = t[65] ^ x[6];
  assign t[52] = t[66] ^ x[7];
  assign t[53] = t[67] ^ x[11];
  assign t[54] = t[68] ^ x[8];
  assign t[55] = t[69] ^ x[9];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[16];
  assign t[63] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[64] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[65] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[66] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[67] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[71] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[72] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[73] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[74] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[75] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[76] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[29] | t[10]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[31]);
  assign y = (t[0] & ~t[13] & ~t[21]) | (~t[0] & t[13] & ~t[21]) | (~t[0] & ~t[13] & t[21]) | (t[0] & t[13] & t[21]);
endmodule

module R2ind121(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[24] | t[25]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[9] & t[11]);
  assign t[19] = ~(t[20] & t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[21] & t[8]);
  assign t[21] = ~(t[26] & t[25]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[29] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[29] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[29] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[29] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[29] & ~t[33]) | (~t[29] & t[33]);
  assign t[27] = t[35] ^ x[10];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[52] & ~t[53] & t[54] & ~t[55] & t[56]) | (~t[51] & t[52] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[51] & t[52] & ~t[55] & ~t[56]) | (~t[50] & t[52] & t[53] & ~t[54] & t[55]) | (t[52] & ~t[53] & t[55] & ~t[56]);
  assign t[39] = (t[51] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (~t[50] & t[51] & ~t[53] & ~t[54] & ~t[56]) | (~t[50] & t[51] & ~t[52] & ~t[55] & ~t[56]) | (t[50] & ~t[51] & t[52] & t[53] & ~t[56]) | (t[50] & ~t[51] & t[54] & t[55] & ~t[56]) | (t[51] & ~t[53] & ~t[55] & t[56]) | (~t[51] & t[53] & t[55] & t[56]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & t[51] & t[52] & ~t[53] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[53] & ~t[54] & t[55] & t[56]) | (~t[51] & ~t[52] & t[53] & ~t[54] & ~t[55]) | (~t[50] & ~t[52] & t[53] & ~t[55] & ~t[56]) | (~t[50] & ~t[51] & t[53] & ~t[54] & ~t[56]) | (~t[51] & t[52] & t[53] & t[54] & ~t[55]) | (~t[52] & t[53] & t[54] & ~t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[50] & t[51] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[51] & ~t[52] & t[55] & ~t[56]) | (~t[51] & t[52] & ~t[53] & t[54] & t[55]) | (t[52] & ~t[54] & t[55] & ~t[56]);
  assign t[43] = t[57] ^ x[10];
  assign t[44] = t[58] ^ x[5];
  assign t[45] = t[59] ^ x[6];
  assign t[46] = t[60] ^ x[7];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[8];
  assign t[49] = t[63] ^ x[9];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[20];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[22];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[59] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[63] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[64] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[65] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[66] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[67] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[68] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[7] = ~(t[23] | t[10]);
  assign t[8] = ~(t[24]);
  assign t[9] = ~(t[25]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind122(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[24]);
  assign t[12] = ~(t[22] | t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[9] & t[11]);
  assign t[19] = t[6] | t[21];
  assign t[1] = ~t[3];
  assign t[20] = (t[25] & ~t[26]) | (~t[25] & t[26]);
  assign t[21] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[22] = (t[27] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[27] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[23] = (t[27] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[27] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[24] = (t[27] & ~t[31]) | (~t[27] & t[31]);
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[18];
  assign t[29] = t[37] ^ x[19];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[20];
  assign t[31] = t[39] ^ x[21];
  assign t[32] = t[40] ^ x[22];
  assign t[33] = (t[41] & ~t[43] & ~t[44] & ~t[45] & ~t[46]) | (t[41] & ~t[42] & ~t[44] & ~t[45] & ~t[47]) | (t[41] & ~t[42] & ~t[43] & ~t[46] & ~t[47]) | (~t[41] & t[42] & t[43] & t[44] & ~t[47]) | (~t[41] & t[42] & t[45] & t[46] & ~t[47]) | (t[41] & ~t[43] & ~t[45] & t[47]) | (~t[41] & t[43] & t[45] & t[47]);
  assign t[34] = (t[41] & t[42] & ~t[43] & ~t[45] & t[46] & ~t[47]) | (t[41] & t[43] & ~t[44] & ~t[45] & ~t[46] & t[47]) | (~t[42] & ~t[43] & t[45] & ~t[46] & ~t[47]) | (~t[41] & ~t[43] & ~t[44] & t[45] & ~t[46]) | (~t[41] & ~t[42] & ~t[44] & t[45] & ~t[47]) | (~t[41] & ~t[43] & t[44] & t[45] & t[46]) | (t[44] & t[45] & ~t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[36] = (t[48] & t[49] & ~t[50] & t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[50] & ~t[51] & t[52] & ~t[53] & t[54]) | (~t[49] & t[50] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[49] & t[50] & ~t[53] & ~t[54]) | (~t[48] & t[50] & t[51] & ~t[52] & t[53]) | (t[50] & ~t[51] & t[53] & ~t[54]);
  assign t[37] = (t[49] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & t[49] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[49] & ~t[50] & ~t[53] & ~t[54]) | (t[48] & ~t[49] & t[50] & t[51] & ~t[54]) | (t[48] & ~t[49] & t[52] & t[53] & ~t[54]) | (t[49] & ~t[51] & ~t[53] & t[54]) | (~t[49] & t[51] & t[53] & t[54]);
  assign t[38] = (t[48] & t[49] & t[50] & ~t[51] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & ~t[51] & ~t[52] & t[53] & t[54]) | (~t[49] & ~t[50] & t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[50] & t[51] & ~t[53] & ~t[54]) | (~t[48] & ~t[49] & t[51] & ~t[52] & ~t[54]) | (~t[49] & t[50] & t[51] & t[52] & ~t[53]) | (~t[50] & t[51] & t[52] & ~t[54]);
  assign t[39] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[48] & t[49] & ~t[51] & t[52] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & ~t[51] & ~t[52] & t[53]) | (~t[48] & ~t[51] & ~t[52] & t[53] & ~t[54]) | (~t[48] & ~t[49] & ~t[50] & t[53] & ~t[54]) | (~t[49] & t[50] & ~t[51] & t[52] & t[53]) | (t[50] & ~t[52] & t[53] & ~t[54]);
  assign t[41] = t[55] ^ x[10];
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[7];
  assign t[45] = t[59] ^ x[11];
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[17];
  assign t[49] = t[63] ^ x[19];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[21];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[16];
  assign t[55] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[56] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[57] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[58] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[59] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[63] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[64] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[65] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[66] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[67] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[68] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[21] | t[10]);
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[23]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind123(x, y);
 input [25:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[22]);
  assign t[11] = ~(t[12] ^ t[13]);
  assign t[12] = ~t[14];
  assign t[13] = t[4] ? x[23] : x[22];
  assign t[14] = x[2] ? x[24] : t[15];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = ~(t[8] & t[18]);
  assign t[17] = ~(t[19] & t[25]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(t[20] & t[10]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = (t[26] & ~t[27]) | (~t[26] & t[27]);
  assign t[22] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[23] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[24] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[25] = (t[28] & ~t[33]) | (~t[28] & t[33]);
  assign t[26] = t[34] ^ x[10];
  assign t[27] = t[35] ^ x[11];
  assign t[28] = t[36] ^ x[17];
  assign t[29] = t[37] ^ x[18];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[19];
  assign t[31] = t[39] ^ x[20];
  assign t[32] = t[40] ^ x[21];
  assign t[33] = t[41] ^ x[25];
  assign t[34] = (t[42] & ~t[44] & ~t[45] & ~t[46] & ~t[47]) | (t[42] & ~t[43] & ~t[45] & ~t[46] & ~t[48]) | (t[42] & ~t[43] & ~t[44] & ~t[47] & ~t[48]) | (~t[42] & t[43] & t[44] & t[45] & ~t[48]) | (~t[42] & t[43] & t[46] & t[47] & ~t[48]) | (t[42] & ~t[44] & ~t[46] & t[48]) | (~t[42] & t[44] & t[46] & t[48]);
  assign t[35] = (t[42] & t[43] & ~t[44] & ~t[46] & t[47] & ~t[48]) | (t[42] & t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[48]) | (~t[42] & ~t[44] & ~t[45] & t[46] & ~t[47]) | (~t[42] & ~t[43] & ~t[45] & t[46] & ~t[48]) | (~t[42] & ~t[44] & t[45] & t[46] & t[47]) | (t[45] & t[46] & ~t[47] & ~t[48]);
  assign t[36] = (t[49] & ~t[51] & ~t[52] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & ~t[52] & ~t[53] & ~t[55]) | (t[49] & ~t[50] & ~t[51] & ~t[54] & ~t[55]) | (~t[49] & t[50] & t[51] & t[52] & ~t[55]) | (~t[49] & t[50] & t[53] & t[54] & ~t[55]) | (t[49] & ~t[51] & ~t[53] & t[55]) | (~t[49] & t[51] & t[53] & t[55]);
  assign t[37] = (t[50] & ~t[51] & ~t[52] & ~t[53] & ~t[54]) | (~t[49] & t[50] & ~t[52] & ~t[53] & ~t[55]) | (~t[49] & t[50] & ~t[51] & ~t[54] & ~t[55]) | (t[49] & ~t[50] & t[51] & t[52] & ~t[55]) | (t[49] & ~t[50] & t[53] & t[54] & ~t[55]) | (t[50] & ~t[52] & ~t[54] & t[55]) | (~t[50] & t[52] & t[54] & t[55]);
  assign t[38] = (t[49] & t[50] & t[51] & ~t[52] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[52] & ~t[53] & t[54] & t[55]) | (~t[50] & ~t[51] & t[52] & ~t[53] & ~t[54]) | (~t[49] & ~t[51] & t[52] & ~t[54] & ~t[55]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[55]) | (~t[50] & t[51] & t[52] & t[53] & ~t[54]) | (~t[51] & t[52] & t[53] & ~t[55]);
  assign t[39] = (t[49] & t[50] & ~t[51] & ~t[53] & t[54] & ~t[55]) | (t[49] & t[51] & ~t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[51] & t[53] & ~t[54] & ~t[55]) | (~t[49] & ~t[51] & ~t[52] & t[53] & ~t[54]) | (~t[49] & ~t[50] & ~t[52] & t[53] & ~t[55]) | (~t[49] & ~t[51] & t[52] & t[53] & t[54]) | (t[52] & t[53] & ~t[54] & ~t[55]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[49] & t[50] & ~t[52] & t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & t[52] & ~t[53] & ~t[54] & t[55]) | (~t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[49] & ~t[50] & ~t[51] & t[54] & ~t[55]) | (~t[50] & t[51] & ~t[52] & t[53] & t[54]) | (t[51] & ~t[53] & t[54] & ~t[55]);
  assign t[41] = (t[49] & t[50] & ~t[51] & t[52] & ~t[53] & ~t[55]) | (t[49] & ~t[51] & ~t[52] & t[53] & ~t[54] & t[55]) | (~t[50] & t[51] & ~t[52] & ~t[53] & ~t[55]) | (~t[49] & t[51] & ~t[52] & ~t[53] & ~t[54]) | (~t[49] & ~t[50] & t[51] & ~t[54] & ~t[55]) | (~t[49] & t[51] & t[52] & ~t[53] & t[54]) | (t[51] & ~t[52] & t[54] & ~t[55]);
  assign t[42] = t[56] ^ x[10];
  assign t[43] = t[57] ^ x[5];
  assign t[44] = t[58] ^ x[6];
  assign t[45] = t[59] ^ x[7];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[8];
  assign t[48] = t[62] ^ x[9];
  assign t[49] = t[63] ^ x[17];
  assign t[4] = ~x[2] & t[21];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[25];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[20];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[16];
  assign t[56] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[57] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[58] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[59] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[5] = ~(t[6] & t[7]);
  assign t[60] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[63] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[64] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[65] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[66] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[67] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[68] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[69] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[6] = ~(t[22] & t[8]);
  assign t[7] = ~(t[23] & t[9]);
  assign t[8] = ~(t[24]);
  assign t[9] = ~(t[24] & t[10]);
  assign y = (t[0] & ~t[11]) | (~t[0] & t[11]);
endmodule

module R2ind124(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21]);
  assign t[11] = ~(t[12] ^ t[13]);
  assign t[12] = ~t[14];
  assign t[13] = t[4] ? x[23] : x[22];
  assign t[14] = x[2] ? x[24] : t[15];
  assign t[15] = ~(t[16] & t[17]);
  assign t[16] = ~(t[8] & t[18]);
  assign t[17] = t[19] | t[24];
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[10] | t[8]);
  assign t[1] = ~t[3];
  assign t[20] = (t[25] & ~t[26]) | (~t[25] & t[26]);
  assign t[21] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[22] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[23] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[24] = (t[27] & ~t[32]) | (~t[27] & t[32]);
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[18];
  assign t[29] = t[37] ^ x[19];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[20];
  assign t[31] = t[39] ^ x[21];
  assign t[32] = t[40] ^ x[25];
  assign t[33] = (t[41] & ~t[43] & ~t[44] & ~t[45] & ~t[46]) | (t[41] & ~t[42] & ~t[44] & ~t[45] & ~t[47]) | (t[41] & ~t[42] & ~t[43] & ~t[46] & ~t[47]) | (~t[41] & t[42] & t[43] & t[44] & ~t[47]) | (~t[41] & t[42] & t[45] & t[46] & ~t[47]) | (t[41] & ~t[43] & ~t[45] & t[47]) | (~t[41] & t[43] & t[45] & t[47]);
  assign t[34] = (t[41] & t[42] & ~t[43] & ~t[45] & t[46] & ~t[47]) | (t[41] & t[43] & ~t[44] & ~t[45] & ~t[46] & t[47]) | (~t[42] & ~t[43] & t[45] & ~t[46] & ~t[47]) | (~t[41] & ~t[43] & ~t[44] & t[45] & ~t[46]) | (~t[41] & ~t[42] & ~t[44] & t[45] & ~t[47]) | (~t[41] & ~t[43] & t[44] & t[45] & t[46]) | (t[44] & t[45] & ~t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[36] = (t[49] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & t[49] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[49] & ~t[50] & ~t[53] & ~t[54]) | (t[48] & ~t[49] & t[50] & t[51] & ~t[54]) | (t[48] & ~t[49] & t[52] & t[53] & ~t[54]) | (t[49] & ~t[51] & ~t[53] & t[54]) | (~t[49] & t[51] & t[53] & t[54]);
  assign t[37] = (t[48] & t[49] & t[50] & ~t[51] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & ~t[51] & ~t[52] & t[53] & t[54]) | (~t[49] & ~t[50] & t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[50] & t[51] & ~t[53] & ~t[54]) | (~t[48] & ~t[49] & t[51] & ~t[52] & ~t[54]) | (~t[49] & t[50] & t[51] & t[52] & ~t[53]) | (~t[50] & t[51] & t[52] & ~t[54]);
  assign t[38] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[39] = (t[48] & t[49] & ~t[51] & t[52] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & ~t[51] & ~t[52] & t[53]) | (~t[48] & ~t[51] & ~t[52] & t[53] & ~t[54]) | (~t[48] & ~t[49] & ~t[50] & t[53] & ~t[54]) | (~t[49] & t[50] & ~t[51] & t[52] & t[53]) | (t[50] & ~t[52] & t[53] & ~t[54]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[48] & t[49] & ~t[50] & t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[50] & ~t[51] & t[52] & ~t[53] & t[54]) | (~t[49] & t[50] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[49] & t[50] & ~t[53] & ~t[54]) | (~t[48] & t[50] & t[51] & ~t[52] & t[53]) | (t[50] & ~t[51] & t[53] & ~t[54]);
  assign t[41] = t[55] ^ x[10];
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[7];
  assign t[45] = t[59] ^ x[11];
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[17];
  assign t[49] = t[63] ^ x[18];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[64] ^ x[25];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[20];
  assign t[53] = t[67] ^ x[21];
  assign t[54] = t[68] ^ x[16];
  assign t[55] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[56] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[57] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[58] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[59] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[5] = ~(t[6] & t[7]);
  assign t[60] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[63] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[64] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[65] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[66] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[67] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[68] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[6] = ~(t[21] & t[8]);
  assign t[7] = ~(t[22] & t[9]);
  assign t[8] = ~(t[23]);
  assign t[9] = ~(t[23] & t[10]);
  assign y = (t[0] & ~t[11]) | (~t[0] & t[11]);
endmodule

module R2ind125(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[23] & t[22]);
  assign t[12] = ~(t[24]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[24] : x[23];
  assign t[16] = x[2] ? x[25] : t[17];
  assign t[17] = ~(t[6] & t[18]);
  assign t[18] = t[19] | t[21];
  assign t[19] = ~(t[12] | t[8]);
  assign t[1] = ~t[3];
  assign t[20] = (t[25] & ~t[26]) | (~t[25] & t[26]);
  assign t[21] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[22] = (t[27] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[27] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[23] = (t[27] & ~t[31]) | (~t[27] & t[31]);
  assign t[24] = (t[27] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[27] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[25] = t[33] ^ x[10];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[18];
  assign t[29] = t[37] ^ x[19];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[20];
  assign t[31] = t[39] ^ x[21];
  assign t[32] = t[40] ^ x[22];
  assign t[33] = (t[41] & ~t[43] & ~t[44] & ~t[45] & ~t[46]) | (t[41] & ~t[42] & ~t[44] & ~t[45] & ~t[47]) | (t[41] & ~t[42] & ~t[43] & ~t[46] & ~t[47]) | (~t[41] & t[42] & t[43] & t[44] & ~t[47]) | (~t[41] & t[42] & t[45] & t[46] & ~t[47]) | (t[41] & ~t[43] & ~t[45] & t[47]) | (~t[41] & t[43] & t[45] & t[47]);
  assign t[34] = (t[41] & t[42] & ~t[43] & ~t[45] & t[46] & ~t[47]) | (t[41] & t[43] & ~t[44] & ~t[45] & ~t[46] & t[47]) | (~t[42] & ~t[43] & t[45] & ~t[46] & ~t[47]) | (~t[41] & ~t[43] & ~t[44] & t[45] & ~t[46]) | (~t[41] & ~t[42] & ~t[44] & t[45] & ~t[47]) | (~t[41] & ~t[43] & t[44] & t[45] & t[46]) | (t[44] & t[45] & ~t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (t[48] & ~t[49] & ~t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[49] & ~t[50] & ~t[53] & ~t[54]) | (~t[48] & t[49] & t[50] & t[51] & ~t[54]) | (~t[48] & t[49] & t[52] & t[53] & ~t[54]) | (t[48] & ~t[50] & ~t[52] & t[54]) | (~t[48] & t[50] & t[52] & t[54]);
  assign t[36] = (t[48] & t[49] & ~t[50] & t[51] & ~t[52] & ~t[54]) | (t[48] & ~t[50] & ~t[51] & t[52] & ~t[53] & t[54]) | (~t[49] & t[50] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[49] & t[50] & ~t[53] & ~t[54]) | (~t[48] & t[50] & t[51] & ~t[52] & t[53]) | (t[50] & ~t[51] & t[53] & ~t[54]);
  assign t[37] = (t[49] & ~t[50] & ~t[51] & ~t[52] & ~t[53]) | (~t[48] & t[49] & ~t[51] & ~t[52] & ~t[54]) | (~t[48] & t[49] & ~t[50] & ~t[53] & ~t[54]) | (t[48] & ~t[49] & t[50] & t[51] & ~t[54]) | (t[48] & ~t[49] & t[52] & t[53] & ~t[54]) | (t[49] & ~t[51] & ~t[53] & t[54]) | (~t[49] & t[51] & t[53] & t[54]);
  assign t[38] = (t[48] & t[49] & t[50] & ~t[51] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & ~t[51] & ~t[52] & t[53] & t[54]) | (~t[49] & ~t[50] & t[51] & ~t[52] & ~t[53]) | (~t[48] & ~t[50] & t[51] & ~t[53] & ~t[54]) | (~t[48] & ~t[49] & t[51] & ~t[52] & ~t[54]) | (~t[49] & t[50] & t[51] & t[52] & ~t[53]) | (~t[50] & t[51] & t[52] & ~t[54]);
  assign t[39] = (t[48] & t[49] & ~t[50] & ~t[52] & t[53] & ~t[54]) | (t[48] & t[50] & ~t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & t[52] & ~t[53] & ~t[54]) | (~t[48] & ~t[50] & ~t[51] & t[52] & ~t[53]) | (~t[48] & ~t[49] & ~t[51] & t[52] & ~t[54]) | (~t[48] & ~t[50] & t[51] & t[52] & t[53]) | (t[51] & t[52] & ~t[53] & ~t[54]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[48] & t[49] & ~t[51] & t[52] & ~t[53] & ~t[54]) | (t[49] & ~t[50] & t[51] & ~t[52] & ~t[53] & t[54]) | (~t[49] & ~t[50] & ~t[51] & ~t[52] & t[53]) | (~t[48] & ~t[51] & ~t[52] & t[53] & ~t[54]) | (~t[48] & ~t[49] & ~t[50] & t[53] & ~t[54]) | (~t[49] & t[50] & ~t[51] & t[52] & t[53]) | (t[50] & ~t[52] & t[53] & ~t[54]);
  assign t[41] = t[55] ^ x[10];
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[7];
  assign t[45] = t[59] ^ x[11];
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[17];
  assign t[49] = t[63] ^ x[19];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[21];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[16];
  assign t[55] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[56] = (x[4] & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0);
  assign t[57] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[58] = (x[4] & ~1'b0) | (~x[4] & 1'b0);
  assign t[59] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[5] = ~(t[6] & t[7]);
  assign t[60] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[61] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[62] = (x[12] & ~x[13] & ~x[14]) | (~x[12] & x[13] & ~x[14]) | (~x[12] & ~x[13] & x[14]) | (x[12] & x[13] & x[14]);
  assign t[63] = (x[12] & ~x[13] & ~x[15]) | (~x[12] & x[13] & ~x[15]) | (~x[12] & ~x[13] & x[15]) | (x[12] & x[13] & x[15]);
  assign t[64] = (x[12] & ~x[14]) | (~x[12] & x[14]);
  assign t[65] = (x[12] & ~x[15]) | (~x[12] & x[15]);
  assign t[66] = (x[13] & ~x[14]) | (~x[13] & x[14]);
  assign t[67] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[68] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[21]);
  assign t[8] = ~(t[22]);
  assign t[9] = ~(t[23]);
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind126(x, y);
 input [28:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[35]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[36]);
  assign t[14] = ~(t[34] | t[35]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[34] & t[11]);
  assign t[21] = ~(t[36] & t[22]);
  assign t[22] = ~(t[35] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[36] & t[35]);
  assign t[32] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[33] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[34] = (t[37] & ~t[42] & ~t[44]) | (~t[41] & t[42] & ~t[43]) | (~t[37] & ~t[42] & t[44]) | (t[41] & t[42] & t[43]);
  assign t[35] = (t[37] & ~t[42] & ~t[43]) | (~t[41] & t[42] & ~t[44]) | (~t[37] & ~t[42] & t[43]) | (t[41] & t[42] & t[44]);
  assign t[36] = (t[37] & ~t[43]) | (~t[37] & t[43]);
  assign t[37] = t[45] ^ x[9];
  assign t[38] = t[46] ^ x[10];
  assign t[39] = t[47] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[18];
  assign t[41] = t[49] ^ x[19];
  assign t[42] = t[50] ^ x[20];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[22];
  assign t[45] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[46] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[8];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[12];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[15];
  assign t[66] = t[80] ^ x[16];
  assign t[67] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[68] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[69] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[71] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[72] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[73] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[75] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[76] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[77] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[79] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = ~(t[32] | t[12]);
  assign t[9] = ~x[2] & t[33];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind127(x, y);
 input [28:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[34]);
  assign t[14] = ~(t[32] | t[33]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32] & t[11]);
  assign t[21] = ~(t[34] & t[22]);
  assign t[22] = ~(t[33] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[27] : x[26];
  assign t[26] = x[2] ? x[28] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = t[7] | t[30];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[31] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[32] = (t[35] & ~t[40] & ~t[42]) | (~t[39] & t[40] & ~t[41]) | (~t[35] & ~t[40] & t[42]) | (t[39] & t[40] & t[41]);
  assign t[33] = (t[35] & ~t[40] & ~t[41]) | (~t[39] & t[40] & ~t[42]) | (~t[35] & ~t[40] & t[41]) | (t[39] & t[40] & t[42]);
  assign t[34] = (t[35] & ~t[41]) | (~t[35] & t[41]);
  assign t[35] = t[43] ^ x[9];
  assign t[36] = t[44] ^ x[10];
  assign t[37] = t[45] ^ x[17];
  assign t[38] = t[46] ^ x[18];
  assign t[39] = t[47] ^ x[19];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = t[48] ^ x[20];
  assign t[41] = t[49] ^ x[21];
  assign t[42] = t[50] ^ x[22];
  assign t[43] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[44] = (t[51] & t[52] & ~t[53] & t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[53] & ~t[54] & t[55] & ~t[56] & t[57]) | (~t[52] & t[53] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[52] & t[53] & ~t[56] & ~t[57]) | (~t[51] & t[53] & t[54] & ~t[55] & t[56]) | (t[53] & ~t[54] & t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[60] & ~t[61] & ~t[62] & ~t[63]) | (t[58] & ~t[59] & ~t[61] & ~t[62] & ~t[64]) | (t[58] & ~t[59] & ~t[60] & ~t[63] & ~t[64]) | (~t[58] & t[59] & t[60] & t[61] & ~t[64]) | (~t[58] & t[59] & t[62] & t[63] & ~t[64]) | (t[58] & ~t[60] & ~t[62] & t[64]) | (~t[58] & t[60] & t[62] & t[64]);
  assign t[46] = (t[58] & t[59] & ~t[60] & ~t[62] & t[63] & ~t[64]) | (t[58] & t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[64]) | (~t[58] & ~t[60] & ~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[59] & ~t[61] & t[62] & ~t[64]) | (~t[58] & ~t[60] & t[61] & t[62] & t[63]) | (t[61] & t[62] & ~t[63] & ~t[64]);
  assign t[47] = (t[52] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (~t[51] & t[52] & ~t[54] & ~t[55] & ~t[57]) | (~t[51] & t[52] & ~t[53] & ~t[56] & ~t[57]) | (t[51] & ~t[52] & t[53] & t[54] & ~t[57]) | (t[51] & ~t[52] & t[55] & t[56] & ~t[57]) | (t[52] & ~t[54] & ~t[56] & t[57]) | (~t[52] & t[54] & t[56] & t[57]);
  assign t[48] = (t[51] & t[52] & t[53] & ~t[54] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[54] & ~t[55] & t[56] & t[57]) | (~t[52] & ~t[53] & t[54] & ~t[55] & ~t[56]) | (~t[51] & ~t[53] & t[54] & ~t[56] & ~t[57]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[57]) | (~t[52] & t[53] & t[54] & t[55] & ~t[56]) | (~t[53] & t[54] & t[55] & ~t[57]);
  assign t[49] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[4] = ~(t[6]);
  assign t[50] = (t[51] & t[52] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[51] & ~t[52] & ~t[53] & t[56] & ~t[57]) | (~t[52] & t[53] & ~t[54] & t[55] & t[56]) | (t[53] & ~t[55] & t[56] & ~t[57]);
  assign t[51] = t[65] ^ x[9];
  assign t[52] = t[66] ^ x[19];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[8];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[12];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[66] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[67] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[68] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[69] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[71] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[74] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[75] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[76] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[77] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[78] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[30] | t[12]);
  assign t[9] = ~x[2] & t[31];
  assign y = (t[0] & ~t[15] & ~t[23]) | (~t[0] & t[15] & ~t[23]) | (~t[0] & ~t[15] & t[23]) | (t[0] & t[15] & t[23]);
endmodule

module R2ind128(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[28]);
  assign t[14] = ~(t[26] | t[27]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = ~(t[22] & t[24]);
  assign t[22] = ~(t[23] & t[10]);
  assign t[23] = ~(t[28] & t[27]);
  assign t[24] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[29] & ~t[34] & ~t[36]) | (~t[33] & t[34] & ~t[35]) | (~t[29] & ~t[34] & t[36]) | (t[33] & t[34] & t[35]);
  assign t[27] = (t[29] & ~t[34] & ~t[35]) | (~t[33] & t[34] & ~t[36]) | (~t[29] & ~t[34] & t[35]) | (t[33] & t[34] & t[36]);
  assign t[28] = (t[29] & ~t[35]) | (~t[29] & t[35]);
  assign t[29] = t[37] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[10];
  assign t[31] = t[39] ^ x[17];
  assign t[32] = t[40] ^ x[18];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[20];
  assign t[35] = t[43] ^ x[21];
  assign t[36] = t[44] ^ x[22];
  assign t[37] = (t[45] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[46] & ~t[47] & ~t[50] & ~t[51]) | (~t[45] & t[46] & t[47] & t[48] & ~t[51]) | (~t[45] & t[46] & t[49] & t[50] & ~t[51]) | (t[45] & ~t[47] & ~t[49] & t[51]) | (~t[45] & t[47] & t[49] & t[51]);
  assign t[38] = (t[45] & t[46] & ~t[47] & t[48] & ~t[49] & ~t[51]) | (t[45] & ~t[47] & ~t[48] & t[49] & ~t[50] & t[51]) | (~t[46] & t[47] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[46] & t[47] & ~t[50] & ~t[51]) | (~t[45] & t[47] & t[48] & ~t[49] & t[50]) | (t[47] & ~t[48] & t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[41] = (t[46] & ~t[47] & ~t[48] & ~t[49] & ~t[50]) | (~t[45] & t[46] & ~t[48] & ~t[49] & ~t[51]) | (~t[45] & t[46] & ~t[47] & ~t[50] & ~t[51]) | (t[45] & ~t[46] & t[47] & t[48] & ~t[51]) | (t[45] & ~t[46] & t[49] & t[50] & ~t[51]) | (t[46] & ~t[48] & ~t[50] & t[51]) | (~t[46] & t[48] & t[50] & t[51]);
  assign t[42] = (t[45] & t[46] & t[47] & ~t[48] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[48] & ~t[49] & t[50] & t[51]) | (~t[46] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (~t[45] & ~t[47] & t[48] & ~t[50] & ~t[51]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[51]) | (~t[46] & t[47] & t[48] & t[49] & ~t[50]) | (~t[47] & t[48] & t[49] & ~t[51]);
  assign t[43] = (t[45] & t[46] & ~t[47] & ~t[49] & t[50] & ~t[51]) | (t[45] & t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[51]) | (~t[45] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[45] & ~t[46] & ~t[48] & t[49] & ~t[51]) | (~t[45] & ~t[47] & t[48] & t[49] & t[50]) | (t[48] & t[49] & ~t[50] & ~t[51]);
  assign t[44] = (t[45] & t[46] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[45] & ~t[46] & ~t[47] & t[50] & ~t[51]) | (~t[46] & t[47] & ~t[48] & t[49] & t[50]) | (t[47] & ~t[49] & t[50] & ~t[51]);
  assign t[45] = t[59] ^ x[9];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[20];
  assign t[49] = t[63] ^ x[21];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[22];
  assign t[51] = t[65] ^ x[8];
  assign t[52] = t[66] ^ x[17];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[13];
  assign t[55] = t[69] ^ x[14];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[61] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[62] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[63] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[64] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[65] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[68] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[69] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[72] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[24] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind129(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[24] | t[25]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[11] & t[13]);
  assign t[21] = t[7] | t[22];
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[25] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[26] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[22] | t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind130(x, y);
 input [25:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = ~(t[26] & t[12]);
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = ~(t[21] & t[27]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[22] & t[12]);
  assign t[22] = ~(t[24] & t[26]);
  assign t[23] = (t[28] & ~t[30] & ~t[32]) | (~t[29] & t[30] & ~t[31]) | (~t[28] & ~t[30] & t[32]) | (t[29] & t[30] & t[31]);
  assign t[24] = (t[28] & ~t[31]) | (~t[28] & t[31]);
  assign t[25] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[26] = (t[28] & ~t[30] & ~t[31]) | (~t[29] & t[30] & ~t[32]) | (~t[28] & ~t[30] & t[31]) | (t[29] & t[30] & t[32]);
  assign t[27] = (t[28] & ~t[35]) | (~t[28] & t[35]);
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[13];
  assign t[33] = t[41] ^ x[20];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[45] & ~t[46] & ~t[49] & ~t[50]) | (~t[44] & t[45] & t[46] & t[47] & ~t[50]) | (~t[44] & t[45] & t[48] & t[49] & ~t[50]) | (t[44] & ~t[46] & ~t[48] & t[50]) | (~t[44] & t[46] & t[48] & t[50]);
  assign t[37] = (t[45] & ~t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & t[45] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[45] & ~t[46] & ~t[49] & ~t[50]) | (t[44] & ~t[45] & t[46] & t[47] & ~t[50]) | (t[44] & ~t[45] & t[48] & t[49] & ~t[50]) | (t[45] & ~t[47] & ~t[49] & t[50]) | (~t[45] & t[47] & t[49] & t[50]);
  assign t[38] = (t[44] & t[45] & t[46] & ~t[47] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & ~t[47] & ~t[48] & t[49] & t[50]) | (~t[45] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[46] & t[47] & ~t[49] & ~t[50]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[50]) | (~t[45] & t[46] & t[47] & t[48] & ~t[49]) | (~t[46] & t[47] & t[48] & ~t[50]);
  assign t[39] = (t[44] & t[45] & ~t[46] & ~t[48] & t[49] & ~t[50]) | (t[44] & t[46] & ~t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & t[48] & ~t[49] & ~t[50]) | (~t[44] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[44] & ~t[45] & ~t[47] & t[48] & ~t[50]) | (~t[44] & ~t[46] & t[47] & t[48] & t[49]) | (t[47] & t[48] & ~t[49] & ~t[50]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[44] & t[45] & ~t[47] & t[48] & ~t[49] & ~t[50]) | (t[45] & ~t[46] & t[47] & ~t[48] & ~t[49] & t[50]) | (~t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[47] & ~t[48] & t[49] & ~t[50]) | (~t[44] & ~t[45] & ~t[46] & t[49] & ~t[50]) | (~t[45] & t[46] & ~t[47] & t[48] & t[49]) | (t[46] & ~t[48] & t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[53] & ~t[54] & ~t[55] & ~t[56]) | (t[51] & ~t[52] & ~t[54] & ~t[55] & ~t[57]) | (t[51] & ~t[52] & ~t[53] & ~t[56] & ~t[57]) | (~t[51] & t[52] & t[53] & t[54] & ~t[57]) | (~t[51] & t[52] & t[55] & t[56] & ~t[57]) | (t[51] & ~t[53] & ~t[55] & t[57]) | (~t[51] & t[53] & t[55] & t[57]);
  assign t[42] = (t[51] & t[52] & ~t[53] & ~t[55] & t[56] & ~t[57]) | (t[51] & t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[57]) | (~t[51] & ~t[53] & ~t[54] & t[55] & ~t[56]) | (~t[51] & ~t[52] & ~t[54] & t[55] & ~t[57]) | (~t[51] & ~t[53] & t[54] & t[55] & t[56]) | (t[54] & t[55] & ~t[56] & ~t[57]);
  assign t[43] = (t[44] & t[45] & ~t[46] & t[47] & ~t[48] & ~t[50]) | (t[44] & ~t[46] & ~t[47] & t[48] & ~t[49] & t[50]) | (~t[45] & t[46] & ~t[47] & ~t[48] & ~t[50]) | (~t[44] & t[46] & ~t[47] & ~t[48] & ~t[49]) | (~t[44] & ~t[45] & t[46] & ~t[49] & ~t[50]) | (~t[44] & t[46] & t[47] & ~t[48] & t[49]) | (t[46] & ~t[47] & t[49] & ~t[50]);
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[25];
  assign t[47] = t[61] ^ x[11];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[13];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[8];
  assign t[51] = t[65] ^ x[20];
  assign t[52] = t[66] ^ x[15];
  assign t[53] = t[67] ^ x[16];
  assign t[54] = t[68] ^ x[17];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[19];
  assign t[58] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[59] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[61] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[62] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[63] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[64] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[71] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[23] & t[10]);
  assign t[8] = ~(t[24] & t[11]);
  assign t[9] = ~x[2] & t[25];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind131(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[25]);
  assign t[11] = ~(t[25] & t[12]);
  assign t[12] = ~(t[22]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[23] : x[22];
  assign t[16] = x[2] ? x[24] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[10] & t[20]);
  assign t[19] = t[21] | t[26];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[12] | t[10]);
  assign t[22] = (t[27] & ~t[29] & ~t[31]) | (~t[28] & t[29] & ~t[30]) | (~t[27] & ~t[29] & t[31]) | (t[28] & t[29] & t[30]);
  assign t[23] = (t[27] & ~t[30]) | (~t[27] & t[30]);
  assign t[24] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[25] = (t[27] & ~t[29] & ~t[30]) | (~t[28] & t[29] & ~t[31]) | (~t[27] & ~t[29] & t[30]) | (t[28] & t[29] & t[31]);
  assign t[26] = (t[27] & ~t[34]) | (~t[27] & t[34]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[12];
  assign t[31] = t[39] ^ x[13];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[25];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[37] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[38] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[39] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[41] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[42] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[10];
  assign t[45] = t[59] ^ x[25];
  assign t[46] = t[60] ^ x[11];
  assign t[47] = t[61] ^ x[12];
  assign t[48] = t[62] ^ x[13];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[20];
  assign t[51] = t[65] ^ x[15];
  assign t[52] = t[66] ^ x[16];
  assign t[53] = t[67] ^ x[17];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[18];
  assign t[56] = t[70] ^ x[19];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0);
  assign t[66] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[67] = (x[14] & ~1'b0) | (~x[14] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[22] & t[10]);
  assign t[8] = ~(t[23] & t[11]);
  assign t[9] = ~x[2] & t[24];
  assign y = (t[0] & ~t[13]) | (~t[0] & t[13]);
endmodule

module R2ind132(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = ~(t[25]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] & t[24]);
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[24] : x[23];
  assign t[18] = x[2] ? x[25] : t[19];
  assign t[19] = ~(t[7] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = t[21] | t[22];
  assign t[21] = ~(t[14] | t[10]);
  assign t[22] = (t[27] & ~t[28]) | (~t[27] & t[28]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[27] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[27] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[25] = (t[27] & ~t[33]) | (~t[27] & t[33]);
  assign t[26] = (t[27] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[27] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[10];
  assign t[29] = t[37] ^ x[17];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[18];
  assign t[31] = t[39] ^ x[19];
  assign t[32] = t[40] ^ x[20];
  assign t[33] = t[41] ^ x[21];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[36] = (t[43] & t[44] & ~t[45] & t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[45] & ~t[46] & t[47] & ~t[48] & t[49]) | (~t[44] & t[45] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[44] & t[45] & ~t[48] & ~t[49]) | (~t[43] & t[45] & t[46] & ~t[47] & t[48]) | (t[45] & ~t[46] & t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[38] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[39] = (t[44] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (~t[43] & t[44] & ~t[46] & ~t[47] & ~t[49]) | (~t[43] & t[44] & ~t[45] & ~t[48] & ~t[49]) | (t[43] & ~t[44] & t[45] & t[46] & ~t[49]) | (t[43] & ~t[44] & t[47] & t[48] & ~t[49]) | (t[44] & ~t[46] & ~t[48] & t[49]) | (~t[44] & t[46] & t[48] & t[49]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[43] & t[44] & t[45] & ~t[46] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & ~t[46] & ~t[47] & t[48] & t[49]) | (~t[44] & ~t[45] & t[46] & ~t[47] & ~t[48]) | (~t[43] & ~t[45] & t[46] & ~t[48] & ~t[49]) | (~t[43] & ~t[44] & t[46] & ~t[47] & ~t[49]) | (~t[44] & t[45] & t[46] & t[47] & ~t[48]) | (~t[45] & t[46] & t[47] & ~t[49]);
  assign t[41] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[42] = (t[43] & t[44] & ~t[46] & t[47] & ~t[48] & ~t[49]) | (t[44] & ~t[45] & t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & ~t[46] & ~t[47] & t[48]) | (~t[43] & ~t[46] & ~t[47] & t[48] & ~t[49]) | (~t[43] & ~t[44] & ~t[45] & t[48] & ~t[49]) | (~t[44] & t[45] & ~t[46] & t[47] & t[48]) | (t[45] & ~t[47] & t[48] & ~t[49]);
  assign t[43] = t[57] ^ x[9];
  assign t[44] = t[58] ^ x[19];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = t[62] ^ x[22];
  assign t[49] = t[63] ^ x[8];
  assign t[4] = ~(t[6]);
  assign t[50] = t[64] ^ x[17];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[13];
  assign t[53] = t[67] ^ x[14];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[15];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = (x[4] & ~x[5] & ~x[6]) | (~x[4] & x[5] & ~x[6]) | (~x[4] & ~x[5] & x[6]) | (x[4] & x[5] & x[6]);
  assign t[58] = (x[4] & ~x[5] & ~x[7]) | (~x[4] & x[5] & ~x[7]) | (~x[4] & ~x[5] & x[7]) | (x[4] & x[5] & x[7]);
  assign t[59] = (x[4] & ~x[6]) | (~x[4] & x[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~x[7]) | (~x[4] & x[7]);
  assign t[61] = (x[5] & ~x[6]) | (~x[5] & x[6]);
  assign t[62] = (x[5] & ~x[7]) | (~x[5] & x[7]);
  assign t[63] = (x[6] & ~x[7]) | (~x[6] & x[7]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0);
  assign t[66] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[67] = (x[11] & ~1'b0) | (~x[11] & 1'b0);
  assign t[68] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[69] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[6] = ~(t[9]);
  assign t[70] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[22]);
  assign t[9] = ~x[2] & t[23];
  assign y = (t[0] & ~t[15]) | (~t[0] & t[15]);
endmodule

module R2ind133(x, y);
 input [42:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[121] ^ x[9];
  assign t[101] = t[122] ^ x[10];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[27];
  assign t[104] = t[125] ^ x[19];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[29];
  assign t[107] = t[128] ^ x[30];
  assign t[108] = t[129] ^ x[17];
  assign t[109] = t[130] ^ x[25];
  assign t[10] = ~x[2] & t[58];
  assign t[110] = t[131] ^ x[31];
  assign t[111] = t[132] ^ x[26];
  assign t[112] = t[133] ^ x[32];
  assign t[113] = t[134] ^ x[33];
  assign t[114] = t[135] ^ x[34];
  assign t[115] = t[136] ^ x[24];
  assign t[116] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[117] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[118] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[119] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[11] = ~(t[14] | t[15]);
  assign t[120] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[121] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[124] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[125] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[126] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[127] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[128] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[129] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[131] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[132] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[133] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[134] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[135] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[136] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = ~(t[59] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[60] | t[21]);
  assign t[16] = ~(t[61]);
  assign t[17] = ~(t[62]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[63]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[64]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[65]);
  assign t[23] = ~(t[61] | t[62]);
  assign t[24] = ~(t[66]);
  assign t[25] = ~(t[63] | t[64]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[10] ? x[36] : x[35];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[37] : t[33];
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[61] & t[17]);
  assign t[36] = ~(t[65] & t[39]);
  assign t[37] = ~(t[63] & t[20]);
  assign t[38] = ~(t[66] & t[40]);
  assign t[39] = ~(t[62] & t[16]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[64] & t[19]);
  assign t[41] = ~(t[42] ^ t[43]);
  assign t[42] = ~t[44];
  assign t[43] = t[4] ? x[40] : x[39];
  assign t[44] = ~(t[45] ^ t[46]);
  assign t[45] = ~t[47];
  assign t[46] = x[2] ? x[41] : t[48];
  assign t[47] = x[2] ? x[42] : t[49];
  assign t[48] = ~(t[50] & t[51]);
  assign t[49] = ~(t[52] & t[53]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[17] & t[22]);
  assign t[51] = ~(t[54] & t[59]);
  assign t[52] = ~(t[20] & t[24]);
  assign t[53] = ~(t[55] & t[60]);
  assign t[54] = ~(t[56] & t[16]);
  assign t[55] = ~(t[57] & t[19]);
  assign t[56] = ~(t[65] & t[62]);
  assign t[57] = ~(t[66] & t[64]);
  assign t[58] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[59] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[5] = ~t[8];
  assign t[60] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[61] = (t[69] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[69] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[62] = (t[69] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[69] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[63] = (t[71] & ~t[78] & ~t[80]) | (~t[77] & t[78] & ~t[79]) | (~t[71] & ~t[78] & t[80]) | (t[77] & t[78] & t[79]);
  assign t[64] = (t[71] & ~t[78] & ~t[79]) | (~t[77] & t[78] & ~t[80]) | (~t[71] & ~t[78] & t[79]) | (t[77] & t[78] & t[80]);
  assign t[65] = (t[69] & ~t[75]) | (~t[69] & t[75]);
  assign t[66] = (t[71] & ~t[79]) | (~t[71] & t[79]);
  assign t[67] = t[81] ^ x[11];
  assign t[68] = t[82] ^ x[12];
  assign t[69] = t[83] ^ x[18];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[84] ^ x[19];
  assign t[71] = t[85] ^ x[25];
  assign t[72] = t[86] ^ x[26];
  assign t[73] = t[87] ^ x[27];
  assign t[74] = t[88] ^ x[28];
  assign t[75] = t[89] ^ x[29];
  assign t[76] = t[90] ^ x[30];
  assign t[77] = t[91] ^ x[31];
  assign t[78] = t[92] ^ x[32];
  assign t[79] = t[93] ^ x[33];
  assign t[7] = ~(t[10]);
  assign t[80] = t[94] ^ x[34];
  assign t[81] = (t[95] & ~t[97] & ~t[98] & ~t[99] & ~t[100]) | (t[95] & ~t[96] & ~t[98] & ~t[99] & ~t[101]) | (t[95] & ~t[96] & ~t[97] & ~t[100] & ~t[101]) | (~t[95] & t[96] & t[97] & t[98] & ~t[101]) | (~t[95] & t[96] & t[99] & t[100] & ~t[101]) | (t[95] & ~t[97] & ~t[99] & t[101]) | (~t[95] & t[97] & t[99] & t[101]);
  assign t[82] = (t[95] & t[96] & ~t[97] & ~t[99] & t[100] & ~t[101]) | (t[95] & t[97] & ~t[98] & ~t[99] & ~t[100] & t[101]) | (~t[96] & ~t[97] & t[99] & ~t[100] & ~t[101]) | (~t[95] & ~t[97] & ~t[98] & t[99] & ~t[100]) | (~t[95] & ~t[96] & ~t[98] & t[99] & ~t[101]) | (~t[95] & ~t[97] & t[98] & t[99] & t[100]) | (t[98] & t[99] & ~t[100] & ~t[101]);
  assign t[83] = (t[102] & ~t[104] & ~t[105] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & ~t[105] & ~t[106] & ~t[108]) | (t[102] & ~t[103] & ~t[104] & ~t[107] & ~t[108]) | (~t[102] & t[103] & t[104] & t[105] & ~t[108]) | (~t[102] & t[103] & t[106] & t[107] & ~t[108]) | (t[102] & ~t[104] & ~t[106] & t[108]) | (~t[102] & t[104] & t[106] & t[108]);
  assign t[84] = (t[102] & t[103] & ~t[104] & t[105] & ~t[106] & ~t[108]) | (t[102] & ~t[104] & ~t[105] & t[106] & ~t[107] & t[108]) | (~t[103] & t[104] & ~t[105] & ~t[106] & ~t[108]) | (~t[102] & t[104] & ~t[105] & ~t[106] & ~t[107]) | (~t[102] & ~t[103] & t[104] & ~t[107] & ~t[108]) | (~t[102] & t[104] & t[105] & ~t[106] & t[107]) | (t[104] & ~t[105] & t[107] & ~t[108]);
  assign t[85] = (t[109] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[110] & ~t[111] & ~t[114] & ~t[115]) | (~t[109] & t[110] & t[111] & t[112] & ~t[115]) | (~t[109] & t[110] & t[113] & t[114] & ~t[115]) | (t[109] & ~t[111] & ~t[113] & t[115]) | (~t[109] & t[111] & t[113] & t[115]);
  assign t[86] = (t[109] & t[110] & ~t[111] & t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[111] & ~t[112] & t[113] & ~t[114] & t[115]) | (~t[110] & t[111] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[110] & t[111] & ~t[114] & ~t[115]) | (~t[109] & t[111] & t[112] & ~t[113] & t[114]) | (t[111] & ~t[112] & t[114] & ~t[115]);
  assign t[87] = (t[103] & ~t[104] & ~t[105] & ~t[106] & ~t[107]) | (~t[102] & t[103] & ~t[105] & ~t[106] & ~t[108]) | (~t[102] & t[103] & ~t[104] & ~t[107] & ~t[108]) | (t[102] & ~t[103] & t[104] & t[105] & ~t[108]) | (t[102] & ~t[103] & t[106] & t[107] & ~t[108]) | (t[103] & ~t[105] & ~t[107] & t[108]) | (~t[103] & t[105] & t[107] & t[108]);
  assign t[88] = (t[102] & t[103] & t[104] & ~t[105] & ~t[107] & ~t[108]) | (t[103] & ~t[104] & ~t[105] & ~t[106] & t[107] & t[108]) | (~t[103] & ~t[104] & t[105] & ~t[106] & ~t[107]) | (~t[102] & ~t[104] & t[105] & ~t[107] & ~t[108]) | (~t[102] & ~t[103] & t[105] & ~t[106] & ~t[108]) | (~t[103] & t[104] & t[105] & t[106] & ~t[107]) | (~t[104] & t[105] & t[106] & ~t[108]);
  assign t[89] = (t[102] & t[103] & ~t[104] & ~t[106] & t[107] & ~t[108]) | (t[102] & t[104] & ~t[105] & ~t[106] & ~t[107] & t[108]) | (~t[103] & ~t[104] & t[106] & ~t[107] & ~t[108]) | (~t[102] & ~t[104] & ~t[105] & t[106] & ~t[107]) | (~t[102] & ~t[103] & ~t[105] & t[106] & ~t[108]) | (~t[102] & ~t[104] & t[105] & t[106] & t[107]) | (t[105] & t[106] & ~t[107] & ~t[108]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = (t[102] & t[103] & ~t[105] & t[106] & ~t[107] & ~t[108]) | (t[103] & ~t[104] & t[105] & ~t[106] & ~t[107] & t[108]) | (~t[103] & ~t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[105] & ~t[106] & t[107] & ~t[108]) | (~t[102] & ~t[103] & ~t[104] & t[107] & ~t[108]) | (~t[103] & t[104] & ~t[105] & t[106] & t[107]) | (t[104] & ~t[106] & t[107] & ~t[108]);
  assign t[91] = (t[110] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & t[110] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[110] & ~t[111] & ~t[114] & ~t[115]) | (t[109] & ~t[110] & t[111] & t[112] & ~t[115]) | (t[109] & ~t[110] & t[113] & t[114] & ~t[115]) | (t[110] & ~t[112] & ~t[114] & t[115]) | (~t[110] & t[112] & t[114] & t[115]);
  assign t[92] = (t[109] & t[110] & t[111] & ~t[112] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[112] & ~t[113] & t[114] & t[115]) | (~t[110] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[111] & t[112] & ~t[114] & ~t[115]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[115]) | (~t[110] & t[111] & t[112] & t[113] & ~t[114]) | (~t[111] & t[112] & t[113] & ~t[115]);
  assign t[93] = (t[109] & t[110] & ~t[111] & ~t[113] & t[114] & ~t[115]) | (t[109] & t[111] & ~t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & t[113] & ~t[114] & ~t[115]) | (~t[109] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[109] & ~t[110] & ~t[112] & t[113] & ~t[115]) | (~t[109] & ~t[111] & t[112] & t[113] & t[114]) | (t[112] & t[113] & ~t[114] & ~t[115]);
  assign t[94] = (t[109] & t[110] & ~t[112] & t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[109] & ~t[110] & ~t[111] & t[114] & ~t[115]) | (~t[110] & t[111] & ~t[112] & t[113] & t[114]) | (t[111] & ~t[113] & t[114] & ~t[115]);
  assign t[95] = t[116] ^ x[11];
  assign t[96] = t[117] ^ x[6];
  assign t[97] = t[118] ^ x[7];
  assign t[98] = t[119] ^ x[8];
  assign t[99] = t[120] ^ x[12];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[26] & ~t[41]) | (~t[0] & t[26] & ~t[41]) | (~t[0] & ~t[26] & t[41]) | (t[0] & t[26] & t[41]);
endmodule

module R2ind134(x, y);
 input [42:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[121] ^ x[19];
  assign t[101] = t[122] ^ x[28];
  assign t[102] = t[123] ^ x[29];
  assign t[103] = t[124] ^ x[30];
  assign t[104] = t[125] ^ x[17];
  assign t[105] = t[126] ^ x[25];
  assign t[106] = t[127] ^ x[31];
  assign t[107] = t[128] ^ x[26];
  assign t[108] = t[129] ^ x[32];
  assign t[109] = t[130] ^ x[33];
  assign t[10] = ~x[2] & t[54];
  assign t[110] = t[131] ^ x[34];
  assign t[111] = t[132] ^ x[24];
  assign t[112] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[113] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[114] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[115] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[120] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[121] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[122] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[123] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[124] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[125] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[126] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[127] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[128] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[129] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[131] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[132] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = ~(t[55] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[56] | t[21]);
  assign t[16] = ~(t[57]);
  assign t[17] = ~(t[58]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[59]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[60]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[61]);
  assign t[23] = ~(t[57] | t[58]);
  assign t[24] = ~(t[62]);
  assign t[25] = ~(t[59] | t[60]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[10] ? x[36] : x[35];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[37] : t[33];
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[57] & t[17]);
  assign t[36] = ~(t[61] & t[39]);
  assign t[37] = ~(t[59] & t[20]);
  assign t[38] = ~(t[62] & t[40]);
  assign t[39] = ~(t[58] & t[16]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[60] & t[19]);
  assign t[41] = ~(t[42] ^ t[43]);
  assign t[42] = ~t[44];
  assign t[43] = t[4] ? x[40] : x[39];
  assign t[44] = ~(t[45] ^ t[46]);
  assign t[45] = ~t[47];
  assign t[46] = x[2] ? x[41] : t[48];
  assign t[47] = x[2] ? x[42] : t[49];
  assign t[48] = ~(t[50] & t[51]);
  assign t[49] = ~(t[52] & t[53]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[17] & t[22]);
  assign t[51] = t[12] | t[55];
  assign t[52] = ~(t[20] & t[24]);
  assign t[53] = t[14] | t[56];
  assign t[54] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[55] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[56] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[57] = (t[65] & ~t[70] & ~t[72]) | (~t[69] & t[70] & ~t[71]) | (~t[65] & ~t[70] & t[72]) | (t[69] & t[70] & t[71]);
  assign t[58] = (t[65] & ~t[70] & ~t[71]) | (~t[69] & t[70] & ~t[72]) | (~t[65] & ~t[70] & t[71]) | (t[69] & t[70] & t[72]);
  assign t[59] = (t[67] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[67] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[5] = ~t[8];
  assign t[60] = (t[67] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[67] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[61] = (t[65] & ~t[71]) | (~t[65] & t[71]);
  assign t[62] = (t[67] & ~t[75]) | (~t[67] & t[75]);
  assign t[63] = t[77] ^ x[11];
  assign t[64] = t[78] ^ x[12];
  assign t[65] = t[79] ^ x[18];
  assign t[66] = t[80] ^ x[19];
  assign t[67] = t[81] ^ x[25];
  assign t[68] = t[82] ^ x[26];
  assign t[69] = t[83] ^ x[27];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[84] ^ x[28];
  assign t[71] = t[85] ^ x[29];
  assign t[72] = t[86] ^ x[30];
  assign t[73] = t[87] ^ x[31];
  assign t[74] = t[88] ^ x[32];
  assign t[75] = t[89] ^ x[33];
  assign t[76] = t[90] ^ x[34];
  assign t[77] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[78] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[79] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[7] = ~(t[10]);
  assign t[80] = (t[98] & t[99] & ~t[100] & t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[100] & ~t[101] & t[102] & ~t[103] & t[104]) | (~t[99] & t[100] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[99] & t[100] & ~t[103] & ~t[104]) | (~t[98] & t[100] & t[101] & ~t[102] & t[103]) | (t[100] & ~t[101] & t[103] & ~t[104]);
  assign t[81] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[82] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[83] = (t[99] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & t[99] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[99] & ~t[100] & ~t[103] & ~t[104]) | (t[98] & ~t[99] & t[100] & t[101] & ~t[104]) | (t[98] & ~t[99] & t[102] & t[103] & ~t[104]) | (t[99] & ~t[101] & ~t[103] & t[104]) | (~t[99] & t[101] & t[103] & t[104]);
  assign t[84] = (t[98] & t[99] & t[100] & ~t[101] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[101] & ~t[102] & t[103] & t[104]) | (~t[99] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[100] & t[101] & ~t[103] & ~t[104]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[104]) | (~t[99] & t[100] & t[101] & t[102] & ~t[103]) | (~t[100] & t[101] & t[102] & ~t[104]);
  assign t[85] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[86] = (t[98] & t[99] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[98] & ~t[99] & ~t[100] & t[103] & ~t[104]) | (~t[99] & t[100] & ~t[101] & t[102] & t[103]) | (t[100] & ~t[102] & t[103] & ~t[104]);
  assign t[87] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[88] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[89] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[91] = t[112] ^ x[11];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[7];
  assign t[94] = t[115] ^ x[8];
  assign t[95] = t[116] ^ x[12];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[10];
  assign t[98] = t[119] ^ x[18];
  assign t[99] = t[120] ^ x[27];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[26] & ~t[41]) | (~t[0] & t[26] & ~t[41]) | (~t[0] & ~t[26] & t[41]) | (t[0] & t[26] & t[41]);
endmodule

module R2ind135(x, y);
 input [38:0] x;
 output y;

 wire [121:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[121] ^ x[24];
  assign t[101] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[102] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[103] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[104] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[107] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[108] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[109] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[10] = ~x[2] & t[43];
  assign t[110] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[111] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[112] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[113] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[114] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[115] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[116] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[117] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[118] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[119] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[120] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[121] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[44] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[45] | t[21]);
  assign t[16] = ~(t[46]);
  assign t[17] = ~(t[47]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[48]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[49]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[50]);
  assign t[23] = ~(t[46] | t[47]);
  assign t[24] = ~(t[51]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[4] ? x[36] : x[35];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[37] : t[33];
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[17] & t[22]);
  assign t[36] = ~(t[39] & t[44]);
  assign t[37] = ~(t[20] & t[24]);
  assign t[38] = ~(t[40] & t[45]);
  assign t[39] = ~(t[41] & t[16]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[42] & t[19]);
  assign t[41] = ~(t[50] & t[47]);
  assign t[42] = ~(t[51] & t[49]);
  assign t[43] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[44] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[54] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[54] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[47] = (t[54] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[54] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[48] = (t[56] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[56] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[49] = (t[56] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[56] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[54] & ~t[60]) | (~t[54] & t[60]);
  assign t[51] = (t[56] & ~t[64]) | (~t[56] & t[64]);
  assign t[52] = t[66] ^ x[11];
  assign t[53] = t[67] ^ x[12];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[19];
  assign t[56] = t[70] ^ x[25];
  assign t[57] = t[71] ^ x[26];
  assign t[58] = t[72] ^ x[27];
  assign t[59] = t[73] ^ x[28];
  assign t[5] = ~t[8];
  assign t[60] = t[74] ^ x[29];
  assign t[61] = t[75] ^ x[30];
  assign t[62] = t[76] ^ x[31];
  assign t[63] = t[77] ^ x[32];
  assign t[64] = t[78] ^ x[33];
  assign t[65] = t[79] ^ x[34];
  assign t[66] = (t[80] & ~t[82] & ~t[83] & ~t[84] & ~t[85]) | (t[80] & ~t[81] & ~t[83] & ~t[84] & ~t[86]) | (t[80] & ~t[81] & ~t[82] & ~t[85] & ~t[86]) | (~t[80] & t[81] & t[82] & t[83] & ~t[86]) | (~t[80] & t[81] & t[84] & t[85] & ~t[86]) | (t[80] & ~t[82] & ~t[84] & t[86]) | (~t[80] & t[82] & t[84] & t[86]);
  assign t[67] = (t[80] & t[81] & ~t[82] & ~t[84] & t[85] & ~t[86]) | (t[80] & t[82] & ~t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[82] & t[84] & ~t[85] & ~t[86]) | (~t[80] & ~t[82] & ~t[83] & t[84] & ~t[85]) | (~t[80] & ~t[81] & ~t[83] & t[84] & ~t[86]) | (~t[80] & ~t[82] & t[83] & t[84] & t[85]) | (t[83] & t[84] & ~t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[89] & ~t[90] & ~t[91] & ~t[92]) | (t[87] & ~t[88] & ~t[90] & ~t[91] & ~t[93]) | (t[87] & ~t[88] & ~t[89] & ~t[92] & ~t[93]) | (~t[87] & t[88] & t[89] & t[90] & ~t[93]) | (~t[87] & t[88] & t[91] & t[92] & ~t[93]) | (t[87] & ~t[89] & ~t[91] & t[93]) | (~t[87] & t[89] & t[91] & t[93]);
  assign t[69] = (t[87] & t[88] & ~t[89] & t[90] & ~t[91] & ~t[93]) | (t[87] & ~t[89] & ~t[90] & t[91] & ~t[92] & t[93]) | (~t[88] & t[89] & ~t[90] & ~t[91] & ~t[93]) | (~t[87] & t[89] & ~t[90] & ~t[91] & ~t[92]) | (~t[87] & ~t[88] & t[89] & ~t[92] & ~t[93]) | (~t[87] & t[89] & t[90] & ~t[91] & t[92]) | (t[89] & ~t[90] & t[92] & ~t[93]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[94] & ~t[96] & ~t[97] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & ~t[97] & ~t[98] & ~t[100]) | (t[94] & ~t[95] & ~t[96] & ~t[99] & ~t[100]) | (~t[94] & t[95] & t[96] & t[97] & ~t[100]) | (~t[94] & t[95] & t[98] & t[99] & ~t[100]) | (t[94] & ~t[96] & ~t[98] & t[100]) | (~t[94] & t[96] & t[98] & t[100]);
  assign t[71] = (t[94] & t[95] & ~t[96] & t[97] & ~t[98] & ~t[100]) | (t[94] & ~t[96] & ~t[97] & t[98] & ~t[99] & t[100]) | (~t[95] & t[96] & ~t[97] & ~t[98] & ~t[100]) | (~t[94] & t[96] & ~t[97] & ~t[98] & ~t[99]) | (~t[94] & ~t[95] & t[96] & ~t[99] & ~t[100]) | (~t[94] & t[96] & t[97] & ~t[98] & t[99]) | (t[96] & ~t[97] & t[99] & ~t[100]);
  assign t[72] = (t[88] & ~t[89] & ~t[90] & ~t[91] & ~t[92]) | (~t[87] & t[88] & ~t[90] & ~t[91] & ~t[93]) | (~t[87] & t[88] & ~t[89] & ~t[92] & ~t[93]) | (t[87] & ~t[88] & t[89] & t[90] & ~t[93]) | (t[87] & ~t[88] & t[91] & t[92] & ~t[93]) | (t[88] & ~t[90] & ~t[92] & t[93]) | (~t[88] & t[90] & t[92] & t[93]);
  assign t[73] = (t[87] & t[88] & t[89] & ~t[90] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & ~t[90] & ~t[91] & t[92] & t[93]) | (~t[88] & ~t[89] & t[90] & ~t[91] & ~t[92]) | (~t[87] & ~t[89] & t[90] & ~t[92] & ~t[93]) | (~t[87] & ~t[88] & t[90] & ~t[91] & ~t[93]) | (~t[88] & t[89] & t[90] & t[91] & ~t[92]) | (~t[89] & t[90] & t[91] & ~t[93]);
  assign t[74] = (t[87] & t[88] & ~t[89] & ~t[91] & t[92] & ~t[93]) | (t[87] & t[89] & ~t[90] & ~t[91] & ~t[92] & t[93]) | (~t[88] & ~t[89] & t[91] & ~t[92] & ~t[93]) | (~t[87] & ~t[89] & ~t[90] & t[91] & ~t[92]) | (~t[87] & ~t[88] & ~t[90] & t[91] & ~t[93]) | (~t[87] & ~t[89] & t[90] & t[91] & t[92]) | (t[90] & t[91] & ~t[92] & ~t[93]);
  assign t[75] = (t[87] & t[88] & ~t[90] & t[91] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & t[90] & ~t[91] & ~t[92] & t[93]) | (~t[88] & ~t[89] & ~t[90] & ~t[91] & t[92]) | (~t[87] & ~t[90] & ~t[91] & t[92] & ~t[93]) | (~t[87] & ~t[88] & ~t[89] & t[92] & ~t[93]) | (~t[88] & t[89] & ~t[90] & t[91] & t[92]) | (t[89] & ~t[91] & t[92] & ~t[93]);
  assign t[76] = (t[95] & ~t[96] & ~t[97] & ~t[98] & ~t[99]) | (~t[94] & t[95] & ~t[97] & ~t[98] & ~t[100]) | (~t[94] & t[95] & ~t[96] & ~t[99] & ~t[100]) | (t[94] & ~t[95] & t[96] & t[97] & ~t[100]) | (t[94] & ~t[95] & t[98] & t[99] & ~t[100]) | (t[95] & ~t[97] & ~t[99] & t[100]) | (~t[95] & t[97] & t[99] & t[100]);
  assign t[77] = (t[94] & t[95] & t[96] & ~t[97] & ~t[99] & ~t[100]) | (t[95] & ~t[96] & ~t[97] & ~t[98] & t[99] & t[100]) | (~t[95] & ~t[96] & t[97] & ~t[98] & ~t[99]) | (~t[94] & ~t[96] & t[97] & ~t[99] & ~t[100]) | (~t[94] & ~t[95] & t[97] & ~t[98] & ~t[100]) | (~t[95] & t[96] & t[97] & t[98] & ~t[99]) | (~t[96] & t[97] & t[98] & ~t[100]);
  assign t[78] = (t[94] & t[95] & ~t[96] & ~t[98] & t[99] & ~t[100]) | (t[94] & t[96] & ~t[97] & ~t[98] & ~t[99] & t[100]) | (~t[95] & ~t[96] & t[98] & ~t[99] & ~t[100]) | (~t[94] & ~t[96] & ~t[97] & t[98] & ~t[99]) | (~t[94] & ~t[95] & ~t[97] & t[98] & ~t[100]) | (~t[94] & ~t[96] & t[97] & t[98] & t[99]) | (t[97] & t[98] & ~t[99] & ~t[100]);
  assign t[79] = (t[94] & t[95] & ~t[97] & t[98] & ~t[99] & ~t[100]) | (t[95] & ~t[96] & t[97] & ~t[98] & ~t[99] & t[100]) | (~t[95] & ~t[96] & ~t[97] & ~t[98] & t[99]) | (~t[94] & ~t[97] & ~t[98] & t[99] & ~t[100]) | (~t[94] & ~t[95] & ~t[96] & t[99] & ~t[100]) | (~t[95] & t[96] & ~t[97] & t[98] & t[99]) | (t[96] & ~t[98] & t[99] & ~t[100]);
  assign t[7] = ~(t[10]);
  assign t[80] = t[101] ^ x[11];
  assign t[81] = t[102] ^ x[6];
  assign t[82] = t[103] ^ x[7];
  assign t[83] = t[104] ^ x[8];
  assign t[84] = t[105] ^ x[12];
  assign t[85] = t[106] ^ x[9];
  assign t[86] = t[107] ^ x[10];
  assign t[87] = t[108] ^ x[18];
  assign t[88] = t[109] ^ x[27];
  assign t[89] = t[110] ^ x[19];
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = t[111] ^ x[28];
  assign t[91] = t[112] ^ x[29];
  assign t[92] = t[113] ^ x[30];
  assign t[93] = t[114] ^ x[17];
  assign t[94] = t[115] ^ x[25];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[26];
  assign t[97] = t[118] ^ x[32];
  assign t[98] = t[119] ^ x[33];
  assign t[99] = t[120] ^ x[34];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[26]) | (~t[0] & t[26]);
endmodule

module R2ind136(x, y);
 input [38:0] x;
 output y;

 wire [117:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[105] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[106] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[107] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[108] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[109] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[10] = ~x[2] & t[39];
  assign t[110] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[111] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[112] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[113] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[114] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[115] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[116] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[117] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[40] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[41] | t[21]);
  assign t[16] = ~(t[42]);
  assign t[17] = ~(t[43]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[44]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[45]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[46]);
  assign t[23] = ~(t[42] | t[43]);
  assign t[24] = ~(t[47]);
  assign t[25] = ~(t[44] | t[45]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[4] ? x[36] : x[35];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[37] : t[33];
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[17] & t[22]);
  assign t[36] = t[12] | t[40];
  assign t[37] = ~(t[20] & t[24]);
  assign t[38] = t[14] | t[41];
  assign t[39] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[41] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[42] = (t[50] & ~t[55] & ~t[57]) | (~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[55] & t[57]) | (t[54] & t[55] & t[56]);
  assign t[43] = (t[50] & ~t[55] & ~t[56]) | (~t[54] & t[55] & ~t[57]) | (~t[50] & ~t[55] & t[56]) | (t[54] & t[55] & t[57]);
  assign t[44] = (t[52] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[52] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[45] = (t[52] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[52] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[46] = (t[50] & ~t[56]) | (~t[50] & t[56]);
  assign t[47] = (t[52] & ~t[60]) | (~t[52] & t[60]);
  assign t[48] = t[62] ^ x[11];
  assign t[49] = t[63] ^ x[12];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[25];
  assign t[53] = t[67] ^ x[26];
  assign t[54] = t[68] ^ x[27];
  assign t[55] = t[69] ^ x[28];
  assign t[56] = t[70] ^ x[29];
  assign t[57] = t[71] ^ x[30];
  assign t[58] = t[72] ^ x[31];
  assign t[59] = t[73] ^ x[32];
  assign t[5] = ~t[8];
  assign t[60] = t[74] ^ x[33];
  assign t[61] = t[75] ^ x[34];
  assign t[62] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[63] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[65] = (t[83] & t[84] & ~t[85] & t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[85] & ~t[86] & t[87] & ~t[88] & t[89]) | (~t[84] & t[85] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[84] & t[85] & ~t[88] & ~t[89]) | (~t[83] & t[85] & t[86] & ~t[87] & t[88]) | (t[85] & ~t[86] & t[88] & ~t[89]);
  assign t[66] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[67] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[68] = (t[84] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & t[84] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[84] & ~t[85] & ~t[88] & ~t[89]) | (t[83] & ~t[84] & t[85] & t[86] & ~t[89]) | (t[83] & ~t[84] & t[87] & t[88] & ~t[89]) | (t[84] & ~t[86] & ~t[88] & t[89]) | (~t[84] & t[86] & t[88] & t[89]);
  assign t[69] = (t[83] & t[84] & t[85] & ~t[86] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[86] & ~t[87] & t[88] & t[89]) | (~t[84] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[85] & t[86] & ~t[88] & ~t[89]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[89]) | (~t[84] & t[85] & t[86] & t[87] & ~t[88]) | (~t[85] & t[86] & t[87] & ~t[89]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[71] = (t[83] & t[84] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[84] & ~t[85] & t[88] & ~t[89]) | (~t[84] & t[85] & ~t[86] & t[87] & t[88]) | (t[85] & ~t[87] & t[88] & ~t[89]);
  assign t[72] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[73] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[76] = t[97] ^ x[11];
  assign t[77] = t[98] ^ x[6];
  assign t[78] = t[99] ^ x[7];
  assign t[79] = t[100] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[101] ^ x[12];
  assign t[81] = t[102] ^ x[9];
  assign t[82] = t[103] ^ x[10];
  assign t[83] = t[104] ^ x[18];
  assign t[84] = t[105] ^ x[27];
  assign t[85] = t[106] ^ x[19];
  assign t[86] = t[107] ^ x[28];
  assign t[87] = t[108] ^ x[29];
  assign t[88] = t[109] ^ x[30];
  assign t[89] = t[110] ^ x[17];
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = t[111] ^ x[25];
  assign t[91] = t[112] ^ x[31];
  assign t[92] = t[113] ^ x[26];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[33];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[24];
  assign t[97] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[98] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[99] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[26]) | (~t[0] & t[26]);
endmodule

module R2ind137(x, y);
 input [38:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[101] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[102] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[42] & t[14]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[114] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[115] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[116] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[117] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[118] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[119] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[11] = ~(t[43] & t[15]);
  assign t[12] = ~(t[44] & t[16]);
  assign t[13] = ~(t[45] & t[17]);
  assign t[14] = ~(t[46]);
  assign t[15] = ~(t[46] & t[18]);
  assign t[16] = ~(t[47]);
  assign t[17] = ~(t[47] & t[19]);
  assign t[18] = ~(t[42]);
  assign t[19] = ~(t[44]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = ~t[23];
  assign t[22] = t[24] ? x[34] : x[33];
  assign t[23] = ~(t[25] ^ t[26]);
  assign t[24] = ~(t[27]);
  assign t[25] = ~t[28];
  assign t[26] = x[2] ? x[35] : t[29];
  assign t[27] = ~(t[4]);
  assign t[28] = x[2] ? x[36] : t[30];
  assign t[29] = ~(t[31] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[33] & t[34]);
  assign t[31] = ~(t[14] & t[35]);
  assign t[32] = ~(t[36] & t[48]);
  assign t[33] = ~(t[16] & t[37]);
  assign t[34] = ~(t[38] & t[49]);
  assign t[35] = ~(t[43]);
  assign t[36] = ~(t[39] & t[18]);
  assign t[37] = ~(t[45]);
  assign t[38] = ~(t[40] & t[19]);
  assign t[39] = ~(t[43] & t[46]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[45] & t[47]);
  assign t[41] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[42] = (t[52] & ~t[54] & ~t[56]) | (~t[53] & t[54] & ~t[55]) | (~t[52] & ~t[54] & t[56]) | (t[53] & t[54] & t[55]);
  assign t[43] = (t[52] & ~t[55]) | (~t[52] & t[55]);
  assign t[44] = (t[57] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[57] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[45] = (t[57] & ~t[60]) | (~t[57] & t[60]);
  assign t[46] = (t[52] & ~t[54] & ~t[55]) | (~t[53] & t[54] & ~t[56]) | (~t[52] & ~t[54] & t[55]) | (t[53] & t[54] & t[56]);
  assign t[47] = (t[57] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[57] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[48] = (t[52] & ~t[62]) | (~t[52] & t[62]);
  assign t[49] = (t[57] & ~t[63]) | (~t[57] & t[63]);
  assign t[4] = ~x[2] & t[41];
  assign t[50] = t[64] ^ x[9];
  assign t[51] = t[65] ^ x[10];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[19];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[28];
  assign t[58] = t[72] ^ x[29];
  assign t[59] = t[73] ^ x[30];
  assign t[5] = ~t[7];
  assign t[60] = t[74] ^ x[31];
  assign t[61] = t[75] ^ x[32];
  assign t[62] = t[76] ^ x[37];
  assign t[63] = t[77] ^ x[38];
  assign t[64] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[65] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = x[2] ? x[11] : t[8];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[72] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[73] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[74] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[76] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[9];
  assign t[79] = t[100] ^ x[4];
  assign t[7] = x[2] ? x[12] : t[9];
  assign t[80] = t[101] ^ x[5];
  assign t[81] = t[102] ^ x[6];
  assign t[82] = t[103] ^ x[10];
  assign t[83] = t[104] ^ x[7];
  assign t[84] = t[105] ^ x[8];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[37];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = ~(t[10] & t[11]);
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[28];
  assign t[93] = t[114] ^ x[29];
  assign t[94] = t[115] ^ x[38];
  assign t[95] = t[116] ^ x[30];
  assign t[96] = t[117] ^ x[31];
  assign t[97] = t[118] ^ x[32];
  assign t[98] = t[119] ^ x[27];
  assign t[99] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0] & ~t[20]) | (~t[0] & t[20]);
endmodule

module R2ind138(x, y);
 input [38:0] x;
 output y;

 wire [117:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[105] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[106] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[107] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[108] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[109] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[10] = ~(t[40] & t[14]);
  assign t[110] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[111] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[112] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[113] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[114] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[115] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[116] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[11] = ~(t[41] & t[15]);
  assign t[12] = ~(t[42] & t[16]);
  assign t[13] = ~(t[43] & t[17]);
  assign t[14] = ~(t[44]);
  assign t[15] = ~(t[44] & t[18]);
  assign t[16] = ~(t[45]);
  assign t[17] = ~(t[45] & t[19]);
  assign t[18] = ~(t[40]);
  assign t[19] = ~(t[42]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = ~t[23];
  assign t[22] = t[24] ? x[34] : x[33];
  assign t[23] = ~(t[25] ^ t[26]);
  assign t[24] = ~(t[27]);
  assign t[25] = ~t[28];
  assign t[26] = x[2] ? x[35] : t[29];
  assign t[27] = ~(t[4]);
  assign t[28] = x[2] ? x[36] : t[30];
  assign t[29] = ~(t[31] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[33] & t[34]);
  assign t[31] = ~(t[14] & t[35]);
  assign t[32] = t[36] | t[46];
  assign t[33] = ~(t[16] & t[37]);
  assign t[34] = t[38] | t[47];
  assign t[35] = ~(t[41]);
  assign t[36] = ~(t[18] | t[14]);
  assign t[37] = ~(t[43]);
  assign t[38] = ~(t[19] | t[16]);
  assign t[39] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50] & ~t[52] & ~t[54]) | (~t[51] & t[52] & ~t[53]) | (~t[50] & ~t[52] & t[54]) | (t[51] & t[52] & t[53]);
  assign t[41] = (t[50] & ~t[53]) | (~t[50] & t[53]);
  assign t[42] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = (t[50] & ~t[52] & ~t[53]) | (~t[51] & t[52] & ~t[54]) | (~t[50] & ~t[52] & t[53]) | (t[51] & t[52] & t[54]);
  assign t[45] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[46] = (t[50] & ~t[60]) | (~t[50] & t[60]);
  assign t[47] = (t[55] & ~t[61]) | (~t[55] & t[61]);
  assign t[48] = t[62] ^ x[9];
  assign t[49] = t[63] ^ x[10];
  assign t[4] = ~x[2] & t[39];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[20];
  assign t[53] = t[67] ^ x[21];
  assign t[54] = t[68] ^ x[22];
  assign t[55] = t[69] ^ x[28];
  assign t[56] = t[70] ^ x[29];
  assign t[57] = t[71] ^ x[30];
  assign t[58] = t[72] ^ x[31];
  assign t[59] = t[73] ^ x[32];
  assign t[5] = ~t[7];
  assign t[60] = t[74] ^ x[37];
  assign t[61] = t[75] ^ x[38];
  assign t[62] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[63] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[65] = (t[84] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & t[84] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[84] & ~t[85] & ~t[88] & ~t[89]) | (t[83] & ~t[84] & t[85] & t[86] & ~t[89]) | (t[83] & ~t[84] & t[87] & t[88] & ~t[89]) | (t[84] & ~t[86] & ~t[88] & t[89]) | (~t[84] & t[86] & t[88] & t[89]);
  assign t[66] = (t[83] & t[84] & t[85] & ~t[86] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[86] & ~t[87] & t[88] & t[89]) | (~t[84] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[85] & t[86] & ~t[88] & ~t[89]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[89]) | (~t[84] & t[85] & t[86] & t[87] & ~t[88]) | (~t[85] & t[86] & t[87] & ~t[89]);
  assign t[67] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[68] = (t[83] & t[84] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[84] & ~t[85] & t[88] & ~t[89]) | (~t[84] & t[85] & ~t[86] & t[87] & t[88]) | (t[85] & ~t[87] & t[88] & ~t[89]);
  assign t[69] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[6] = x[2] ? x[11] : t[8];
  assign t[70] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[71] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[72] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[73] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[74] = (t[83] & t[84] & ~t[85] & t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[85] & ~t[86] & t[87] & ~t[88] & t[89]) | (~t[84] & t[85] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[84] & t[85] & ~t[88] & ~t[89]) | (~t[83] & t[85] & t[86] & ~t[87] & t[88]) | (t[85] & ~t[86] & t[88] & ~t[89]);
  assign t[75] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[76] = t[97] ^ x[9];
  assign t[77] = t[98] ^ x[4];
  assign t[78] = t[99] ^ x[5];
  assign t[79] = t[100] ^ x[6];
  assign t[7] = x[2] ? x[12] : t[9];
  assign t[80] = t[101] ^ x[10];
  assign t[81] = t[102] ^ x[7];
  assign t[82] = t[103] ^ x[8];
  assign t[83] = t[104] ^ x[18];
  assign t[84] = t[105] ^ x[19];
  assign t[85] = t[106] ^ x[37];
  assign t[86] = t[107] ^ x[20];
  assign t[87] = t[108] ^ x[21];
  assign t[88] = t[109] ^ x[22];
  assign t[89] = t[110] ^ x[17];
  assign t[8] = ~(t[10] & t[11]);
  assign t[90] = t[111] ^ x[28];
  assign t[91] = t[112] ^ x[29];
  assign t[92] = t[113] ^ x[38];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[31];
  assign t[95] = t[116] ^ x[32];
  assign t[96] = t[117] ^ x[27];
  assign t[97] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[98] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[99] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0] & ~t[20]) | (~t[0] & t[20]);
endmodule

module R2ind139(x, y);
 input [38:0] x;
 output y;

 wire [117:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[105] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[106] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[107] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[108] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[109] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[10] = ~x[2] & t[39];
  assign t[110] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[111] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[112] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[113] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[114] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[115] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[116] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[117] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[40]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[41]);
  assign t[16] = ~(t[42]);
  assign t[17] = ~(t[43]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[44]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[45]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[43] & t[42]);
  assign t[23] = ~(t[46]);
  assign t[24] = ~(t[45] & t[44]);
  assign t[25] = ~(t[47]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[4] ? x[36] : x[35];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[37] : t[33];
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[12] & t[35]);
  assign t[34] = ~(t[14] & t[36]);
  assign t[35] = t[37] | t[40];
  assign t[36] = t[38] | t[41];
  assign t[37] = ~(t[23] | t[16]);
  assign t[38] = ~(t[25] | t[19]);
  assign t[39] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[41] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[42] = (t[50] & ~t[55] & ~t[56]) | (~t[54] & t[55] & ~t[57]) | (~t[50] & ~t[55] & t[56]) | (t[54] & t[55] & t[57]);
  assign t[43] = (t[50] & ~t[56]) | (~t[50] & t[56]);
  assign t[44] = (t[52] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[52] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[45] = (t[52] & ~t[60]) | (~t[52] & t[60]);
  assign t[46] = (t[50] & ~t[55] & ~t[57]) | (~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[55] & t[57]) | (t[54] & t[55] & t[56]);
  assign t[47] = (t[52] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[52] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[48] = t[62] ^ x[11];
  assign t[49] = t[63] ^ x[12];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[25];
  assign t[53] = t[67] ^ x[26];
  assign t[54] = t[68] ^ x[27];
  assign t[55] = t[69] ^ x[28];
  assign t[56] = t[70] ^ x[29];
  assign t[57] = t[71] ^ x[30];
  assign t[58] = t[72] ^ x[31];
  assign t[59] = t[73] ^ x[32];
  assign t[5] = ~t[8];
  assign t[60] = t[74] ^ x[33];
  assign t[61] = t[75] ^ x[34];
  assign t[62] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[63] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[65] = (t[83] & t[84] & ~t[85] & t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[85] & ~t[86] & t[87] & ~t[88] & t[89]) | (~t[84] & t[85] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[84] & t[85] & ~t[88] & ~t[89]) | (~t[83] & t[85] & t[86] & ~t[87] & t[88]) | (t[85] & ~t[86] & t[88] & ~t[89]);
  assign t[66] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[67] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[68] = (t[84] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & t[84] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[84] & ~t[85] & ~t[88] & ~t[89]) | (t[83] & ~t[84] & t[85] & t[86] & ~t[89]) | (t[83] & ~t[84] & t[87] & t[88] & ~t[89]) | (t[84] & ~t[86] & ~t[88] & t[89]) | (~t[84] & t[86] & t[88] & t[89]);
  assign t[69] = (t[83] & t[84] & t[85] & ~t[86] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[86] & ~t[87] & t[88] & t[89]) | (~t[84] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[85] & t[86] & ~t[88] & ~t[89]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[89]) | (~t[84] & t[85] & t[86] & t[87] & ~t[88]) | (~t[85] & t[86] & t[87] & ~t[89]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[71] = (t[83] & t[84] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[84] & ~t[85] & t[88] & ~t[89]) | (~t[84] & t[85] & ~t[86] & t[87] & t[88]) | (t[85] & ~t[87] & t[88] & ~t[89]);
  assign t[72] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[73] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[76] = t[97] ^ x[11];
  assign t[77] = t[98] ^ x[6];
  assign t[78] = t[99] ^ x[7];
  assign t[79] = t[100] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[101] ^ x[12];
  assign t[81] = t[102] ^ x[9];
  assign t[82] = t[103] ^ x[10];
  assign t[83] = t[104] ^ x[18];
  assign t[84] = t[105] ^ x[27];
  assign t[85] = t[106] ^ x[19];
  assign t[86] = t[107] ^ x[28];
  assign t[87] = t[108] ^ x[29];
  assign t[88] = t[109] ^ x[30];
  assign t[89] = t[110] ^ x[17];
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = t[111] ^ x[25];
  assign t[91] = t[112] ^ x[31];
  assign t[92] = t[113] ^ x[26];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[33];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[24];
  assign t[97] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[98] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[99] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0] & ~t[26]) | (~t[0] & t[26]);
endmodule

module R2ind140(x, y);
 input [42:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[121] ^ x[7];
  assign t[101] = t[122] ^ x[8];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[27];
  assign t[104] = t[125] ^ x[19];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[29];
  assign t[107] = t[128] ^ x[30];
  assign t[108] = t[129] ^ x[17];
  assign t[109] = t[130] ^ x[25];
  assign t[10] = ~(t[14] | t[15]);
  assign t[110] = t[131] ^ x[31];
  assign t[111] = t[132] ^ x[26];
  assign t[112] = t[133] ^ x[32];
  assign t[113] = t[134] ^ x[33];
  assign t[114] = t[135] ^ x[34];
  assign t[115] = t[136] ^ x[24];
  assign t[116] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[117] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[118] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[119] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[11] = ~(t[59] | t[16]);
  assign t[120] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[121] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[124] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[125] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[126] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[127] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[128] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[129] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[131] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[132] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[133] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[134] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[135] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[136] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = ~(t[60] | t[19]);
  assign t[14] = ~(t[61]);
  assign t[15] = ~(t[62]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[63]);
  assign t[18] = ~(t[64]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[65]);
  assign t[21] = ~(t[61] | t[62]);
  assign t[22] = ~(t[66]);
  assign t[23] = ~(t[63] | t[64]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~t[27];
  assign t[26] = t[28] ? x[36] : x[35];
  assign t[27] = ~(t[29] ^ t[30]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~t[32];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = x[2] ? x[37] : t[33];
  assign t[31] = ~(t[4]);
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[61] & t[15]);
  assign t[36] = ~(t[65] & t[39]);
  assign t[37] = ~(t[63] & t[18]);
  assign t[38] = ~(t[66] & t[40]);
  assign t[39] = ~(t[62] & t[14]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[64] & t[17]);
  assign t[41] = ~(t[42] ^ t[43]);
  assign t[42] = ~t[44];
  assign t[43] = t[28] ? x[40] : x[39];
  assign t[44] = ~(t[45] ^ t[46]);
  assign t[45] = ~t[47];
  assign t[46] = x[2] ? x[41] : t[48];
  assign t[47] = x[2] ? x[42] : t[49];
  assign t[48] = ~(t[50] & t[51]);
  assign t[49] = ~(t[52] & t[53]);
  assign t[4] = ~x[2] & t[58];
  assign t[50] = ~(t[15] & t[20]);
  assign t[51] = ~(t[54] & t[59]);
  assign t[52] = ~(t[18] & t[22]);
  assign t[53] = ~(t[55] & t[60]);
  assign t[54] = ~(t[56] & t[14]);
  assign t[55] = ~(t[57] & t[17]);
  assign t[56] = ~(t[65] & t[62]);
  assign t[57] = ~(t[66] & t[64]);
  assign t[58] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[59] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[5] = ~t[7];
  assign t[60] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[61] = (t[69] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[69] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[62] = (t[69] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[69] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[63] = (t[71] & ~t[78] & ~t[80]) | (~t[77] & t[78] & ~t[79]) | (~t[71] & ~t[78] & t[80]) | (t[77] & t[78] & t[79]);
  assign t[64] = (t[71] & ~t[78] & ~t[79]) | (~t[77] & t[78] & ~t[80]) | (~t[71] & ~t[78] & t[79]) | (t[77] & t[78] & t[80]);
  assign t[65] = (t[69] & ~t[75]) | (~t[69] & t[75]);
  assign t[66] = (t[71] & ~t[79]) | (~t[71] & t[79]);
  assign t[67] = t[81] ^ x[9];
  assign t[68] = t[82] ^ x[10];
  assign t[69] = t[83] ^ x[18];
  assign t[6] = x[2] ? x[11] : t[8];
  assign t[70] = t[84] ^ x[19];
  assign t[71] = t[85] ^ x[25];
  assign t[72] = t[86] ^ x[26];
  assign t[73] = t[87] ^ x[27];
  assign t[74] = t[88] ^ x[28];
  assign t[75] = t[89] ^ x[29];
  assign t[76] = t[90] ^ x[30];
  assign t[77] = t[91] ^ x[31];
  assign t[78] = t[92] ^ x[32];
  assign t[79] = t[93] ^ x[33];
  assign t[7] = x[2] ? x[12] : t[9];
  assign t[80] = t[94] ^ x[34];
  assign t[81] = (t[95] & ~t[97] & ~t[98] & ~t[99] & ~t[100]) | (t[95] & ~t[96] & ~t[98] & ~t[99] & ~t[101]) | (t[95] & ~t[96] & ~t[97] & ~t[100] & ~t[101]) | (~t[95] & t[96] & t[97] & t[98] & ~t[101]) | (~t[95] & t[96] & t[99] & t[100] & ~t[101]) | (t[95] & ~t[97] & ~t[99] & t[101]) | (~t[95] & t[97] & t[99] & t[101]);
  assign t[82] = (t[95] & t[96] & ~t[97] & ~t[99] & t[100] & ~t[101]) | (t[95] & t[97] & ~t[98] & ~t[99] & ~t[100] & t[101]) | (~t[96] & ~t[97] & t[99] & ~t[100] & ~t[101]) | (~t[95] & ~t[97] & ~t[98] & t[99] & ~t[100]) | (~t[95] & ~t[96] & ~t[98] & t[99] & ~t[101]) | (~t[95] & ~t[97] & t[98] & t[99] & t[100]) | (t[98] & t[99] & ~t[100] & ~t[101]);
  assign t[83] = (t[102] & ~t[104] & ~t[105] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & ~t[105] & ~t[106] & ~t[108]) | (t[102] & ~t[103] & ~t[104] & ~t[107] & ~t[108]) | (~t[102] & t[103] & t[104] & t[105] & ~t[108]) | (~t[102] & t[103] & t[106] & t[107] & ~t[108]) | (t[102] & ~t[104] & ~t[106] & t[108]) | (~t[102] & t[104] & t[106] & t[108]);
  assign t[84] = (t[102] & t[103] & ~t[104] & t[105] & ~t[106] & ~t[108]) | (t[102] & ~t[104] & ~t[105] & t[106] & ~t[107] & t[108]) | (~t[103] & t[104] & ~t[105] & ~t[106] & ~t[108]) | (~t[102] & t[104] & ~t[105] & ~t[106] & ~t[107]) | (~t[102] & ~t[103] & t[104] & ~t[107] & ~t[108]) | (~t[102] & t[104] & t[105] & ~t[106] & t[107]) | (t[104] & ~t[105] & t[107] & ~t[108]);
  assign t[85] = (t[109] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[110] & ~t[111] & ~t[114] & ~t[115]) | (~t[109] & t[110] & t[111] & t[112] & ~t[115]) | (~t[109] & t[110] & t[113] & t[114] & ~t[115]) | (t[109] & ~t[111] & ~t[113] & t[115]) | (~t[109] & t[111] & t[113] & t[115]);
  assign t[86] = (t[109] & t[110] & ~t[111] & t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[111] & ~t[112] & t[113] & ~t[114] & t[115]) | (~t[110] & t[111] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[110] & t[111] & ~t[114] & ~t[115]) | (~t[109] & t[111] & t[112] & ~t[113] & t[114]) | (t[111] & ~t[112] & t[114] & ~t[115]);
  assign t[87] = (t[103] & ~t[104] & ~t[105] & ~t[106] & ~t[107]) | (~t[102] & t[103] & ~t[105] & ~t[106] & ~t[108]) | (~t[102] & t[103] & ~t[104] & ~t[107] & ~t[108]) | (t[102] & ~t[103] & t[104] & t[105] & ~t[108]) | (t[102] & ~t[103] & t[106] & t[107] & ~t[108]) | (t[103] & ~t[105] & ~t[107] & t[108]) | (~t[103] & t[105] & t[107] & t[108]);
  assign t[88] = (t[102] & t[103] & t[104] & ~t[105] & ~t[107] & ~t[108]) | (t[103] & ~t[104] & ~t[105] & ~t[106] & t[107] & t[108]) | (~t[103] & ~t[104] & t[105] & ~t[106] & ~t[107]) | (~t[102] & ~t[104] & t[105] & ~t[107] & ~t[108]) | (~t[102] & ~t[103] & t[105] & ~t[106] & ~t[108]) | (~t[103] & t[104] & t[105] & t[106] & ~t[107]) | (~t[104] & t[105] & t[106] & ~t[108]);
  assign t[89] = (t[102] & t[103] & ~t[104] & ~t[106] & t[107] & ~t[108]) | (t[102] & t[104] & ~t[105] & ~t[106] & ~t[107] & t[108]) | (~t[103] & ~t[104] & t[106] & ~t[107] & ~t[108]) | (~t[102] & ~t[104] & ~t[105] & t[106] & ~t[107]) | (~t[102] & ~t[103] & ~t[105] & t[106] & ~t[108]) | (~t[102] & ~t[104] & t[105] & t[106] & t[107]) | (t[105] & t[106] & ~t[107] & ~t[108]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[90] = (t[102] & t[103] & ~t[105] & t[106] & ~t[107] & ~t[108]) | (t[103] & ~t[104] & t[105] & ~t[106] & ~t[107] & t[108]) | (~t[103] & ~t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[105] & ~t[106] & t[107] & ~t[108]) | (~t[102] & ~t[103] & ~t[104] & t[107] & ~t[108]) | (~t[103] & t[104] & ~t[105] & t[106] & t[107]) | (t[104] & ~t[106] & t[107] & ~t[108]);
  assign t[91] = (t[110] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & t[110] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[110] & ~t[111] & ~t[114] & ~t[115]) | (t[109] & ~t[110] & t[111] & t[112] & ~t[115]) | (t[109] & ~t[110] & t[113] & t[114] & ~t[115]) | (t[110] & ~t[112] & ~t[114] & t[115]) | (~t[110] & t[112] & t[114] & t[115]);
  assign t[92] = (t[109] & t[110] & t[111] & ~t[112] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[112] & ~t[113] & t[114] & t[115]) | (~t[110] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[111] & t[112] & ~t[114] & ~t[115]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[115]) | (~t[110] & t[111] & t[112] & t[113] & ~t[114]) | (~t[111] & t[112] & t[113] & ~t[115]);
  assign t[93] = (t[109] & t[110] & ~t[111] & ~t[113] & t[114] & ~t[115]) | (t[109] & t[111] & ~t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & t[113] & ~t[114] & ~t[115]) | (~t[109] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[109] & ~t[110] & ~t[112] & t[113] & ~t[115]) | (~t[109] & ~t[111] & t[112] & t[113] & t[114]) | (t[112] & t[113] & ~t[114] & ~t[115]);
  assign t[94] = (t[109] & t[110] & ~t[112] & t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[109] & ~t[110] & ~t[111] & t[114] & ~t[115]) | (~t[110] & t[111] & ~t[112] & t[113] & t[114]) | (t[111] & ~t[113] & t[114] & ~t[115]);
  assign t[95] = t[116] ^ x[9];
  assign t[96] = t[117] ^ x[4];
  assign t[97] = t[118] ^ x[5];
  assign t[98] = t[119] ^ x[6];
  assign t[99] = t[120] ^ x[10];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[24] & ~t[41]) | (~t[0] & t[24] & ~t[41]) | (~t[0] & ~t[24] & t[41]) | (t[0] & t[24] & t[41]);
endmodule

module R2ind141(x, y);
 input [42:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[121] ^ x[19];
  assign t[101] = t[122] ^ x[28];
  assign t[102] = t[123] ^ x[29];
  assign t[103] = t[124] ^ x[30];
  assign t[104] = t[125] ^ x[17];
  assign t[105] = t[126] ^ x[25];
  assign t[106] = t[127] ^ x[31];
  assign t[107] = t[128] ^ x[26];
  assign t[108] = t[129] ^ x[32];
  assign t[109] = t[130] ^ x[33];
  assign t[10] = ~(t[14] | t[15]);
  assign t[110] = t[131] ^ x[34];
  assign t[111] = t[132] ^ x[24];
  assign t[112] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[113] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[114] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[115] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[11] = ~(t[55] | t[16]);
  assign t[120] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[121] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[122] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[123] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[124] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[125] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[126] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[127] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[128] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[129] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[131] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[132] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = ~(t[56] | t[19]);
  assign t[14] = ~(t[57]);
  assign t[15] = ~(t[58]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[59]);
  assign t[18] = ~(t[60]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[61]);
  assign t[21] = ~(t[57] | t[58]);
  assign t[22] = ~(t[62]);
  assign t[23] = ~(t[59] | t[60]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~t[27];
  assign t[26] = t[28] ? x[36] : x[35];
  assign t[27] = ~(t[29] ^ t[30]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~t[32];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = x[2] ? x[37] : t[33];
  assign t[31] = ~(t[4]);
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[57] & t[15]);
  assign t[36] = ~(t[61] & t[39]);
  assign t[37] = ~(t[59] & t[18]);
  assign t[38] = ~(t[62] & t[40]);
  assign t[39] = ~(t[58] & t[14]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[60] & t[17]);
  assign t[41] = ~(t[42] ^ t[43]);
  assign t[42] = ~t[44];
  assign t[43] = t[4] ? x[40] : x[39];
  assign t[44] = ~(t[45] ^ t[46]);
  assign t[45] = ~t[47];
  assign t[46] = x[2] ? x[41] : t[48];
  assign t[47] = x[2] ? x[42] : t[49];
  assign t[48] = ~(t[50] & t[51]);
  assign t[49] = ~(t[52] & t[53]);
  assign t[4] = ~x[2] & t[54];
  assign t[50] = ~(t[15] & t[20]);
  assign t[51] = t[10] | t[55];
  assign t[52] = ~(t[18] & t[22]);
  assign t[53] = t[12] | t[56];
  assign t[54] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[55] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[56] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[57] = (t[65] & ~t[70] & ~t[72]) | (~t[69] & t[70] & ~t[71]) | (~t[65] & ~t[70] & t[72]) | (t[69] & t[70] & t[71]);
  assign t[58] = (t[65] & ~t[70] & ~t[71]) | (~t[69] & t[70] & ~t[72]) | (~t[65] & ~t[70] & t[71]) | (t[69] & t[70] & t[72]);
  assign t[59] = (t[67] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[67] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[5] = ~t[7];
  assign t[60] = (t[67] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[67] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[61] = (t[65] & ~t[71]) | (~t[65] & t[71]);
  assign t[62] = (t[67] & ~t[75]) | (~t[67] & t[75]);
  assign t[63] = t[77] ^ x[9];
  assign t[64] = t[78] ^ x[10];
  assign t[65] = t[79] ^ x[18];
  assign t[66] = t[80] ^ x[19];
  assign t[67] = t[81] ^ x[25];
  assign t[68] = t[82] ^ x[26];
  assign t[69] = t[83] ^ x[27];
  assign t[6] = x[2] ? x[11] : t[8];
  assign t[70] = t[84] ^ x[28];
  assign t[71] = t[85] ^ x[29];
  assign t[72] = t[86] ^ x[30];
  assign t[73] = t[87] ^ x[31];
  assign t[74] = t[88] ^ x[32];
  assign t[75] = t[89] ^ x[33];
  assign t[76] = t[90] ^ x[34];
  assign t[77] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[78] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[79] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[7] = x[2] ? x[12] : t[9];
  assign t[80] = (t[98] & t[99] & ~t[100] & t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[100] & ~t[101] & t[102] & ~t[103] & t[104]) | (~t[99] & t[100] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[99] & t[100] & ~t[103] & ~t[104]) | (~t[98] & t[100] & t[101] & ~t[102] & t[103]) | (t[100] & ~t[101] & t[103] & ~t[104]);
  assign t[81] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[82] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[83] = (t[99] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & t[99] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[99] & ~t[100] & ~t[103] & ~t[104]) | (t[98] & ~t[99] & t[100] & t[101] & ~t[104]) | (t[98] & ~t[99] & t[102] & t[103] & ~t[104]) | (t[99] & ~t[101] & ~t[103] & t[104]) | (~t[99] & t[101] & t[103] & t[104]);
  assign t[84] = (t[98] & t[99] & t[100] & ~t[101] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[101] & ~t[102] & t[103] & t[104]) | (~t[99] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[100] & t[101] & ~t[103] & ~t[104]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[104]) | (~t[99] & t[100] & t[101] & t[102] & ~t[103]) | (~t[100] & t[101] & t[102] & ~t[104]);
  assign t[85] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[86] = (t[98] & t[99] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[98] & ~t[99] & ~t[100] & t[103] & ~t[104]) | (~t[99] & t[100] & ~t[101] & t[102] & t[103]) | (t[100] & ~t[102] & t[103] & ~t[104]);
  assign t[87] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[88] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[89] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[90] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[91] = t[112] ^ x[9];
  assign t[92] = t[113] ^ x[4];
  assign t[93] = t[114] ^ x[5];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[10];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[8];
  assign t[98] = t[119] ^ x[18];
  assign t[99] = t[120] ^ x[27];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[24] & ~t[41]) | (~t[0] & t[24] & ~t[41]) | (~t[0] & ~t[24] & t[41]) | (t[0] & t[24] & t[41]);
endmodule

module R2ind142(x, y);
 input [38:0] x;
 output y;

 wire [121:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[121] ^ x[24];
  assign t[101] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[102] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[103] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[104] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[107] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[108] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[109] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[110] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[111] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[112] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[113] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[114] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[115] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[116] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[117] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[118] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[119] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[11] = ~(t[44] | t[16]);
  assign t[120] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[121] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[45] | t[19]);
  assign t[14] = ~(t[46]);
  assign t[15] = ~(t[47]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[48]);
  assign t[18] = ~(t[49]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[50]);
  assign t[21] = ~(t[46] | t[47]);
  assign t[22] = ~(t[51]);
  assign t[23] = ~(t[48] | t[49]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~t[27];
  assign t[26] = t[28] ? x[36] : x[35];
  assign t[27] = ~(t[29] ^ t[30]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~t[32];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = x[2] ? x[37] : t[33];
  assign t[31] = ~(t[4]);
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[15] & t[20]);
  assign t[36] = ~(t[39] & t[44]);
  assign t[37] = ~(t[18] & t[22]);
  assign t[38] = ~(t[40] & t[45]);
  assign t[39] = ~(t[41] & t[14]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[42] & t[17]);
  assign t[41] = ~(t[50] & t[47]);
  assign t[42] = ~(t[51] & t[49]);
  assign t[43] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[44] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[54] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[54] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[47] = (t[54] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[54] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[48] = (t[56] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[56] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[49] = (t[56] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[56] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[4] = ~x[2] & t[43];
  assign t[50] = (t[54] & ~t[60]) | (~t[54] & t[60]);
  assign t[51] = (t[56] & ~t[64]) | (~t[56] & t[64]);
  assign t[52] = t[66] ^ x[9];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[18];
  assign t[55] = t[69] ^ x[19];
  assign t[56] = t[70] ^ x[25];
  assign t[57] = t[71] ^ x[26];
  assign t[58] = t[72] ^ x[27];
  assign t[59] = t[73] ^ x[28];
  assign t[5] = ~t[7];
  assign t[60] = t[74] ^ x[29];
  assign t[61] = t[75] ^ x[30];
  assign t[62] = t[76] ^ x[31];
  assign t[63] = t[77] ^ x[32];
  assign t[64] = t[78] ^ x[33];
  assign t[65] = t[79] ^ x[34];
  assign t[66] = (t[80] & ~t[82] & ~t[83] & ~t[84] & ~t[85]) | (t[80] & ~t[81] & ~t[83] & ~t[84] & ~t[86]) | (t[80] & ~t[81] & ~t[82] & ~t[85] & ~t[86]) | (~t[80] & t[81] & t[82] & t[83] & ~t[86]) | (~t[80] & t[81] & t[84] & t[85] & ~t[86]) | (t[80] & ~t[82] & ~t[84] & t[86]) | (~t[80] & t[82] & t[84] & t[86]);
  assign t[67] = (t[80] & t[81] & ~t[82] & ~t[84] & t[85] & ~t[86]) | (t[80] & t[82] & ~t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[82] & t[84] & ~t[85] & ~t[86]) | (~t[80] & ~t[82] & ~t[83] & t[84] & ~t[85]) | (~t[80] & ~t[81] & ~t[83] & t[84] & ~t[86]) | (~t[80] & ~t[82] & t[83] & t[84] & t[85]) | (t[83] & t[84] & ~t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[89] & ~t[90] & ~t[91] & ~t[92]) | (t[87] & ~t[88] & ~t[90] & ~t[91] & ~t[93]) | (t[87] & ~t[88] & ~t[89] & ~t[92] & ~t[93]) | (~t[87] & t[88] & t[89] & t[90] & ~t[93]) | (~t[87] & t[88] & t[91] & t[92] & ~t[93]) | (t[87] & ~t[89] & ~t[91] & t[93]) | (~t[87] & t[89] & t[91] & t[93]);
  assign t[69] = (t[87] & t[88] & ~t[89] & t[90] & ~t[91] & ~t[93]) | (t[87] & ~t[89] & ~t[90] & t[91] & ~t[92] & t[93]) | (~t[88] & t[89] & ~t[90] & ~t[91] & ~t[93]) | (~t[87] & t[89] & ~t[90] & ~t[91] & ~t[92]) | (~t[87] & ~t[88] & t[89] & ~t[92] & ~t[93]) | (~t[87] & t[89] & t[90] & ~t[91] & t[92]) | (t[89] & ~t[90] & t[92] & ~t[93]);
  assign t[6] = x[2] ? x[11] : t[8];
  assign t[70] = (t[94] & ~t[96] & ~t[97] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & ~t[97] & ~t[98] & ~t[100]) | (t[94] & ~t[95] & ~t[96] & ~t[99] & ~t[100]) | (~t[94] & t[95] & t[96] & t[97] & ~t[100]) | (~t[94] & t[95] & t[98] & t[99] & ~t[100]) | (t[94] & ~t[96] & ~t[98] & t[100]) | (~t[94] & t[96] & t[98] & t[100]);
  assign t[71] = (t[94] & t[95] & ~t[96] & t[97] & ~t[98] & ~t[100]) | (t[94] & ~t[96] & ~t[97] & t[98] & ~t[99] & t[100]) | (~t[95] & t[96] & ~t[97] & ~t[98] & ~t[100]) | (~t[94] & t[96] & ~t[97] & ~t[98] & ~t[99]) | (~t[94] & ~t[95] & t[96] & ~t[99] & ~t[100]) | (~t[94] & t[96] & t[97] & ~t[98] & t[99]) | (t[96] & ~t[97] & t[99] & ~t[100]);
  assign t[72] = (t[88] & ~t[89] & ~t[90] & ~t[91] & ~t[92]) | (~t[87] & t[88] & ~t[90] & ~t[91] & ~t[93]) | (~t[87] & t[88] & ~t[89] & ~t[92] & ~t[93]) | (t[87] & ~t[88] & t[89] & t[90] & ~t[93]) | (t[87] & ~t[88] & t[91] & t[92] & ~t[93]) | (t[88] & ~t[90] & ~t[92] & t[93]) | (~t[88] & t[90] & t[92] & t[93]);
  assign t[73] = (t[87] & t[88] & t[89] & ~t[90] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & ~t[90] & ~t[91] & t[92] & t[93]) | (~t[88] & ~t[89] & t[90] & ~t[91] & ~t[92]) | (~t[87] & ~t[89] & t[90] & ~t[92] & ~t[93]) | (~t[87] & ~t[88] & t[90] & ~t[91] & ~t[93]) | (~t[88] & t[89] & t[90] & t[91] & ~t[92]) | (~t[89] & t[90] & t[91] & ~t[93]);
  assign t[74] = (t[87] & t[88] & ~t[89] & ~t[91] & t[92] & ~t[93]) | (t[87] & t[89] & ~t[90] & ~t[91] & ~t[92] & t[93]) | (~t[88] & ~t[89] & t[91] & ~t[92] & ~t[93]) | (~t[87] & ~t[89] & ~t[90] & t[91] & ~t[92]) | (~t[87] & ~t[88] & ~t[90] & t[91] & ~t[93]) | (~t[87] & ~t[89] & t[90] & t[91] & t[92]) | (t[90] & t[91] & ~t[92] & ~t[93]);
  assign t[75] = (t[87] & t[88] & ~t[90] & t[91] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & t[90] & ~t[91] & ~t[92] & t[93]) | (~t[88] & ~t[89] & ~t[90] & ~t[91] & t[92]) | (~t[87] & ~t[90] & ~t[91] & t[92] & ~t[93]) | (~t[87] & ~t[88] & ~t[89] & t[92] & ~t[93]) | (~t[88] & t[89] & ~t[90] & t[91] & t[92]) | (t[89] & ~t[91] & t[92] & ~t[93]);
  assign t[76] = (t[95] & ~t[96] & ~t[97] & ~t[98] & ~t[99]) | (~t[94] & t[95] & ~t[97] & ~t[98] & ~t[100]) | (~t[94] & t[95] & ~t[96] & ~t[99] & ~t[100]) | (t[94] & ~t[95] & t[96] & t[97] & ~t[100]) | (t[94] & ~t[95] & t[98] & t[99] & ~t[100]) | (t[95] & ~t[97] & ~t[99] & t[100]) | (~t[95] & t[97] & t[99] & t[100]);
  assign t[77] = (t[94] & t[95] & t[96] & ~t[97] & ~t[99] & ~t[100]) | (t[95] & ~t[96] & ~t[97] & ~t[98] & t[99] & t[100]) | (~t[95] & ~t[96] & t[97] & ~t[98] & ~t[99]) | (~t[94] & ~t[96] & t[97] & ~t[99] & ~t[100]) | (~t[94] & ~t[95] & t[97] & ~t[98] & ~t[100]) | (~t[95] & t[96] & t[97] & t[98] & ~t[99]) | (~t[96] & t[97] & t[98] & ~t[100]);
  assign t[78] = (t[94] & t[95] & ~t[96] & ~t[98] & t[99] & ~t[100]) | (t[94] & t[96] & ~t[97] & ~t[98] & ~t[99] & t[100]) | (~t[95] & ~t[96] & t[98] & ~t[99] & ~t[100]) | (~t[94] & ~t[96] & ~t[97] & t[98] & ~t[99]) | (~t[94] & ~t[95] & ~t[97] & t[98] & ~t[100]) | (~t[94] & ~t[96] & t[97] & t[98] & t[99]) | (t[97] & t[98] & ~t[99] & ~t[100]);
  assign t[79] = (t[94] & t[95] & ~t[97] & t[98] & ~t[99] & ~t[100]) | (t[95] & ~t[96] & t[97] & ~t[98] & ~t[99] & t[100]) | (~t[95] & ~t[96] & ~t[97] & ~t[98] & t[99]) | (~t[94] & ~t[97] & ~t[98] & t[99] & ~t[100]) | (~t[94] & ~t[95] & ~t[96] & t[99] & ~t[100]) | (~t[95] & t[96] & ~t[97] & t[98] & t[99]) | (t[96] & ~t[98] & t[99] & ~t[100]);
  assign t[7] = x[2] ? x[12] : t[9];
  assign t[80] = t[101] ^ x[9];
  assign t[81] = t[102] ^ x[4];
  assign t[82] = t[103] ^ x[5];
  assign t[83] = t[104] ^ x[6];
  assign t[84] = t[105] ^ x[10];
  assign t[85] = t[106] ^ x[7];
  assign t[86] = t[107] ^ x[8];
  assign t[87] = t[108] ^ x[18];
  assign t[88] = t[109] ^ x[27];
  assign t[89] = t[110] ^ x[19];
  assign t[8] = ~(t[10] | t[11]);
  assign t[90] = t[111] ^ x[28];
  assign t[91] = t[112] ^ x[29];
  assign t[92] = t[113] ^ x[30];
  assign t[93] = t[114] ^ x[17];
  assign t[94] = t[115] ^ x[25];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[26];
  assign t[97] = t[118] ^ x[32];
  assign t[98] = t[119] ^ x[33];
  assign t[99] = t[120] ^ x[34];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[24]) | (~t[0] & t[24]);
endmodule

module R2ind143(x, y);
 input [38:0] x;
 output y;

 wire [115:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[103] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[104] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[105] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[106] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[107] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[108] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[109] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[110] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[111] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[112] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[113] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[114] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[115] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[11] = ~(t[38] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[39] | t[19]);
  assign t[14] = ~(t[40]);
  assign t[15] = ~(t[41]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[42]);
  assign t[18] = ~(t[43]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[44]);
  assign t[21] = ~(t[40] | t[41]);
  assign t[22] = ~(t[45]);
  assign t[23] = ~(t[42] | t[43]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~t[27];
  assign t[26] = t[4] ? x[36] : x[35];
  assign t[27] = ~(t[28] ^ t[29]);
  assign t[28] = ~t[30];
  assign t[29] = x[2] ? x[37] : t[31];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = x[2] ? x[38] : t[32];
  assign t[31] = ~(t[33] & t[34]);
  assign t[32] = ~(t[35] & t[36]);
  assign t[33] = ~(t[15] & t[20]);
  assign t[34] = t[10] | t[38];
  assign t[35] = ~(t[18] & t[22]);
  assign t[36] = t[12] | t[39];
  assign t[37] = (t[46] & ~t[47]) | (~t[46] & t[47]);
  assign t[38] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[39] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[48] & ~t[53] & ~t[55]) | (~t[52] & t[53] & ~t[54]) | (~t[48] & ~t[53] & t[55]) | (t[52] & t[53] & t[54]);
  assign t[41] = (t[48] & ~t[53] & ~t[54]) | (~t[52] & t[53] & ~t[55]) | (~t[48] & ~t[53] & t[54]) | (t[52] & t[53] & t[55]);
  assign t[42] = (t[50] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[50] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[43] = (t[50] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[50] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[44] = (t[48] & ~t[54]) | (~t[48] & t[54]);
  assign t[45] = (t[50] & ~t[58]) | (~t[50] & t[58]);
  assign t[46] = t[60] ^ x[9];
  assign t[47] = t[61] ^ x[10];
  assign t[48] = t[62] ^ x[18];
  assign t[49] = t[63] ^ x[19];
  assign t[4] = ~x[2] & t[37];
  assign t[50] = t[64] ^ x[25];
  assign t[51] = t[65] ^ x[26];
  assign t[52] = t[66] ^ x[27];
  assign t[53] = t[67] ^ x[28];
  assign t[54] = t[68] ^ x[29];
  assign t[55] = t[69] ^ x[30];
  assign t[56] = t[70] ^ x[31];
  assign t[57] = t[71] ^ x[32];
  assign t[58] = t[72] ^ x[33];
  assign t[59] = t[73] ^ x[34];
  assign t[5] = ~t[7];
  assign t[60] = (t[74] & ~t[76] & ~t[77] & ~t[78] & ~t[79]) | (t[74] & ~t[75] & ~t[77] & ~t[78] & ~t[80]) | (t[74] & ~t[75] & ~t[76] & ~t[79] & ~t[80]) | (~t[74] & t[75] & t[76] & t[77] & ~t[80]) | (~t[74] & t[75] & t[78] & t[79] & ~t[80]) | (t[74] & ~t[76] & ~t[78] & t[80]) | (~t[74] & t[76] & t[78] & t[80]);
  assign t[61] = (t[74] & t[75] & ~t[76] & ~t[78] & t[79] & ~t[80]) | (t[74] & t[76] & ~t[77] & ~t[78] & ~t[79] & t[80]) | (~t[75] & ~t[76] & t[78] & ~t[79] & ~t[80]) | (~t[74] & ~t[76] & ~t[77] & t[78] & ~t[79]) | (~t[74] & ~t[75] & ~t[77] & t[78] & ~t[80]) | (~t[74] & ~t[76] & t[77] & t[78] & t[79]) | (t[77] & t[78] & ~t[79] & ~t[80]);
  assign t[62] = (t[81] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (t[81] & ~t[82] & ~t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[82] & ~t[83] & ~t[86] & ~t[87]) | (~t[81] & t[82] & t[83] & t[84] & ~t[87]) | (~t[81] & t[82] & t[85] & t[86] & ~t[87]) | (t[81] & ~t[83] & ~t[85] & t[87]) | (~t[81] & t[83] & t[85] & t[87]);
  assign t[63] = (t[81] & t[82] & ~t[83] & t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[83] & ~t[84] & t[85] & ~t[86] & t[87]) | (~t[82] & t[83] & ~t[84] & ~t[85] & ~t[87]) | (~t[81] & t[83] & ~t[84] & ~t[85] & ~t[86]) | (~t[81] & ~t[82] & t[83] & ~t[86] & ~t[87]) | (~t[81] & t[83] & t[84] & ~t[85] & t[86]) | (t[83] & ~t[84] & t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[90] & ~t[91] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & ~t[91] & ~t[92] & ~t[94]) | (t[88] & ~t[89] & ~t[90] & ~t[93] & ~t[94]) | (~t[88] & t[89] & t[90] & t[91] & ~t[94]) | (~t[88] & t[89] & t[92] & t[93] & ~t[94]) | (t[88] & ~t[90] & ~t[92] & t[94]) | (~t[88] & t[90] & t[92] & t[94]);
  assign t[65] = (t[88] & t[89] & ~t[90] & t[91] & ~t[92] & ~t[94]) | (t[88] & ~t[90] & ~t[91] & t[92] & ~t[93] & t[94]) | (~t[89] & t[90] & ~t[91] & ~t[92] & ~t[94]) | (~t[88] & t[90] & ~t[91] & ~t[92] & ~t[93]) | (~t[88] & ~t[89] & t[90] & ~t[93] & ~t[94]) | (~t[88] & t[90] & t[91] & ~t[92] & t[93]) | (t[90] & ~t[91] & t[93] & ~t[94]);
  assign t[66] = (t[82] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (~t[81] & t[82] & ~t[84] & ~t[85] & ~t[87]) | (~t[81] & t[82] & ~t[83] & ~t[86] & ~t[87]) | (t[81] & ~t[82] & t[83] & t[84] & ~t[87]) | (t[81] & ~t[82] & t[85] & t[86] & ~t[87]) | (t[82] & ~t[84] & ~t[86] & t[87]) | (~t[82] & t[84] & t[86] & t[87]);
  assign t[67] = (t[81] & t[82] & t[83] & ~t[84] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & ~t[84] & ~t[85] & t[86] & t[87]) | (~t[82] & ~t[83] & t[84] & ~t[85] & ~t[86]) | (~t[81] & ~t[83] & t[84] & ~t[86] & ~t[87]) | (~t[81] & ~t[82] & t[84] & ~t[85] & ~t[87]) | (~t[82] & t[83] & t[84] & t[85] & ~t[86]) | (~t[83] & t[84] & t[85] & ~t[87]);
  assign t[68] = (t[81] & t[82] & ~t[83] & ~t[85] & t[86] & ~t[87]) | (t[81] & t[83] & ~t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & t[85] & ~t[86] & ~t[87]) | (~t[81] & ~t[83] & ~t[84] & t[85] & ~t[86]) | (~t[81] & ~t[82] & ~t[84] & t[85] & ~t[87]) | (~t[81] & ~t[83] & t[84] & t[85] & t[86]) | (t[84] & t[85] & ~t[86] & ~t[87]);
  assign t[69] = (t[81] & t[82] & ~t[84] & t[85] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[84] & ~t[85] & t[86] & ~t[87]) | (~t[81] & ~t[82] & ~t[83] & t[86] & ~t[87]) | (~t[82] & t[83] & ~t[84] & t[85] & t[86]) | (t[83] & ~t[85] & t[86] & ~t[87]);
  assign t[6] = x[2] ? x[11] : t[8];
  assign t[70] = (t[89] & ~t[90] & ~t[91] & ~t[92] & ~t[93]) | (~t[88] & t[89] & ~t[91] & ~t[92] & ~t[94]) | (~t[88] & t[89] & ~t[90] & ~t[93] & ~t[94]) | (t[88] & ~t[89] & t[90] & t[91] & ~t[94]) | (t[88] & ~t[89] & t[92] & t[93] & ~t[94]) | (t[89] & ~t[91] & ~t[93] & t[94]) | (~t[89] & t[91] & t[93] & t[94]);
  assign t[71] = (t[88] & t[89] & t[90] & ~t[91] & ~t[93] & ~t[94]) | (t[89] & ~t[90] & ~t[91] & ~t[92] & t[93] & t[94]) | (~t[89] & ~t[90] & t[91] & ~t[92] & ~t[93]) | (~t[88] & ~t[90] & t[91] & ~t[93] & ~t[94]) | (~t[88] & ~t[89] & t[91] & ~t[92] & ~t[94]) | (~t[89] & t[90] & t[91] & t[92] & ~t[93]) | (~t[90] & t[91] & t[92] & ~t[94]);
  assign t[72] = (t[88] & t[89] & ~t[90] & ~t[92] & t[93] & ~t[94]) | (t[88] & t[90] & ~t[91] & ~t[92] & ~t[93] & t[94]) | (~t[89] & ~t[90] & t[92] & ~t[93] & ~t[94]) | (~t[88] & ~t[90] & ~t[91] & t[92] & ~t[93]) | (~t[88] & ~t[89] & ~t[91] & t[92] & ~t[94]) | (~t[88] & ~t[90] & t[91] & t[92] & t[93]) | (t[91] & t[92] & ~t[93] & ~t[94]);
  assign t[73] = (t[88] & t[89] & ~t[91] & t[92] & ~t[93] & ~t[94]) | (t[89] & ~t[90] & t[91] & ~t[92] & ~t[93] & t[94]) | (~t[89] & ~t[90] & ~t[91] & ~t[92] & t[93]) | (~t[88] & ~t[91] & ~t[92] & t[93] & ~t[94]) | (~t[88] & ~t[89] & ~t[90] & t[93] & ~t[94]) | (~t[89] & t[90] & ~t[91] & t[92] & t[93]) | (t[90] & ~t[92] & t[93] & ~t[94]);
  assign t[74] = t[95] ^ x[9];
  assign t[75] = t[96] ^ x[4];
  assign t[76] = t[97] ^ x[5];
  assign t[77] = t[98] ^ x[6];
  assign t[78] = t[99] ^ x[10];
  assign t[79] = t[100] ^ x[7];
  assign t[7] = x[2] ? x[12] : t[9];
  assign t[80] = t[101] ^ x[8];
  assign t[81] = t[102] ^ x[18];
  assign t[82] = t[103] ^ x[27];
  assign t[83] = t[104] ^ x[19];
  assign t[84] = t[105] ^ x[28];
  assign t[85] = t[106] ^ x[29];
  assign t[86] = t[107] ^ x[30];
  assign t[87] = t[108] ^ x[17];
  assign t[88] = t[109] ^ x[25];
  assign t[89] = t[110] ^ x[31];
  assign t[8] = ~(t[10] | t[11]);
  assign t[90] = t[111] ^ x[26];
  assign t[91] = t[112] ^ x[32];
  assign t[92] = t[113] ^ x[33];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[24];
  assign t[95] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[96] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[97] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[98] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[99] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[24]) | (~t[0] & t[24]);
endmodule

module R2ind144(x, y);
 input [38:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[101] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[102] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~x[2] & t[41];
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[114] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[115] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[116] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[117] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[118] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[119] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[42] & t[16]);
  assign t[13] = ~(t[43] & t[17]);
  assign t[14] = ~(t[44] & t[18]);
  assign t[15] = ~(t[45] & t[19]);
  assign t[16] = ~(t[46]);
  assign t[17] = ~(t[46] & t[20]);
  assign t[18] = ~(t[47]);
  assign t[19] = ~(t[47] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[42]);
  assign t[21] = ~(t[44]);
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = ~t[25];
  assign t[24] = t[4] ? x[34] : x[33];
  assign t[25] = ~(t[26] ^ t[27]);
  assign t[26] = ~t[28];
  assign t[27] = x[2] ? x[35] : t[29];
  assign t[28] = x[2] ? x[36] : t[30];
  assign t[29] = ~(t[31] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[33] & t[34]);
  assign t[31] = ~(t[16] & t[35]);
  assign t[32] = ~(t[36] & t[48]);
  assign t[33] = ~(t[18] & t[37]);
  assign t[34] = ~(t[38] & t[49]);
  assign t[35] = ~(t[43]);
  assign t[36] = ~(t[39] & t[20]);
  assign t[37] = ~(t[45]);
  assign t[38] = ~(t[40] & t[21]);
  assign t[39] = ~(t[43] & t[46]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[45] & t[47]);
  assign t[41] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[42] = (t[52] & ~t[54] & ~t[56]) | (~t[53] & t[54] & ~t[55]) | (~t[52] & ~t[54] & t[56]) | (t[53] & t[54] & t[55]);
  assign t[43] = (t[52] & ~t[55]) | (~t[52] & t[55]);
  assign t[44] = (t[57] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[57] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[45] = (t[57] & ~t[60]) | (~t[57] & t[60]);
  assign t[46] = (t[52] & ~t[54] & ~t[55]) | (~t[53] & t[54] & ~t[56]) | (~t[52] & ~t[54] & t[55]) | (t[53] & t[54] & t[56]);
  assign t[47] = (t[57] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[57] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[48] = (t[52] & ~t[62]) | (~t[52] & t[62]);
  assign t[49] = (t[57] & ~t[63]) | (~t[57] & t[63]);
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[11];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[19];
  assign t[54] = t[68] ^ x[20];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[28];
  assign t[58] = t[72] ^ x[29];
  assign t[59] = t[73] ^ x[30];
  assign t[5] = ~t[8];
  assign t[60] = t[74] ^ x[31];
  assign t[61] = t[75] ^ x[32];
  assign t[62] = t[76] ^ x[37];
  assign t[63] = t[77] ^ x[38];
  assign t[64] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[65] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[72] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[73] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[74] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[76] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[11];
  assign t[79] = t[100] ^ x[6];
  assign t[7] = ~(t[10]);
  assign t[80] = t[101] ^ x[7];
  assign t[81] = t[102] ^ x[8];
  assign t[82] = t[103] ^ x[12];
  assign t[83] = t[104] ^ x[9];
  assign t[84] = t[105] ^ x[10];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[37];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[28];
  assign t[93] = t[114] ^ x[29];
  assign t[94] = t[115] ^ x[38];
  assign t[95] = t[116] ^ x[30];
  assign t[96] = t[117] ^ x[31];
  assign t[97] = t[118] ^ x[32];
  assign t[98] = t[119] ^ x[27];
  assign t[99] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0] & ~t[22]) | (~t[0] & t[22]);
endmodule

module R2ind145(x, y);
 input [38:0] x;
 output y;

 wire [117:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[105] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[106] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[107] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[108] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[109] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[10] = ~x[2] & t[39];
  assign t[110] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[111] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[112] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[113] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[114] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[115] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[116] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[40] & t[16]);
  assign t[13] = ~(t[41] & t[17]);
  assign t[14] = ~(t[42] & t[18]);
  assign t[15] = ~(t[43] & t[19]);
  assign t[16] = ~(t[44]);
  assign t[17] = ~(t[44] & t[20]);
  assign t[18] = ~(t[45]);
  assign t[19] = ~(t[45] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40]);
  assign t[21] = ~(t[42]);
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = ~t[25];
  assign t[24] = t[10] ? x[34] : x[33];
  assign t[25] = ~(t[26] ^ t[27]);
  assign t[26] = ~t[28];
  assign t[27] = x[2] ? x[35] : t[29];
  assign t[28] = x[2] ? x[36] : t[30];
  assign t[29] = ~(t[31] & t[32]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[33] & t[34]);
  assign t[31] = ~(t[16] & t[35]);
  assign t[32] = t[36] | t[46];
  assign t[33] = ~(t[18] & t[37]);
  assign t[34] = t[38] | t[47];
  assign t[35] = ~(t[41]);
  assign t[36] = ~(t[20] | t[16]);
  assign t[37] = ~(t[43]);
  assign t[38] = ~(t[21] | t[18]);
  assign t[39] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50] & ~t[52] & ~t[54]) | (~t[51] & t[52] & ~t[53]) | (~t[50] & ~t[52] & t[54]) | (t[51] & t[52] & t[53]);
  assign t[41] = (t[50] & ~t[53]) | (~t[50] & t[53]);
  assign t[42] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = (t[50] & ~t[52] & ~t[53]) | (~t[51] & t[52] & ~t[54]) | (~t[50] & ~t[52] & t[53]) | (t[51] & t[52] & t[54]);
  assign t[45] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[46] = (t[50] & ~t[60]) | (~t[50] & t[60]);
  assign t[47] = (t[55] & ~t[61]) | (~t[55] & t[61]);
  assign t[48] = t[62] ^ x[11];
  assign t[49] = t[63] ^ x[12];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[20];
  assign t[53] = t[67] ^ x[21];
  assign t[54] = t[68] ^ x[22];
  assign t[55] = t[69] ^ x[28];
  assign t[56] = t[70] ^ x[29];
  assign t[57] = t[71] ^ x[30];
  assign t[58] = t[72] ^ x[31];
  assign t[59] = t[73] ^ x[32];
  assign t[5] = ~t[8];
  assign t[60] = t[74] ^ x[37];
  assign t[61] = t[75] ^ x[38];
  assign t[62] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[63] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[65] = (t[84] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & t[84] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[84] & ~t[85] & ~t[88] & ~t[89]) | (t[83] & ~t[84] & t[85] & t[86] & ~t[89]) | (t[83] & ~t[84] & t[87] & t[88] & ~t[89]) | (t[84] & ~t[86] & ~t[88] & t[89]) | (~t[84] & t[86] & t[88] & t[89]);
  assign t[66] = (t[83] & t[84] & t[85] & ~t[86] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[86] & ~t[87] & t[88] & t[89]) | (~t[84] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[85] & t[86] & ~t[88] & ~t[89]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[89]) | (~t[84] & t[85] & t[86] & t[87] & ~t[88]) | (~t[85] & t[86] & t[87] & ~t[89]);
  assign t[67] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[68] = (t[83] & t[84] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[84] & ~t[85] & t[88] & ~t[89]) | (~t[84] & t[85] & ~t[86] & t[87] & t[88]) | (t[85] & ~t[87] & t[88] & ~t[89]);
  assign t[69] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[71] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[72] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[73] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[74] = (t[83] & t[84] & ~t[85] & t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[85] & ~t[86] & t[87] & ~t[88] & t[89]) | (~t[84] & t[85] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[84] & t[85] & ~t[88] & ~t[89]) | (~t[83] & t[85] & t[86] & ~t[87] & t[88]) | (t[85] & ~t[86] & t[88] & ~t[89]);
  assign t[75] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[76] = t[97] ^ x[11];
  assign t[77] = t[98] ^ x[6];
  assign t[78] = t[99] ^ x[7];
  assign t[79] = t[100] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[101] ^ x[12];
  assign t[81] = t[102] ^ x[9];
  assign t[82] = t[103] ^ x[10];
  assign t[83] = t[104] ^ x[18];
  assign t[84] = t[105] ^ x[19];
  assign t[85] = t[106] ^ x[37];
  assign t[86] = t[107] ^ x[20];
  assign t[87] = t[108] ^ x[21];
  assign t[88] = t[109] ^ x[22];
  assign t[89] = t[110] ^ x[17];
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = t[111] ^ x[28];
  assign t[91] = t[112] ^ x[29];
  assign t[92] = t[113] ^ x[38];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[31];
  assign t[95] = t[116] ^ x[32];
  assign t[96] = t[117] ^ x[27];
  assign t[97] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[98] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[99] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0] & ~t[22]) | (~t[0] & t[22]);
endmodule

module R2ind146(x, y);
 input [38:0] x;
 output y;

 wire [117:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[105] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[106] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[107] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[108] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[109] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[10] = ~x[2] & t[39];
  assign t[110] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[111] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[112] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[113] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[114] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[115] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[116] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[117] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[40]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[41]);
  assign t[16] = ~(t[42]);
  assign t[17] = ~(t[43]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[44]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[45]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[43] & t[42]);
  assign t[23] = ~(t[46]);
  assign t[24] = ~(t[45] & t[44]);
  assign t[25] = ~(t[47]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[10] ? x[36] : x[35];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[37] : t[33];
  assign t[32] = x[2] ? x[38] : t[34];
  assign t[33] = ~(t[12] & t[35]);
  assign t[34] = ~(t[14] & t[36]);
  assign t[35] = t[37] | t[40];
  assign t[36] = t[38] | t[41];
  assign t[37] = ~(t[23] | t[16]);
  assign t[38] = ~(t[25] | t[19]);
  assign t[39] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[41] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[42] = (t[50] & ~t[55] & ~t[56]) | (~t[54] & t[55] & ~t[57]) | (~t[50] & ~t[55] & t[56]) | (t[54] & t[55] & t[57]);
  assign t[43] = (t[50] & ~t[56]) | (~t[50] & t[56]);
  assign t[44] = (t[52] & ~t[59] & ~t[60]) | (~t[58] & t[59] & ~t[61]) | (~t[52] & ~t[59] & t[60]) | (t[58] & t[59] & t[61]);
  assign t[45] = (t[52] & ~t[60]) | (~t[52] & t[60]);
  assign t[46] = (t[50] & ~t[55] & ~t[57]) | (~t[54] & t[55] & ~t[56]) | (~t[50] & ~t[55] & t[57]) | (t[54] & t[55] & t[56]);
  assign t[47] = (t[52] & ~t[59] & ~t[61]) | (~t[58] & t[59] & ~t[60]) | (~t[52] & ~t[59] & t[61]) | (t[58] & t[59] & t[60]);
  assign t[48] = t[62] ^ x[11];
  assign t[49] = t[63] ^ x[12];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[25];
  assign t[53] = t[67] ^ x[26];
  assign t[54] = t[68] ^ x[27];
  assign t[55] = t[69] ^ x[28];
  assign t[56] = t[70] ^ x[29];
  assign t[57] = t[71] ^ x[30];
  assign t[58] = t[72] ^ x[31];
  assign t[59] = t[73] ^ x[32];
  assign t[5] = ~t[8];
  assign t[60] = t[74] ^ x[33];
  assign t[61] = t[75] ^ x[34];
  assign t[62] = (t[76] & ~t[78] & ~t[79] & ~t[80] & ~t[81]) | (t[76] & ~t[77] & ~t[79] & ~t[80] & ~t[82]) | (t[76] & ~t[77] & ~t[78] & ~t[81] & ~t[82]) | (~t[76] & t[77] & t[78] & t[79] & ~t[82]) | (~t[76] & t[77] & t[80] & t[81] & ~t[82]) | (t[76] & ~t[78] & ~t[80] & t[82]) | (~t[76] & t[78] & t[80] & t[82]);
  assign t[63] = (t[76] & t[77] & ~t[78] & ~t[80] & t[81] & ~t[82]) | (t[76] & t[78] & ~t[79] & ~t[80] & ~t[81] & t[82]) | (~t[77] & ~t[78] & t[80] & ~t[81] & ~t[82]) | (~t[76] & ~t[78] & ~t[79] & t[80] & ~t[81]) | (~t[76] & ~t[77] & ~t[79] & t[80] & ~t[82]) | (~t[76] & ~t[78] & t[79] & t[80] & t[81]) | (t[79] & t[80] & ~t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[65] = (t[83] & t[84] & ~t[85] & t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[85] & ~t[86] & t[87] & ~t[88] & t[89]) | (~t[84] & t[85] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[84] & t[85] & ~t[88] & ~t[89]) | (~t[83] & t[85] & t[86] & ~t[87] & t[88]) | (t[85] & ~t[86] & t[88] & ~t[89]);
  assign t[66] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[67] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[68] = (t[84] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & t[84] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[84] & ~t[85] & ~t[88] & ~t[89]) | (t[83] & ~t[84] & t[85] & t[86] & ~t[89]) | (t[83] & ~t[84] & t[87] & t[88] & ~t[89]) | (t[84] & ~t[86] & ~t[88] & t[89]) | (~t[84] & t[86] & t[88] & t[89]);
  assign t[69] = (t[83] & t[84] & t[85] & ~t[86] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[86] & ~t[87] & t[88] & t[89]) | (~t[84] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[85] & t[86] & ~t[88] & ~t[89]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[89]) | (~t[84] & t[85] & t[86] & t[87] & ~t[88]) | (~t[85] & t[86] & t[87] & ~t[89]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[71] = (t[83] & t[84] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[84] & ~t[85] & t[88] & ~t[89]) | (~t[84] & t[85] & ~t[86] & t[87] & t[88]) | (t[85] & ~t[87] & t[88] & ~t[89]);
  assign t[72] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[73] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[76] = t[97] ^ x[11];
  assign t[77] = t[98] ^ x[6];
  assign t[78] = t[99] ^ x[7];
  assign t[79] = t[100] ^ x[8];
  assign t[7] = ~(t[10]);
  assign t[80] = t[101] ^ x[12];
  assign t[81] = t[102] ^ x[9];
  assign t[82] = t[103] ^ x[10];
  assign t[83] = t[104] ^ x[18];
  assign t[84] = t[105] ^ x[27];
  assign t[85] = t[106] ^ x[19];
  assign t[86] = t[107] ^ x[28];
  assign t[87] = t[108] ^ x[29];
  assign t[88] = t[109] ^ x[30];
  assign t[89] = t[110] ^ x[17];
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = t[111] ^ x[25];
  assign t[91] = t[112] ^ x[31];
  assign t[92] = t[113] ^ x[26];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[33];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[24];
  assign t[97] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[98] = (x[5] & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0);
  assign t[99] = (x[5] & ~1'b0) | (~x[5] & 1'b0);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0] & ~t[26]) | (~t[0] & t[26]);
endmodule

module R2ind147(x, y);
 input [66:0] x;
 output y;

 wire [199:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[130] & ~t[132] & ~t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[133] & ~t[134] & ~t[136]) | (t[130] & ~t[131] & ~t[132] & ~t[135] & ~t[136]) | (~t[130] & t[131] & t[132] & t[133] & ~t[136]) | (~t[130] & t[131] & t[134] & t[135] & ~t[136]) | (t[130] & ~t[132] & ~t[134] & t[136]) | (~t[130] & t[132] & t[134] & t[136]);
  assign t[101] = (t[130] & t[131] & ~t[132] & ~t[134] & t[135] & ~t[136]) | (t[130] & t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[136]) | (~t[130] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[130] & ~t[131] & ~t[133] & t[134] & ~t[136]) | (~t[130] & ~t[132] & t[133] & t[134] & t[135]) | (t[133] & t[134] & ~t[135] & ~t[136]);
  assign t[102] = (t[137] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & ~t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[138] & ~t[139] & ~t[142] & ~t[143]) | (~t[137] & t[138] & t[139] & t[140] & ~t[143]) | (~t[137] & t[138] & t[141] & t[142] & ~t[143]) | (t[137] & ~t[139] & ~t[141] & t[143]) | (~t[137] & t[139] & t[141] & t[143]);
  assign t[103] = (t[137] & t[138] & ~t[139] & t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[139] & ~t[140] & t[141] & ~t[142] & t[143]) | (~t[138] & t[139] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[138] & t[139] & ~t[142] & ~t[143]) | (~t[137] & t[139] & t[140] & ~t[141] & t[142]) | (t[139] & ~t[140] & t[142] & ~t[143]);
  assign t[104] = (t[124] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & t[124] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[124] & ~t[125] & ~t[128] & ~t[129]) | (t[123] & ~t[124] & t[125] & t[126] & ~t[129]) | (t[123] & ~t[124] & t[127] & t[128] & ~t[129]) | (t[124] & ~t[126] & ~t[128] & t[129]) | (~t[124] & t[126] & t[128] & t[129]);
  assign t[105] = (t[123] & t[124] & t[125] & ~t[126] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[126] & ~t[127] & t[128] & t[129]) | (~t[124] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[125] & t[126] & ~t[128] & ~t[129]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[129]) | (~t[124] & t[125] & t[126] & t[127] & ~t[128]) | (~t[125] & t[126] & t[127] & ~t[129]);
  assign t[106] = (t[123] & t[124] & ~t[125] & ~t[127] & t[128] & ~t[129]) | (t[123] & t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[129]) | (~t[123] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[123] & ~t[124] & ~t[126] & t[127] & ~t[129]) | (~t[123] & ~t[125] & t[126] & t[127] & t[128]) | (t[126] & t[127] & ~t[128] & ~t[129]);
  assign t[107] = (t[123] & t[124] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[123] & ~t[124] & ~t[125] & t[128] & ~t[129]) | (~t[124] & t[125] & ~t[126] & t[127] & t[128]) | (t[125] & ~t[127] & t[128] & ~t[129]);
  assign t[108] = (t[138] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & t[138] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[138] & ~t[139] & ~t[142] & ~t[143]) | (t[137] & ~t[138] & t[139] & t[140] & ~t[143]) | (t[137] & ~t[138] & t[141] & t[142] & ~t[143]) | (t[138] & ~t[140] & ~t[142] & t[143]) | (~t[138] & t[140] & t[142] & t[143]);
  assign t[109] = (t[137] & t[138] & t[139] & ~t[140] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[140] & ~t[141] & t[142] & t[143]) | (~t[138] & ~t[139] & t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[139] & t[140] & ~t[142] & ~t[143]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[143]) | (~t[138] & t[139] & t[140] & t[141] & ~t[142]) | (~t[139] & t[140] & t[141] & ~t[143]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (t[137] & t[138] & ~t[139] & ~t[141] & t[142] & ~t[143]) | (t[137] & t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[143]) | (~t[137] & ~t[139] & ~t[140] & t[141] & ~t[142]) | (~t[137] & ~t[138] & ~t[140] & t[141] & ~t[143]) | (~t[137] & ~t[139] & t[140] & t[141] & t[142]) | (t[140] & t[141] & ~t[142] & ~t[143]);
  assign t[111] = (t[137] & t[138] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[137] & ~t[138] & ~t[139] & t[142] & ~t[143]) | (~t[138] & t[139] & ~t[140] & t[141] & t[142]) | (t[139] & ~t[141] & t[142] & ~t[143]);
  assign t[112] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[113] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[114] = (t[151] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & ~t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[152] & ~t[153] & ~t[156] & ~t[157]) | (~t[151] & t[152] & t[153] & t[154] & ~t[157]) | (~t[151] & t[152] & t[155] & t[156] & ~t[157]) | (t[151] & ~t[153] & ~t[155] & t[157]) | (~t[151] & t[153] & t[155] & t[157]);
  assign t[115] = (t[151] & t[152] & ~t[153] & ~t[155] & t[156] & ~t[157]) | (t[151] & t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[157]) | (~t[151] & ~t[153] & ~t[154] & t[155] & ~t[156]) | (~t[151] & ~t[152] & ~t[154] & t[155] & ~t[157]) | (~t[151] & ~t[153] & t[154] & t[155] & t[156]) | (t[154] & t[155] & ~t[156] & ~t[157]);
  assign t[116] = t[158] ^ x[9];
  assign t[117] = t[159] ^ x[4];
  assign t[118] = t[160] ^ x[5];
  assign t[119] = t[161] ^ x[6];
  assign t[11] = ~(t[15]);
  assign t[120] = t[162] ^ x[10];
  assign t[121] = t[163] ^ x[7];
  assign t[122] = t[164] ^ x[8];
  assign t[123] = t[165] ^ x[18];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[19];
  assign t[126] = t[168] ^ x[36];
  assign t[127] = t[169] ^ x[37];
  assign t[128] = t[170] ^ x[38];
  assign t[129] = t[171] ^ x[17];
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = t[172] ^ x[26];
  assign t[131] = t[173] ^ x[21];
  assign t[132] = t[174] ^ x[22];
  assign t[133] = t[175] ^ x[23];
  assign t[134] = t[176] ^ x[27];
  assign t[135] = t[177] ^ x[24];
  assign t[136] = t[178] ^ x[25];
  assign t[137] = t[179] ^ x[33];
  assign t[138] = t[180] ^ x[39];
  assign t[139] = t[181] ^ x[34];
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = t[182] ^ x[40];
  assign t[141] = t[183] ^ x[41];
  assign t[142] = t[184] ^ x[42];
  assign t[143] = t[185] ^ x[32];
  assign t[144] = t[186] ^ x[51];
  assign t[145] = t[187] ^ x[46];
  assign t[146] = t[188] ^ x[47];
  assign t[147] = t[189] ^ x[48];
  assign t[148] = t[190] ^ x[52];
  assign t[149] = t[191] ^ x[49];
  assign t[14] = ~(t[65] | t[20]);
  assign t[150] = t[192] ^ x[50];
  assign t[151] = t[193] ^ x[63];
  assign t[152] = t[194] ^ x[58];
  assign t[153] = t[195] ^ x[59];
  assign t[154] = t[196] ^ x[60];
  assign t[155] = t[197] ^ x[64];
  assign t[156] = t[198] ^ x[61];
  assign t[157] = t[199] ^ x[62];
  assign t[158] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[159] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[66];
  assign t[160] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[161] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[164] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[165] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[166] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[167] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[168] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[169] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[16] = ~(t[21] | t[22]);
  assign t[170] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[171] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[172] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[173] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[174] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[175] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[176] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[177] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[178] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[179] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[17] = ~(t[67] | t[23]);
  assign t[180] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[181] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[182] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[183] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[184] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[185] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[186] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[187] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[188] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[189] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[18] = ~(t[68]);
  assign t[190] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[192] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[193] = (x[57] & ~1'b0 & ~1'b0) | (~x[57] & 1'b0 & ~1'b0) | (~x[57] & ~1'b0 & 1'b0) | (x[57] & 1'b0 & 1'b0);
  assign t[194] = (x[57] & ~1'b0 & ~1'b0) | (~x[57] & 1'b0 & ~1'b0) | (~x[57] & ~1'b0 & 1'b0) | (x[57] & 1'b0 & 1'b0);
  assign t[195] = (x[57] & ~1'b0) | (~x[57] & 1'b0);
  assign t[196] = (x[57] & ~1'b0) | (~x[57] & 1'b0);
  assign t[197] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[198] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[199] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = ~(t[69]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[70]);
  assign t[22] = ~(t[71]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[72]);
  assign t[25] = ~(t[68] | t[69]);
  assign t[26] = ~(t[73]);
  assign t[27] = ~(t[70] | t[71]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[74];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[68] & t[19]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[72] & t[43]);
  assign t[41] = ~(t[70] & t[22]);
  assign t[42] = ~(t[73] & t[44]);
  assign t[43] = ~(t[69] & t[18]);
  assign t[44] = ~(t[71] & t[21]);
  assign t[45] = ~(t[46] ^ t[47]);
  assign t[46] = t[48];
  assign t[47] = ~(t[49] ^ t[50]);
  assign t[48] = ~(t[51] ^ t[52]);
  assign t[49] = t[8] ? x[56] : x[55];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = ~x[2] & t[75];
  assign t[51] = ~t[53];
  assign t[52] = x[2] ? x[65] : t[54];
  assign t[53] = x[2] ? x[66] : t[55];
  assign t[54] = ~(t[56] & t[57]);
  assign t[55] = ~(t[58] & t[59]);
  assign t[56] = ~(t[19] & t[24]);
  assign t[57] = ~(t[60] & t[65]);
  assign t[58] = ~(t[22] & t[26]);
  assign t[59] = ~(t[61] & t[67]);
  assign t[5] = ~(~x[2] & ~t[64]);
  assign t[60] = ~(t[62] & t[18]);
  assign t[61] = ~(t[63] & t[21]);
  assign t[62] = ~(t[72] & t[69]);
  assign t[63] = ~(t[73] & t[71]);
  assign t[64] = (t[76] & ~t[77]) | (~t[76] & t[77]);
  assign t[65] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[66] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[67] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[68] = (t[78] & ~t[85] & ~t[87]) | (~t[84] & t[85] & ~t[86]) | (~t[78] & ~t[85] & t[87]) | (t[84] & t[85] & t[86]);
  assign t[69] = (t[78] & ~t[85] & ~t[86]) | (~t[84] & t[85] & ~t[87]) | (~t[78] & ~t[85] & t[86]) | (t[84] & t[85] & t[87]);
  assign t[6] = ~t[9];
  assign t[70] = (t[82] & ~t[89] & ~t[91]) | (~t[88] & t[89] & ~t[90]) | (~t[82] & ~t[89] & t[91]) | (t[88] & t[89] & t[90]);
  assign t[71] = (t[82] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[91]) | (~t[82] & ~t[89] & t[90]) | (t[88] & t[89] & t[91]);
  assign t[72] = (t[78] & ~t[86]) | (~t[78] & t[86]);
  assign t[73] = (t[82] & ~t[90]) | (~t[82] & t[90]);
  assign t[74] = (t[92] & ~t[93]) | (~t[92] & t[93]);
  assign t[75] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[76] = t[96] ^ x[9];
  assign t[77] = t[97] ^ x[10];
  assign t[78] = t[98] ^ x[18];
  assign t[79] = t[99] ^ x[19];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[26];
  assign t[81] = t[101] ^ x[27];
  assign t[82] = t[102] ^ x[33];
  assign t[83] = t[103] ^ x[34];
  assign t[84] = t[104] ^ x[35];
  assign t[85] = t[105] ^ x[36];
  assign t[86] = t[106] ^ x[37];
  assign t[87] = t[107] ^ x[38];
  assign t[88] = t[108] ^ x[39];
  assign t[89] = t[109] ^ x[40];
  assign t[8] = ~(t[11]);
  assign t[90] = t[110] ^ x[41];
  assign t[91] = t[111] ^ x[42];
  assign t[92] = t[112] ^ x[51];
  assign t[93] = t[113] ^ x[52];
  assign t[94] = t[114] ^ x[63];
  assign t[95] = t[115] ^ x[64];
  assign t[96] = (t[116] & ~t[118] & ~t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[119] & ~t[120] & ~t[122]) | (t[116] & ~t[117] & ~t[118] & ~t[121] & ~t[122]) | (~t[116] & t[117] & t[118] & t[119] & ~t[122]) | (~t[116] & t[117] & t[120] & t[121] & ~t[122]) | (t[116] & ~t[118] & ~t[120] & t[122]) | (~t[116] & t[118] & t[120] & t[122]);
  assign t[97] = (t[116] & t[117] & ~t[118] & ~t[120] & t[121] & ~t[122]) | (t[116] & t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[122]) | (~t[116] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[116] & ~t[117] & ~t[119] & t[120] & ~t[122]) | (~t[116] & ~t[118] & t[119] & t[120] & t[121]) | (t[119] & t[120] & ~t[121] & ~t[122]);
  assign t[98] = (t[123] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[124] & ~t[125] & ~t[128] & ~t[129]) | (~t[123] & t[124] & t[125] & t[126] & ~t[129]) | (~t[123] & t[124] & t[127] & t[128] & ~t[129]) | (t[123] & ~t[125] & ~t[127] & t[129]) | (~t[123] & t[125] & t[127] & t[129]);
  assign t[99] = (t[123] & t[124] & ~t[125] & t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[125] & ~t[126] & t[127] & ~t[128] & t[129]) | (~t[124] & t[125] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[124] & t[125] & ~t[128] & ~t[129]) | (~t[123] & t[125] & t[126] & ~t[127] & t[128]) | (t[125] & ~t[126] & t[128] & ~t[129]);
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28] & ~t[45]) | (~t[0] & t[28] & ~t[45]) | (~t[0] & ~t[28] & t[45]) | (t[0] & t[28] & t[45]);
endmodule

module R2ind148(x, y);
 input [58:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[101] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[102] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[103] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[104] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[105] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[106] = t[141] ^ x[9];
  assign t[107] = t[142] ^ x[4];
  assign t[108] = t[143] ^ x[5];
  assign t[109] = t[144] ^ x[6];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[145] ^ x[10];
  assign t[111] = t[146] ^ x[7];
  assign t[112] = t[147] ^ x[8];
  assign t[113] = t[148] ^ x[18];
  assign t[114] = t[149] ^ x[35];
  assign t[115] = t[150] ^ x[19];
  assign t[116] = t[151] ^ x[36];
  assign t[117] = t[152] ^ x[37];
  assign t[118] = t[153] ^ x[38];
  assign t[119] = t[154] ^ x[17];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[26];
  assign t[121] = t[156] ^ x[21];
  assign t[122] = t[157] ^ x[22];
  assign t[123] = t[158] ^ x[23];
  assign t[124] = t[159] ^ x[27];
  assign t[125] = t[160] ^ x[24];
  assign t[126] = t[161] ^ x[25];
  assign t[127] = t[162] ^ x[33];
  assign t[128] = t[163] ^ x[39];
  assign t[129] = t[164] ^ x[34];
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = t[165] ^ x[40];
  assign t[131] = t[166] ^ x[41];
  assign t[132] = t[167] ^ x[42];
  assign t[133] = t[168] ^ x[32];
  assign t[134] = t[169] ^ x[51];
  assign t[135] = t[170] ^ x[46];
  assign t[136] = t[171] ^ x[47];
  assign t[137] = t[172] ^ x[48];
  assign t[138] = t[173] ^ x[52];
  assign t[139] = t[174] ^ x[49];
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = t[175] ^ x[50];
  assign t[141] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[142] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[143] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[144] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[149] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[14] = ~(t[60] | t[20]);
  assign t[150] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[151] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[152] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[153] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[154] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[155] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[156] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[157] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[158] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[61];
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[163] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[164] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[165] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[166] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[167] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[168] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[169] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[16] = ~(t[21] | t[22]);
  assign t[170] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[171] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[172] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[174] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[175] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[17] = ~(t[62] | t[23]);
  assign t[18] = ~(t[63]);
  assign t[19] = ~(t[64]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[65]);
  assign t[22] = ~(t[66]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[67]);
  assign t[25] = ~(t[63] | t[64]);
  assign t[26] = ~(t[68]);
  assign t[27] = ~(t[65] | t[66]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[69];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[63] & t[19]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[67] & t[43]);
  assign t[41] = ~(t[65] & t[22]);
  assign t[42] = ~(t[68] & t[44]);
  assign t[43] = ~(t[64] & t[18]);
  assign t[44] = ~(t[66] & t[21]);
  assign t[45] = ~(t[46] ^ t[47]);
  assign t[46] = t[48];
  assign t[47] = ~t[49];
  assign t[48] = ~(t[50] ^ t[51]);
  assign t[49] = t[8] ? x[56] : x[55];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = ~t[52];
  assign t[51] = x[2] ? x[57] : t[53];
  assign t[52] = x[2] ? x[58] : t[54];
  assign t[53] = ~(t[55] & t[56]);
  assign t[54] = ~(t[57] & t[58]);
  assign t[55] = ~(t[19] & t[24]);
  assign t[56] = t[13] | t[60];
  assign t[57] = ~(t[22] & t[26]);
  assign t[58] = t[16] | t[62];
  assign t[59] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[5] = ~(~x[2] & ~t[59]);
  assign t[60] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[61] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[62] = (t[76] & ~t[77]) | (~t[76] & t[77]);
  assign t[63] = (t[72] & ~t[79] & ~t[81]) | (~t[78] & t[79] & ~t[80]) | (~t[72] & ~t[79] & t[81]) | (t[78] & t[79] & t[80]);
  assign t[64] = (t[72] & ~t[79] & ~t[80]) | (~t[78] & t[79] & ~t[81]) | (~t[72] & ~t[79] & t[80]) | (t[78] & t[79] & t[81]);
  assign t[65] = (t[76] & ~t[83] & ~t[85]) | (~t[82] & t[83] & ~t[84]) | (~t[76] & ~t[83] & t[85]) | (t[82] & t[83] & t[84]);
  assign t[66] = (t[76] & ~t[83] & ~t[84]) | (~t[82] & t[83] & ~t[85]) | (~t[76] & ~t[83] & t[84]) | (t[82] & t[83] & t[85]);
  assign t[67] = (t[72] & ~t[80]) | (~t[72] & t[80]);
  assign t[68] = (t[76] & ~t[84]) | (~t[76] & t[84]);
  assign t[69] = (t[86] & ~t[87]) | (~t[86] & t[87]);
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[9];
  assign t[71] = t[89] ^ x[10];
  assign t[72] = t[90] ^ x[18];
  assign t[73] = t[91] ^ x[19];
  assign t[74] = t[92] ^ x[26];
  assign t[75] = t[93] ^ x[27];
  assign t[76] = t[94] ^ x[33];
  assign t[77] = t[95] ^ x[34];
  assign t[78] = t[96] ^ x[35];
  assign t[79] = t[97] ^ x[36];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[98] ^ x[37];
  assign t[81] = t[99] ^ x[38];
  assign t[82] = t[100] ^ x[39];
  assign t[83] = t[101] ^ x[40];
  assign t[84] = t[102] ^ x[41];
  assign t[85] = t[103] ^ x[42];
  assign t[86] = t[104] ^ x[51];
  assign t[87] = t[105] ^ x[52];
  assign t[88] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[89] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[93] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[94] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[95] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[96] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[97] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[98] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[99] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28] & ~t[45]) | (~t[0] & t[28] & ~t[45]) | (~t[0] & ~t[28] & t[45]) | (t[0] & t[28] & t[45]);
endmodule

module R2ind149(x, y);
 input [54:0] x;
 output y;

 wire [163:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[8];
  assign t[101] = t[136] ^ x[18];
  assign t[102] = t[137] ^ x[35];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[36];
  assign t[105] = t[140] ^ x[37];
  assign t[106] = t[141] ^ x[38];
  assign t[107] = t[142] ^ x[17];
  assign t[108] = t[143] ^ x[26];
  assign t[109] = t[144] ^ x[21];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[145] ^ x[22];
  assign t[111] = t[146] ^ x[23];
  assign t[112] = t[147] ^ x[27];
  assign t[113] = t[148] ^ x[24];
  assign t[114] = t[149] ^ x[25];
  assign t[115] = t[150] ^ x[33];
  assign t[116] = t[151] ^ x[39];
  assign t[117] = t[152] ^ x[34];
  assign t[118] = t[153] ^ x[40];
  assign t[119] = t[154] ^ x[41];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[42];
  assign t[121] = t[156] ^ x[32];
  assign t[122] = t[157] ^ x[51];
  assign t[123] = t[158] ^ x[46];
  assign t[124] = t[159] ^ x[47];
  assign t[125] = t[160] ^ x[48];
  assign t[126] = t[161] ^ x[52];
  assign t[127] = t[162] ^ x[49];
  assign t[128] = t[163] ^ x[50];
  assign t[129] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[131] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[132] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[133] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[134] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[135] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[136] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[137] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[138] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[139] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[141] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[142] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[143] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[144] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[145] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[146] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[149] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = ~(t[48] | t[20]);
  assign t[150] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[151] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[152] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[153] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[154] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[155] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[156] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[157] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[158] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[159] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[15] = ~x[2] & t[49];
  assign t[160] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[50] | t[23]);
  assign t[18] = ~(t[51]);
  assign t[19] = ~(t[52]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[53]);
  assign t[22] = ~(t[54]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[55]);
  assign t[25] = ~(t[51] | t[52]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] | t[54]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[57];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[19] & t[24]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[43] & t[48]);
  assign t[41] = ~(t[22] & t[26]);
  assign t[42] = ~(t[44] & t[50]);
  assign t[43] = ~(t[45] & t[18]);
  assign t[44] = ~(t[46] & t[21]);
  assign t[45] = ~(t[55] & t[52]);
  assign t[46] = ~(t[56] & t[54]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[49] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[60] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[60] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[52] = (t[60] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[60] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[53] = (t[64] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[64] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[54] = (t[64] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[64] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[55] = (t[60] & ~t[68]) | (~t[60] & t[68]);
  assign t[56] = (t[64] & ~t[72]) | (~t[64] & t[72]);
  assign t[57] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[58] = t[76] ^ x[9];
  assign t[59] = t[77] ^ x[10];
  assign t[5] = ~(~x[2] & ~t[47]);
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[26];
  assign t[63] = t[81] ^ x[27];
  assign t[64] = t[82] ^ x[33];
  assign t[65] = t[83] ^ x[34];
  assign t[66] = t[84] ^ x[35];
  assign t[67] = t[85] ^ x[36];
  assign t[68] = t[86] ^ x[37];
  assign t[69] = t[87] ^ x[38];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[39];
  assign t[71] = t[89] ^ x[40];
  assign t[72] = t[90] ^ x[41];
  assign t[73] = t[91] ^ x[42];
  assign t[74] = t[92] ^ x[51];
  assign t[75] = t[93] ^ x[52];
  assign t[76] = (t[94] & ~t[96] & ~t[97] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & ~t[97] & ~t[98] & ~t[100]) | (t[94] & ~t[95] & ~t[96] & ~t[99] & ~t[100]) | (~t[94] & t[95] & t[96] & t[97] & ~t[100]) | (~t[94] & t[95] & t[98] & t[99] & ~t[100]) | (t[94] & ~t[96] & ~t[98] & t[100]) | (~t[94] & t[96] & t[98] & t[100]);
  assign t[77] = (t[94] & t[95] & ~t[96] & ~t[98] & t[99] & ~t[100]) | (t[94] & t[96] & ~t[97] & ~t[98] & ~t[99] & t[100]) | (~t[95] & ~t[96] & t[98] & ~t[99] & ~t[100]) | (~t[94] & ~t[96] & ~t[97] & t[98] & ~t[99]) | (~t[94] & ~t[95] & ~t[97] & t[98] & ~t[100]) | (~t[94] & ~t[96] & t[97] & t[98] & t[99]) | (t[97] & t[98] & ~t[99] & ~t[100]);
  assign t[78] = (t[101] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & ~t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[102] & ~t[103] & ~t[106] & ~t[107]) | (~t[101] & t[102] & t[103] & t[104] & ~t[107]) | (~t[101] & t[102] & t[105] & t[106] & ~t[107]) | (t[101] & ~t[103] & ~t[105] & t[107]) | (~t[101] & t[103] & t[105] & t[107]);
  assign t[79] = (t[101] & t[102] & ~t[103] & t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[103] & ~t[104] & t[105] & ~t[106] & t[107]) | (~t[102] & t[103] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[102] & t[103] & ~t[106] & ~t[107]) | (~t[101] & t[103] & t[104] & ~t[105] & t[106]) | (t[103] & ~t[104] & t[106] & ~t[107]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[81] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[82] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[83] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[84] = (t[102] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & t[102] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[102] & ~t[103] & ~t[106] & ~t[107]) | (t[101] & ~t[102] & t[103] & t[104] & ~t[107]) | (t[101] & ~t[102] & t[105] & t[106] & ~t[107]) | (t[102] & ~t[104] & ~t[106] & t[107]) | (~t[102] & t[104] & t[106] & t[107]);
  assign t[85] = (t[101] & t[102] & t[103] & ~t[104] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & ~t[104] & ~t[105] & t[106] & t[107]) | (~t[102] & ~t[103] & t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[103] & t[104] & ~t[106] & ~t[107]) | (~t[101] & ~t[102] & t[104] & ~t[105] & ~t[107]) | (~t[102] & t[103] & t[104] & t[105] & ~t[106]) | (~t[103] & t[104] & t[105] & ~t[107]);
  assign t[86] = (t[101] & t[102] & ~t[103] & ~t[105] & t[106] & ~t[107]) | (t[101] & t[103] & ~t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & t[105] & ~t[106] & ~t[107]) | (~t[101] & ~t[103] & ~t[104] & t[105] & ~t[106]) | (~t[101] & ~t[102] & ~t[104] & t[105] & ~t[107]) | (~t[101] & ~t[103] & t[104] & t[105] & t[106]) | (t[104] & t[105] & ~t[106] & ~t[107]);
  assign t[87] = (t[101] & t[102] & ~t[104] & t[105] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[104] & ~t[105] & t[106] & ~t[107]) | (~t[101] & ~t[102] & ~t[103] & t[106] & ~t[107]) | (~t[102] & t[103] & ~t[104] & t[105] & t[106]) | (t[103] & ~t[105] & t[106] & ~t[107]);
  assign t[88] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[89] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[8] = ~(t[11]);
  assign t[90] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[91] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[93] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[94] = t[129] ^ x[9];
  assign t[95] = t[130] ^ x[4];
  assign t[96] = t[131] ^ x[5];
  assign t[97] = t[132] ^ x[6];
  assign t[98] = t[133] ^ x[10];
  assign t[99] = t[134] ^ x[7];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind150(x, y);
 input [46:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[128] ^ x[22];
  assign t[101] = t[129] ^ x[23];
  assign t[102] = t[130] ^ x[27];
  assign t[103] = t[131] ^ x[24];
  assign t[104] = t[132] ^ x[25];
  assign t[105] = t[133] ^ x[33];
  assign t[106] = t[134] ^ x[39];
  assign t[107] = t[135] ^ x[34];
  assign t[108] = t[136] ^ x[40];
  assign t[109] = t[137] ^ x[41];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[138] ^ x[42];
  assign t[111] = t[139] ^ x[32];
  assign t[112] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[113] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[114] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[115] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[11] = ~(t[15]);
  assign t[120] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[121] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[122] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[123] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[124] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[125] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[126] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[127] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[128] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[129] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[133] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[134] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[135] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[136] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[137] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[138] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[139] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[43] | t[20]);
  assign t[15] = ~x[2] & t[44];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[45] | t[23]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[47]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[48]);
  assign t[22] = ~(t[49]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[50]);
  assign t[25] = ~(t[46] | t[47]);
  assign t[26] = ~(t[51]);
  assign t[27] = ~(t[48] | t[49]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~t[32];
  assign t[31] = ~(t[33] ^ t[34]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~t[35];
  assign t[34] = x[2] ? x[45] : t[36];
  assign t[35] = x[2] ? x[46] : t[37];
  assign t[36] = ~(t[38] & t[39]);
  assign t[37] = ~(t[40] & t[41]);
  assign t[38] = ~(t[19] & t[24]);
  assign t[39] = t[13] | t[43];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[22] & t[26]);
  assign t[41] = t[16] | t[45];
  assign t[42] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[43] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[44] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[45] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[46] = (t[54] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[54] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[47] = (t[54] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[54] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[48] = (t[58] & ~t[65] & ~t[67]) | (~t[64] & t[65] & ~t[66]) | (~t[58] & ~t[65] & t[67]) | (t[64] & t[65] & t[66]);
  assign t[49] = (t[58] & ~t[65] & ~t[66]) | (~t[64] & t[65] & ~t[67]) | (~t[58] & ~t[65] & t[66]) | (t[64] & t[65] & t[67]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[54] & ~t[62]) | (~t[54] & t[62]);
  assign t[51] = (t[58] & ~t[66]) | (~t[58] & t[66]);
  assign t[52] = t[68] ^ x[9];
  assign t[53] = t[69] ^ x[10];
  assign t[54] = t[70] ^ x[18];
  assign t[55] = t[71] ^ x[19];
  assign t[56] = t[72] ^ x[26];
  assign t[57] = t[73] ^ x[27];
  assign t[58] = t[74] ^ x[33];
  assign t[59] = t[75] ^ x[34];
  assign t[5] = ~(~x[2] & ~t[42]);
  assign t[60] = t[76] ^ x[35];
  assign t[61] = t[77] ^ x[36];
  assign t[62] = t[78] ^ x[37];
  assign t[63] = t[79] ^ x[38];
  assign t[64] = t[80] ^ x[39];
  assign t[65] = t[81] ^ x[40];
  assign t[66] = t[82] ^ x[41];
  assign t[67] = t[83] ^ x[42];
  assign t[68] = (t[84] & ~t[86] & ~t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[87] & ~t[88] & ~t[90]) | (t[84] & ~t[85] & ~t[86] & ~t[89] & ~t[90]) | (~t[84] & t[85] & t[86] & t[87] & ~t[90]) | (~t[84] & t[85] & t[88] & t[89] & ~t[90]) | (t[84] & ~t[86] & ~t[88] & t[90]) | (~t[84] & t[86] & t[88] & t[90]);
  assign t[69] = (t[84] & t[85] & ~t[86] & ~t[88] & t[89] & ~t[90]) | (t[84] & t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[90]) | (~t[84] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[84] & ~t[85] & ~t[87] & t[88] & ~t[90]) | (~t[84] & ~t[86] & t[87] & t[88] & t[89]) | (t[87] & t[88] & ~t[89] & ~t[90]);
  assign t[6] = ~t[9];
  assign t[70] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[71] = (t[91] & t[92] & ~t[93] & t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[93] & ~t[94] & t[95] & ~t[96] & t[97]) | (~t[92] & t[93] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[92] & t[93] & ~t[96] & ~t[97]) | (~t[91] & t[93] & t[94] & ~t[95] & t[96]) | (t[93] & ~t[94] & t[96] & ~t[97]);
  assign t[72] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[73] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[74] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[75] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[76] = (t[92] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & t[92] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[92] & ~t[93] & ~t[96] & ~t[97]) | (t[91] & ~t[92] & t[93] & t[94] & ~t[97]) | (t[91] & ~t[92] & t[95] & t[96] & ~t[97]) | (t[92] & ~t[94] & ~t[96] & t[97]) | (~t[92] & t[94] & t[96] & t[97]);
  assign t[77] = (t[91] & t[92] & t[93] & ~t[94] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[94] & ~t[95] & t[96] & t[97]) | (~t[92] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[93] & t[94] & ~t[96] & ~t[97]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[97]) | (~t[92] & t[93] & t[94] & t[95] & ~t[96]) | (~t[93] & t[94] & t[95] & ~t[97]);
  assign t[78] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[79] = (t[91] & t[92] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[91] & ~t[92] & ~t[93] & t[96] & ~t[97]) | (~t[92] & t[93] & ~t[94] & t[95] & t[96]) | (t[93] & ~t[95] & t[96] & ~t[97]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[81] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[82] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[83] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[84] = t[112] ^ x[9];
  assign t[85] = t[113] ^ x[4];
  assign t[86] = t[114] ^ x[5];
  assign t[87] = t[115] ^ x[6];
  assign t[88] = t[116] ^ x[10];
  assign t[89] = t[117] ^ x[7];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[8];
  assign t[91] = t[119] ^ x[18];
  assign t[92] = t[120] ^ x[35];
  assign t[93] = t[121] ^ x[19];
  assign t[94] = t[122] ^ x[36];
  assign t[95] = t[123] ^ x[37];
  assign t[96] = t[124] ^ x[38];
  assign t[97] = t[125] ^ x[17];
  assign t[98] = t[126] ^ x[26];
  assign t[99] = t[127] ^ x[21];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind151(x, y);
 input [54:0] x;
 output y;

 wire [161:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[19];
  assign t[101] = t[136] ^ x[53];
  assign t[102] = t[137] ^ x[20];
  assign t[103] = t[138] ^ x[21];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[17];
  assign t[106] = t[141] ^ x[29];
  assign t[107] = t[142] ^ x[24];
  assign t[108] = t[143] ^ x[25];
  assign t[109] = t[144] ^ x[26];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[145] ^ x[30];
  assign t[111] = t[146] ^ x[27];
  assign t[112] = t[147] ^ x[28];
  assign t[113] = t[148] ^ x[36];
  assign t[114] = t[149] ^ x[37];
  assign t[115] = t[150] ^ x[54];
  assign t[116] = t[151] ^ x[38];
  assign t[117] = t[152] ^ x[39];
  assign t[118] = t[153] ^ x[40];
  assign t[119] = t[154] ^ x[35];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[49];
  assign t[121] = t[156] ^ x[44];
  assign t[122] = t[157] ^ x[45];
  assign t[123] = t[158] ^ x[46];
  assign t[124] = t[159] ^ x[50];
  assign t[125] = t[160] ^ x[47];
  assign t[126] = t[161] ^ x[48];
  assign t[127] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[128] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[129] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[12] = ~(t[16] & t[17]);
  assign t[130] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[133] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[134] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[135] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[136] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[137] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[138] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[139] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[13] = ~(t[46] & t[18]);
  assign t[140] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[141] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[142] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[143] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[144] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[31] & ~x[32] & ~x[33]) | (~x[31] & x[32] & ~x[33]) | (~x[31] & ~x[32] & x[33]) | (x[31] & x[32] & x[33]);
  assign t[149] = (x[31] & ~x[32] & ~x[34]) | (~x[31] & x[32] & ~x[34]) | (~x[31] & ~x[32] & x[34]) | (x[31] & x[32] & x[34]);
  assign t[14] = ~(t[47] & t[19]);
  assign t[150] = (x[31] & ~x[33]) | (~x[31] & x[33]);
  assign t[151] = (x[31] & ~x[34]) | (~x[31] & x[34]);
  assign t[152] = (x[32] & ~x[33]) | (~x[32] & x[33]);
  assign t[153] = (x[32] & ~x[34]) | (~x[32] & x[34]);
  assign t[154] = (x[33] & ~x[34]) | (~x[33] & x[34]);
  assign t[155] = (x[43] & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0);
  assign t[156] = (x[43] & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0);
  assign t[157] = (x[43] & ~1'b0) | (~x[43] & 1'b0);
  assign t[158] = (x[43] & ~1'b0) | (~x[43] & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[48];
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[16] = ~(t[49] & t[20]);
  assign t[17] = ~(t[50] & t[21]);
  assign t[18] = ~(t[51]);
  assign t[19] = ~(t[51] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[52]);
  assign t[21] = ~(t[52] & t[23]);
  assign t[22] = ~(t[46]);
  assign t[23] = ~(t[49]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27];
  assign t[26] = ~(t[28] ^ t[29]);
  assign t[27] = ~(t[30] ^ t[31]);
  assign t[28] = t[8] ? x[42] : x[41];
  assign t[29] = ~x[2] & t[53];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[51] : t[33];
  assign t[32] = x[2] ? x[52] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[18] & t[39]);
  assign t[36] = ~(t[40] & t[54]);
  assign t[37] = ~(t[20] & t[41]);
  assign t[38] = ~(t[42] & t[55]);
  assign t[39] = ~(t[47]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[43] & t[22]);
  assign t[41] = ~(t[50]);
  assign t[42] = ~(t[44] & t[23]);
  assign t[43] = ~(t[47] & t[51]);
  assign t[44] = ~(t[50] & t[52]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[58] & ~t[60] & ~t[62]) | (~t[59] & t[60] & ~t[61]) | (~t[58] & ~t[60] & t[62]) | (t[59] & t[60] & t[61]);
  assign t[47] = (t[58] & ~t[61]) | (~t[58] & t[61]);
  assign t[48] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[49] = (t[65] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[65] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[65] & ~t[68]) | (~t[65] & t[68]);
  assign t[51] = (t[58] & ~t[60] & ~t[61]) | (~t[59] & t[60] & ~t[62]) | (~t[58] & ~t[60] & t[61]) | (t[59] & t[60] & t[62]);
  assign t[52] = (t[65] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[65] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[53] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[54] = (t[58] & ~t[72]) | (~t[58] & t[72]);
  assign t[55] = (t[65] & ~t[73]) | (~t[65] & t[73]);
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[10];
  assign t[58] = t[76] ^ x[18];
  assign t[59] = t[77] ^ x[19];
  assign t[5] = ~x[2] & t[45];
  assign t[60] = t[78] ^ x[20];
  assign t[61] = t[79] ^ x[21];
  assign t[62] = t[80] ^ x[22];
  assign t[63] = t[81] ^ x[29];
  assign t[64] = t[82] ^ x[30];
  assign t[65] = t[83] ^ x[36];
  assign t[66] = t[84] ^ x[37];
  assign t[67] = t[85] ^ x[38];
  assign t[68] = t[86] ^ x[39];
  assign t[69] = t[87] ^ x[40];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[49];
  assign t[71] = t[89] ^ x[50];
  assign t[72] = t[90] ^ x[53];
  assign t[73] = t[91] ^ x[54];
  assign t[74] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[78] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[79] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[82] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[83] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[84] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[85] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[86] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[87] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[89] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[8] = ~(t[11]);
  assign t[90] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = t[127] ^ x[9];
  assign t[93] = t[128] ^ x[4];
  assign t[94] = t[129] ^ x[5];
  assign t[95] = t[130] ^ x[6];
  assign t[96] = t[131] ^ x[10];
  assign t[97] = t[132] ^ x[7];
  assign t[98] = t[133] ^ x[8];
  assign t[99] = t[134] ^ x[18];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[24]) | (~t[0] & t[24]);
endmodule

module R2ind152(x, y);
 input [46:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[128] ^ x[25];
  assign t[101] = t[129] ^ x[26];
  assign t[102] = t[130] ^ x[30];
  assign t[103] = t[131] ^ x[27];
  assign t[104] = t[132] ^ x[28];
  assign t[105] = t[133] ^ x[36];
  assign t[106] = t[134] ^ x[37];
  assign t[107] = t[135] ^ x[46];
  assign t[108] = t[136] ^ x[38];
  assign t[109] = t[137] ^ x[39];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[138] ^ x[40];
  assign t[111] = t[139] ^ x[35];
  assign t[112] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[113] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[114] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[115] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[11] = ~(t[15]);
  assign t[120] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[121] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[122] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[123] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[124] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[125] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[127] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[128] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[129] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[12] = ~(t[16] & t[17]);
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[133] = (x[31] & ~x[32] & ~x[33]) | (~x[31] & x[32] & ~x[33]) | (~x[31] & ~x[32] & x[33]) | (x[31] & x[32] & x[33]);
  assign t[134] = (x[31] & ~x[32] & ~x[34]) | (~x[31] & x[32] & ~x[34]) | (~x[31] & ~x[32] & x[34]) | (x[31] & x[32] & x[34]);
  assign t[135] = (x[31] & ~x[33]) | (~x[31] & x[33]);
  assign t[136] = (x[31] & ~x[34]) | (~x[31] & x[34]);
  assign t[137] = (x[32] & ~x[33]) | (~x[32] & x[33]);
  assign t[138] = (x[32] & ~x[34]) | (~x[32] & x[34]);
  assign t[139] = (x[33] & ~x[34]) | (~x[33] & x[34]);
  assign t[13] = ~(t[43] & t[18]);
  assign t[14] = ~(t[44] & t[19]);
  assign t[15] = ~x[2] & t[45];
  assign t[16] = ~(t[46] & t[20]);
  assign t[17] = ~(t[47] & t[21]);
  assign t[18] = ~(t[48]);
  assign t[19] = ~(t[48] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[49]);
  assign t[21] = ~(t[49] & t[23]);
  assign t[22] = ~(t[43]);
  assign t[23] = ~(t[46]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27];
  assign t[26] = ~t[28];
  assign t[27] = ~(t[29] ^ t[30]);
  assign t[28] = t[8] ? x[42] : x[41];
  assign t[29] = ~t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = x[2] ? x[43] : t[32];
  assign t[31] = x[2] ? x[44] : t[33];
  assign t[32] = ~(t[34] & t[35]);
  assign t[33] = ~(t[36] & t[37]);
  assign t[34] = ~(t[18] & t[38]);
  assign t[35] = t[39] | t[50];
  assign t[36] = ~(t[20] & t[40]);
  assign t[37] = t[41] | t[51];
  assign t[38] = ~(t[44]);
  assign t[39] = ~(t[22] | t[18]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[47]);
  assign t[41] = ~(t[23] | t[20]);
  assign t[42] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[43] = (t[54] & ~t[56] & ~t[58]) | (~t[55] & t[56] & ~t[57]) | (~t[54] & ~t[56] & t[58]) | (t[55] & t[56] & t[57]);
  assign t[44] = (t[54] & ~t[57]) | (~t[54] & t[57]);
  assign t[45] = (t[59] & ~t[60]) | (~t[59] & t[60]);
  assign t[46] = (t[61] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[61] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[47] = (t[61] & ~t[64]) | (~t[61] & t[64]);
  assign t[48] = (t[54] & ~t[56] & ~t[57]) | (~t[55] & t[56] & ~t[58]) | (~t[54] & ~t[56] & t[57]) | (t[55] & t[56] & t[58]);
  assign t[49] = (t[61] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[61] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[54] & ~t[66]) | (~t[54] & t[66]);
  assign t[51] = (t[61] & ~t[67]) | (~t[61] & t[67]);
  assign t[52] = t[68] ^ x[9];
  assign t[53] = t[69] ^ x[10];
  assign t[54] = t[70] ^ x[18];
  assign t[55] = t[71] ^ x[19];
  assign t[56] = t[72] ^ x[20];
  assign t[57] = t[73] ^ x[21];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[29];
  assign t[5] = ~x[2] & t[42];
  assign t[60] = t[76] ^ x[30];
  assign t[61] = t[77] ^ x[36];
  assign t[62] = t[78] ^ x[37];
  assign t[63] = t[79] ^ x[38];
  assign t[64] = t[80] ^ x[39];
  assign t[65] = t[81] ^ x[40];
  assign t[66] = t[82] ^ x[45];
  assign t[67] = t[83] ^ x[46];
  assign t[68] = (t[84] & ~t[86] & ~t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[87] & ~t[88] & ~t[90]) | (t[84] & ~t[85] & ~t[86] & ~t[89] & ~t[90]) | (~t[84] & t[85] & t[86] & t[87] & ~t[90]) | (~t[84] & t[85] & t[88] & t[89] & ~t[90]) | (t[84] & ~t[86] & ~t[88] & t[90]) | (~t[84] & t[86] & t[88] & t[90]);
  assign t[69] = (t[84] & t[85] & ~t[86] & ~t[88] & t[89] & ~t[90]) | (t[84] & t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[90]) | (~t[84] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[84] & ~t[85] & ~t[87] & t[88] & ~t[90]) | (~t[84] & ~t[86] & t[87] & t[88] & t[89]) | (t[87] & t[88] & ~t[89] & ~t[90]);
  assign t[6] = ~t[9];
  assign t[70] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[71] = (t[92] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & t[92] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[92] & ~t[93] & ~t[96] & ~t[97]) | (t[91] & ~t[92] & t[93] & t[94] & ~t[97]) | (t[91] & ~t[92] & t[95] & t[96] & ~t[97]) | (t[92] & ~t[94] & ~t[96] & t[97]) | (~t[92] & t[94] & t[96] & t[97]);
  assign t[72] = (t[91] & t[92] & t[93] & ~t[94] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[94] & ~t[95] & t[96] & t[97]) | (~t[92] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[93] & t[94] & ~t[96] & ~t[97]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[97]) | (~t[92] & t[93] & t[94] & t[95] & ~t[96]) | (~t[93] & t[94] & t[95] & ~t[97]);
  assign t[73] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[74] = (t[91] & t[92] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[91] & ~t[92] & ~t[93] & t[96] & ~t[97]) | (~t[92] & t[93] & ~t[94] & t[95] & t[96]) | (t[93] & ~t[95] & t[96] & ~t[97]);
  assign t[75] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[76] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[77] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[78] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[79] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[81] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[82] = (t[91] & t[92] & ~t[93] & t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[93] & ~t[94] & t[95] & ~t[96] & t[97]) | (~t[92] & t[93] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[92] & t[93] & ~t[96] & ~t[97]) | (~t[91] & t[93] & t[94] & ~t[95] & t[96]) | (t[93] & ~t[94] & t[96] & ~t[97]);
  assign t[83] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[84] = t[112] ^ x[9];
  assign t[85] = t[113] ^ x[4];
  assign t[86] = t[114] ^ x[5];
  assign t[87] = t[115] ^ x[6];
  assign t[88] = t[116] ^ x[10];
  assign t[89] = t[117] ^ x[7];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[8];
  assign t[91] = t[119] ^ x[18];
  assign t[92] = t[120] ^ x[19];
  assign t[93] = t[121] ^ x[45];
  assign t[94] = t[122] ^ x[20];
  assign t[95] = t[123] ^ x[21];
  assign t[96] = t[124] ^ x[22];
  assign t[97] = t[125] ^ x[17];
  assign t[98] = t[126] ^ x[29];
  assign t[99] = t[127] ^ x[24];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[24]) | (~t[0] & t[24]);
endmodule

module R2ind153(x, y);
 input [46:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[128] ^ x[22];
  assign t[101] = t[129] ^ x[23];
  assign t[102] = t[130] ^ x[27];
  assign t[103] = t[131] ^ x[24];
  assign t[104] = t[132] ^ x[25];
  assign t[105] = t[133] ^ x[33];
  assign t[106] = t[134] ^ x[39];
  assign t[107] = t[135] ^ x[34];
  assign t[108] = t[136] ^ x[40];
  assign t[109] = t[137] ^ x[41];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[138] ^ x[42];
  assign t[111] = t[139] ^ x[32];
  assign t[112] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[113] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[114] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[115] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[116] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[11] = ~(t[15]);
  assign t[120] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[121] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[122] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[123] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[124] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[125] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[126] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[127] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[128] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[129] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[12] = ~(t[16] & t[17]);
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[133] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[134] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[135] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[136] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[137] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[138] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[139] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[43]);
  assign t[15] = ~x[2] & t[44];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[45]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[47]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[48]);
  assign t[22] = ~(t[49]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[47] & t[46]);
  assign t[25] = ~(t[50]);
  assign t[26] = ~(t[49] & t[48]);
  assign t[27] = ~(t[51]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~t[32];
  assign t[31] = ~(t[33] ^ t[34]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~t[35];
  assign t[34] = x[2] ? x[45] : t[36];
  assign t[35] = x[2] ? x[46] : t[37];
  assign t[36] = ~(t[13] & t[38]);
  assign t[37] = ~(t[16] & t[39]);
  assign t[38] = t[40] | t[43];
  assign t[39] = t[41] | t[45];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[25] | t[18]);
  assign t[41] = ~(t[27] | t[21]);
  assign t[42] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[43] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[44] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[45] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[46] = (t[54] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[54] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[47] = (t[54] & ~t[62]) | (~t[54] & t[62]);
  assign t[48] = (t[58] & ~t[65] & ~t[66]) | (~t[64] & t[65] & ~t[67]) | (~t[58] & ~t[65] & t[66]) | (t[64] & t[65] & t[67]);
  assign t[49] = (t[58] & ~t[66]) | (~t[58] & t[66]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[54] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[54] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[51] = (t[58] & ~t[65] & ~t[67]) | (~t[64] & t[65] & ~t[66]) | (~t[58] & ~t[65] & t[67]) | (t[64] & t[65] & t[66]);
  assign t[52] = t[68] ^ x[9];
  assign t[53] = t[69] ^ x[10];
  assign t[54] = t[70] ^ x[18];
  assign t[55] = t[71] ^ x[19];
  assign t[56] = t[72] ^ x[26];
  assign t[57] = t[73] ^ x[27];
  assign t[58] = t[74] ^ x[33];
  assign t[59] = t[75] ^ x[34];
  assign t[5] = ~x[2] & t[42];
  assign t[60] = t[76] ^ x[35];
  assign t[61] = t[77] ^ x[36];
  assign t[62] = t[78] ^ x[37];
  assign t[63] = t[79] ^ x[38];
  assign t[64] = t[80] ^ x[39];
  assign t[65] = t[81] ^ x[40];
  assign t[66] = t[82] ^ x[41];
  assign t[67] = t[83] ^ x[42];
  assign t[68] = (t[84] & ~t[86] & ~t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[87] & ~t[88] & ~t[90]) | (t[84] & ~t[85] & ~t[86] & ~t[89] & ~t[90]) | (~t[84] & t[85] & t[86] & t[87] & ~t[90]) | (~t[84] & t[85] & t[88] & t[89] & ~t[90]) | (t[84] & ~t[86] & ~t[88] & t[90]) | (~t[84] & t[86] & t[88] & t[90]);
  assign t[69] = (t[84] & t[85] & ~t[86] & ~t[88] & t[89] & ~t[90]) | (t[84] & t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[90]) | (~t[84] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[84] & ~t[85] & ~t[87] & t[88] & ~t[90]) | (~t[84] & ~t[86] & t[87] & t[88] & t[89]) | (t[87] & t[88] & ~t[89] & ~t[90]);
  assign t[6] = ~t[9];
  assign t[70] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[71] = (t[91] & t[92] & ~t[93] & t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[93] & ~t[94] & t[95] & ~t[96] & t[97]) | (~t[92] & t[93] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[92] & t[93] & ~t[96] & ~t[97]) | (~t[91] & t[93] & t[94] & ~t[95] & t[96]) | (t[93] & ~t[94] & t[96] & ~t[97]);
  assign t[72] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[73] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[74] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[75] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[76] = (t[92] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & t[92] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[92] & ~t[93] & ~t[96] & ~t[97]) | (t[91] & ~t[92] & t[93] & t[94] & ~t[97]) | (t[91] & ~t[92] & t[95] & t[96] & ~t[97]) | (t[92] & ~t[94] & ~t[96] & t[97]) | (~t[92] & t[94] & t[96] & t[97]);
  assign t[77] = (t[91] & t[92] & t[93] & ~t[94] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[94] & ~t[95] & t[96] & t[97]) | (~t[92] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[93] & t[94] & ~t[96] & ~t[97]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[97]) | (~t[92] & t[93] & t[94] & t[95] & ~t[96]) | (~t[93] & t[94] & t[95] & ~t[97]);
  assign t[78] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[79] = (t[91] & t[92] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[91] & ~t[92] & ~t[93] & t[96] & ~t[97]) | (~t[92] & t[93] & ~t[94] & t[95] & t[96]) | (t[93] & ~t[95] & t[96] & ~t[97]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[81] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[82] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[83] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[84] = t[112] ^ x[9];
  assign t[85] = t[113] ^ x[4];
  assign t[86] = t[114] ^ x[5];
  assign t[87] = t[115] ^ x[6];
  assign t[88] = t[116] ^ x[10];
  assign t[89] = t[117] ^ x[7];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[8];
  assign t[91] = t[119] ^ x[18];
  assign t[92] = t[120] ^ x[35];
  assign t[93] = t[121] ^ x[19];
  assign t[94] = t[122] ^ x[36];
  assign t[95] = t[123] ^ x[37];
  assign t[96] = t[124] ^ x[38];
  assign t[97] = t[125] ^ x[17];
  assign t[98] = t[126] ^ x[26];
  assign t[99] = t[127] ^ x[21];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind154(x, y);
 input [66:0] x;
 output y;

 wire [199:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[130] & ~t[132] & ~t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[133] & ~t[134] & ~t[136]) | (t[130] & ~t[131] & ~t[132] & ~t[135] & ~t[136]) | (~t[130] & t[131] & t[132] & t[133] & ~t[136]) | (~t[130] & t[131] & t[134] & t[135] & ~t[136]) | (t[130] & ~t[132] & ~t[134] & t[136]) | (~t[130] & t[132] & t[134] & t[136]);
  assign t[101] = (t[130] & t[131] & ~t[132] & ~t[134] & t[135] & ~t[136]) | (t[130] & t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[136]) | (~t[130] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[130] & ~t[131] & ~t[133] & t[134] & ~t[136]) | (~t[130] & ~t[132] & t[133] & t[134] & t[135]) | (t[133] & t[134] & ~t[135] & ~t[136]);
  assign t[102] = (t[137] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & ~t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[138] & ~t[139] & ~t[142] & ~t[143]) | (~t[137] & t[138] & t[139] & t[140] & ~t[143]) | (~t[137] & t[138] & t[141] & t[142] & ~t[143]) | (t[137] & ~t[139] & ~t[141] & t[143]) | (~t[137] & t[139] & t[141] & t[143]);
  assign t[103] = (t[137] & t[138] & ~t[139] & t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[139] & ~t[140] & t[141] & ~t[142] & t[143]) | (~t[138] & t[139] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[138] & t[139] & ~t[142] & ~t[143]) | (~t[137] & t[139] & t[140] & ~t[141] & t[142]) | (t[139] & ~t[140] & t[142] & ~t[143]);
  assign t[104] = (t[124] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & t[124] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[124] & ~t[125] & ~t[128] & ~t[129]) | (t[123] & ~t[124] & t[125] & t[126] & ~t[129]) | (t[123] & ~t[124] & t[127] & t[128] & ~t[129]) | (t[124] & ~t[126] & ~t[128] & t[129]) | (~t[124] & t[126] & t[128] & t[129]);
  assign t[105] = (t[123] & t[124] & t[125] & ~t[126] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[126] & ~t[127] & t[128] & t[129]) | (~t[124] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[125] & t[126] & ~t[128] & ~t[129]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[129]) | (~t[124] & t[125] & t[126] & t[127] & ~t[128]) | (~t[125] & t[126] & t[127] & ~t[129]);
  assign t[106] = (t[123] & t[124] & ~t[125] & ~t[127] & t[128] & ~t[129]) | (t[123] & t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[129]) | (~t[123] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[123] & ~t[124] & ~t[126] & t[127] & ~t[129]) | (~t[123] & ~t[125] & t[126] & t[127] & t[128]) | (t[126] & t[127] & ~t[128] & ~t[129]);
  assign t[107] = (t[123] & t[124] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[123] & ~t[124] & ~t[125] & t[128] & ~t[129]) | (~t[124] & t[125] & ~t[126] & t[127] & t[128]) | (t[125] & ~t[127] & t[128] & ~t[129]);
  assign t[108] = (t[138] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & t[138] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[138] & ~t[139] & ~t[142] & ~t[143]) | (t[137] & ~t[138] & t[139] & t[140] & ~t[143]) | (t[137] & ~t[138] & t[141] & t[142] & ~t[143]) | (t[138] & ~t[140] & ~t[142] & t[143]) | (~t[138] & t[140] & t[142] & t[143]);
  assign t[109] = (t[137] & t[138] & t[139] & ~t[140] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[140] & ~t[141] & t[142] & t[143]) | (~t[138] & ~t[139] & t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[139] & t[140] & ~t[142] & ~t[143]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[143]) | (~t[138] & t[139] & t[140] & t[141] & ~t[142]) | (~t[139] & t[140] & t[141] & ~t[143]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (t[137] & t[138] & ~t[139] & ~t[141] & t[142] & ~t[143]) | (t[137] & t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[143]) | (~t[137] & ~t[139] & ~t[140] & t[141] & ~t[142]) | (~t[137] & ~t[138] & ~t[140] & t[141] & ~t[143]) | (~t[137] & ~t[139] & t[140] & t[141] & t[142]) | (t[140] & t[141] & ~t[142] & ~t[143]);
  assign t[111] = (t[137] & t[138] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[137] & ~t[138] & ~t[139] & t[142] & ~t[143]) | (~t[138] & t[139] & ~t[140] & t[141] & t[142]) | (t[139] & ~t[141] & t[142] & ~t[143]);
  assign t[112] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[113] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[114] = (t[151] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & ~t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[152] & ~t[153] & ~t[156] & ~t[157]) | (~t[151] & t[152] & t[153] & t[154] & ~t[157]) | (~t[151] & t[152] & t[155] & t[156] & ~t[157]) | (t[151] & ~t[153] & ~t[155] & t[157]) | (~t[151] & t[153] & t[155] & t[157]);
  assign t[115] = (t[151] & t[152] & ~t[153] & ~t[155] & t[156] & ~t[157]) | (t[151] & t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[157]) | (~t[151] & ~t[153] & ~t[154] & t[155] & ~t[156]) | (~t[151] & ~t[152] & ~t[154] & t[155] & ~t[157]) | (~t[151] & ~t[153] & t[154] & t[155] & t[156]) | (t[154] & t[155] & ~t[156] & ~t[157]);
  assign t[116] = t[158] ^ x[9];
  assign t[117] = t[159] ^ x[4];
  assign t[118] = t[160] ^ x[5];
  assign t[119] = t[161] ^ x[6];
  assign t[11] = ~(t[15]);
  assign t[120] = t[162] ^ x[10];
  assign t[121] = t[163] ^ x[7];
  assign t[122] = t[164] ^ x[8];
  assign t[123] = t[165] ^ x[18];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[19];
  assign t[126] = t[168] ^ x[36];
  assign t[127] = t[169] ^ x[37];
  assign t[128] = t[170] ^ x[38];
  assign t[129] = t[171] ^ x[17];
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = t[172] ^ x[26];
  assign t[131] = t[173] ^ x[21];
  assign t[132] = t[174] ^ x[22];
  assign t[133] = t[175] ^ x[23];
  assign t[134] = t[176] ^ x[27];
  assign t[135] = t[177] ^ x[24];
  assign t[136] = t[178] ^ x[25];
  assign t[137] = t[179] ^ x[33];
  assign t[138] = t[180] ^ x[39];
  assign t[139] = t[181] ^ x[34];
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = t[182] ^ x[40];
  assign t[141] = t[183] ^ x[41];
  assign t[142] = t[184] ^ x[42];
  assign t[143] = t[185] ^ x[32];
  assign t[144] = t[186] ^ x[51];
  assign t[145] = t[187] ^ x[46];
  assign t[146] = t[188] ^ x[47];
  assign t[147] = t[189] ^ x[48];
  assign t[148] = t[190] ^ x[52];
  assign t[149] = t[191] ^ x[49];
  assign t[14] = ~(t[65] | t[20]);
  assign t[150] = t[192] ^ x[50];
  assign t[151] = t[193] ^ x[63];
  assign t[152] = t[194] ^ x[58];
  assign t[153] = t[195] ^ x[59];
  assign t[154] = t[196] ^ x[60];
  assign t[155] = t[197] ^ x[64];
  assign t[156] = t[198] ^ x[61];
  assign t[157] = t[199] ^ x[62];
  assign t[158] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[159] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[66];
  assign t[160] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[161] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[164] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[165] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[166] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[167] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[168] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[169] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[16] = ~(t[21] | t[22]);
  assign t[170] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[171] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[172] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[173] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[174] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[175] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[176] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[177] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[178] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[179] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[17] = ~(t[67] | t[23]);
  assign t[180] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[181] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[182] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[183] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[184] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[185] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[186] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[187] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[188] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[189] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[18] = ~(t[68]);
  assign t[190] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[192] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[193] = (x[57] & ~1'b0 & ~1'b0) | (~x[57] & 1'b0 & ~1'b0) | (~x[57] & ~1'b0 & 1'b0) | (x[57] & 1'b0 & 1'b0);
  assign t[194] = (x[57] & ~1'b0 & ~1'b0) | (~x[57] & 1'b0 & ~1'b0) | (~x[57] & ~1'b0 & 1'b0) | (x[57] & 1'b0 & 1'b0);
  assign t[195] = (x[57] & ~1'b0) | (~x[57] & 1'b0);
  assign t[196] = (x[57] & ~1'b0) | (~x[57] & 1'b0);
  assign t[197] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[198] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[199] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = ~(t[69]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[70]);
  assign t[22] = ~(t[71]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[72]);
  assign t[25] = ~(t[68] | t[69]);
  assign t[26] = ~(t[73]);
  assign t[27] = ~(t[70] | t[71]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[74];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[68] & t[19]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[72] & t[43]);
  assign t[41] = ~(t[70] & t[22]);
  assign t[42] = ~(t[73] & t[44]);
  assign t[43] = ~(t[69] & t[18]);
  assign t[44] = ~(t[71] & t[21]);
  assign t[45] = ~(t[46] ^ t[47]);
  assign t[46] = t[48];
  assign t[47] = ~(t[49] ^ t[50]);
  assign t[48] = ~(t[51] ^ t[52]);
  assign t[49] = t[8] ? x[56] : x[55];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = ~x[2] & t[75];
  assign t[51] = ~t[53];
  assign t[52] = x[2] ? x[65] : t[54];
  assign t[53] = x[2] ? x[66] : t[55];
  assign t[54] = ~(t[56] & t[57]);
  assign t[55] = ~(t[58] & t[59]);
  assign t[56] = ~(t[19] & t[24]);
  assign t[57] = ~(t[60] & t[65]);
  assign t[58] = ~(t[22] & t[26]);
  assign t[59] = ~(t[61] & t[67]);
  assign t[5] = ~(~x[2] & ~t[64]);
  assign t[60] = ~(t[62] & t[18]);
  assign t[61] = ~(t[63] & t[21]);
  assign t[62] = ~(t[72] & t[69]);
  assign t[63] = ~(t[73] & t[71]);
  assign t[64] = (t[76] & ~t[77]) | (~t[76] & t[77]);
  assign t[65] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[66] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[67] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[68] = (t[78] & ~t[85] & ~t[87]) | (~t[84] & t[85] & ~t[86]) | (~t[78] & ~t[85] & t[87]) | (t[84] & t[85] & t[86]);
  assign t[69] = (t[78] & ~t[85] & ~t[86]) | (~t[84] & t[85] & ~t[87]) | (~t[78] & ~t[85] & t[86]) | (t[84] & t[85] & t[87]);
  assign t[6] = ~t[9];
  assign t[70] = (t[82] & ~t[89] & ~t[91]) | (~t[88] & t[89] & ~t[90]) | (~t[82] & ~t[89] & t[91]) | (t[88] & t[89] & t[90]);
  assign t[71] = (t[82] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[91]) | (~t[82] & ~t[89] & t[90]) | (t[88] & t[89] & t[91]);
  assign t[72] = (t[78] & ~t[86]) | (~t[78] & t[86]);
  assign t[73] = (t[82] & ~t[90]) | (~t[82] & t[90]);
  assign t[74] = (t[92] & ~t[93]) | (~t[92] & t[93]);
  assign t[75] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[76] = t[96] ^ x[9];
  assign t[77] = t[97] ^ x[10];
  assign t[78] = t[98] ^ x[18];
  assign t[79] = t[99] ^ x[19];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[26];
  assign t[81] = t[101] ^ x[27];
  assign t[82] = t[102] ^ x[33];
  assign t[83] = t[103] ^ x[34];
  assign t[84] = t[104] ^ x[35];
  assign t[85] = t[105] ^ x[36];
  assign t[86] = t[106] ^ x[37];
  assign t[87] = t[107] ^ x[38];
  assign t[88] = t[108] ^ x[39];
  assign t[89] = t[109] ^ x[40];
  assign t[8] = ~(t[11]);
  assign t[90] = t[110] ^ x[41];
  assign t[91] = t[111] ^ x[42];
  assign t[92] = t[112] ^ x[51];
  assign t[93] = t[113] ^ x[52];
  assign t[94] = t[114] ^ x[63];
  assign t[95] = t[115] ^ x[64];
  assign t[96] = (t[116] & ~t[118] & ~t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[119] & ~t[120] & ~t[122]) | (t[116] & ~t[117] & ~t[118] & ~t[121] & ~t[122]) | (~t[116] & t[117] & t[118] & t[119] & ~t[122]) | (~t[116] & t[117] & t[120] & t[121] & ~t[122]) | (t[116] & ~t[118] & ~t[120] & t[122]) | (~t[116] & t[118] & t[120] & t[122]);
  assign t[97] = (t[116] & t[117] & ~t[118] & ~t[120] & t[121] & ~t[122]) | (t[116] & t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[122]) | (~t[116] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[116] & ~t[117] & ~t[119] & t[120] & ~t[122]) | (~t[116] & ~t[118] & t[119] & t[120] & t[121]) | (t[119] & t[120] & ~t[121] & ~t[122]);
  assign t[98] = (t[123] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[124] & ~t[125] & ~t[128] & ~t[129]) | (~t[123] & t[124] & t[125] & t[126] & ~t[129]) | (~t[123] & t[124] & t[127] & t[128] & ~t[129]) | (t[123] & ~t[125] & ~t[127] & t[129]) | (~t[123] & t[125] & t[127] & t[129]);
  assign t[99] = (t[123] & t[124] & ~t[125] & t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[125] & ~t[126] & t[127] & ~t[128] & t[129]) | (~t[124] & t[125] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[124] & t[125] & ~t[128] & ~t[129]) | (~t[123] & t[125] & t[126] & ~t[127] & t[128]) | (t[125] & ~t[126] & t[128] & ~t[129]);
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28] & ~t[45]) | (~t[0] & t[28] & ~t[45]) | (~t[0] & ~t[28] & t[45]) | (t[0] & t[28] & t[45]);
endmodule

module R2ind155(x, y);
 input [66:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[120] & ~t[121] & ~t[122] & ~t[123] & ~t[124]) | (~t[119] & t[120] & ~t[122] & ~t[123] & ~t[125]) | (~t[119] & t[120] & ~t[121] & ~t[124] & ~t[125]) | (t[119] & ~t[120] & t[121] & t[122] & ~t[125]) | (t[119] & ~t[120] & t[123] & t[124] & ~t[125]) | (t[120] & ~t[122] & ~t[124] & t[125]) | (~t[120] & t[122] & t[124] & t[125]);
  assign t[101] = (t[119] & t[120] & t[121] & ~t[122] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[122] & ~t[123] & t[124] & t[125]) | (~t[120] & ~t[121] & t[122] & ~t[123] & ~t[124]) | (~t[119] & ~t[121] & t[122] & ~t[124] & ~t[125]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[125]) | (~t[120] & t[121] & t[122] & t[123] & ~t[124]) | (~t[121] & t[122] & t[123] & ~t[125]);
  assign t[102] = (t[119] & t[120] & ~t[121] & ~t[123] & t[124] & ~t[125]) | (t[119] & t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[125]) | (~t[119] & ~t[121] & ~t[122] & t[123] & ~t[124]) | (~t[119] & ~t[120] & ~t[122] & t[123] & ~t[125]) | (~t[119] & ~t[121] & t[122] & t[123] & t[124]) | (t[122] & t[123] & ~t[124] & ~t[125]);
  assign t[103] = (t[119] & t[120] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[119] & ~t[120] & ~t[121] & t[124] & ~t[125]) | (~t[120] & t[121] & ~t[122] & t[123] & t[124]) | (t[121] & ~t[123] & t[124] & ~t[125]);
  assign t[104] = (t[134] & ~t[135] & ~t[136] & ~t[137] & ~t[138]) | (~t[133] & t[134] & ~t[136] & ~t[137] & ~t[139]) | (~t[133] & t[134] & ~t[135] & ~t[138] & ~t[139]) | (t[133] & ~t[134] & t[135] & t[136] & ~t[139]) | (t[133] & ~t[134] & t[137] & t[138] & ~t[139]) | (t[134] & ~t[136] & ~t[138] & t[139]) | (~t[134] & t[136] & t[138] & t[139]);
  assign t[105] = (t[133] & t[134] & t[135] & ~t[136] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[136] & ~t[137] & t[138] & t[139]) | (~t[134] & ~t[135] & t[136] & ~t[137] & ~t[138]) | (~t[133] & ~t[135] & t[136] & ~t[138] & ~t[139]) | (~t[133] & ~t[134] & t[136] & ~t[137] & ~t[139]) | (~t[134] & t[135] & t[136] & t[137] & ~t[138]) | (~t[135] & t[136] & t[137] & ~t[139]);
  assign t[106] = (t[133] & t[134] & ~t[135] & ~t[137] & t[138] & ~t[139]) | (t[133] & t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[139]) | (~t[133] & ~t[135] & ~t[136] & t[137] & ~t[138]) | (~t[133] & ~t[134] & ~t[136] & t[137] & ~t[139]) | (~t[133] & ~t[135] & t[136] & t[137] & t[138]) | (t[136] & t[137] & ~t[138] & ~t[139]);
  assign t[107] = (t[133] & t[134] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[135] & ~t[136] & ~t[137] & t[138]) | (~t[133] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[133] & ~t[134] & ~t[135] & t[138] & ~t[139]) | (~t[134] & t[135] & ~t[136] & t[137] & t[138]) | (t[135] & ~t[137] & t[138] & ~t[139]);
  assign t[108] = (t[140] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (t[140] & ~t[141] & ~t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[141] & ~t[142] & ~t[145] & ~t[146]) | (~t[140] & t[141] & t[142] & t[143] & ~t[146]) | (~t[140] & t[141] & t[144] & t[145] & ~t[146]) | (t[140] & ~t[142] & ~t[144] & t[146]) | (~t[140] & t[142] & t[144] & t[146]);
  assign t[109] = (t[140] & t[141] & ~t[142] & ~t[144] & t[145] & ~t[146]) | (t[140] & t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[146]) | (~t[140] & ~t[142] & ~t[143] & t[144] & ~t[145]) | (~t[140] & ~t[141] & ~t[143] & t[144] & ~t[146]) | (~t[140] & ~t[142] & t[143] & t[144] & t[145]) | (t[143] & t[144] & ~t[145] & ~t[146]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (t[147] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (t[147] & ~t[148] & ~t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[148] & ~t[149] & ~t[152] & ~t[153]) | (~t[147] & t[148] & t[149] & t[150] & ~t[153]) | (~t[147] & t[148] & t[151] & t[152] & ~t[153]) | (t[147] & ~t[149] & ~t[151] & t[153]) | (~t[147] & t[149] & t[151] & t[153]);
  assign t[111] = (t[147] & t[148] & ~t[149] & ~t[151] & t[152] & ~t[153]) | (t[147] & t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[153]) | (~t[147] & ~t[149] & ~t[150] & t[151] & ~t[152]) | (~t[147] & ~t[148] & ~t[150] & t[151] & ~t[153]) | (~t[147] & ~t[149] & t[150] & t[151] & t[152]) | (t[150] & t[151] & ~t[152] & ~t[153]);
  assign t[112] = t[154] ^ x[9];
  assign t[113] = t[155] ^ x[4];
  assign t[114] = t[156] ^ x[5];
  assign t[115] = t[157] ^ x[6];
  assign t[116] = t[158] ^ x[10];
  assign t[117] = t[159] ^ x[7];
  assign t[118] = t[160] ^ x[8];
  assign t[119] = t[161] ^ x[18];
  assign t[11] = ~(t[15]);
  assign t[120] = t[162] ^ x[35];
  assign t[121] = t[163] ^ x[19];
  assign t[122] = t[164] ^ x[36];
  assign t[123] = t[165] ^ x[37];
  assign t[124] = t[166] ^ x[38];
  assign t[125] = t[167] ^ x[17];
  assign t[126] = t[168] ^ x[26];
  assign t[127] = t[169] ^ x[21];
  assign t[128] = t[170] ^ x[22];
  assign t[129] = t[171] ^ x[23];
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = t[172] ^ x[27];
  assign t[131] = t[173] ^ x[24];
  assign t[132] = t[174] ^ x[25];
  assign t[133] = t[175] ^ x[33];
  assign t[134] = t[176] ^ x[39];
  assign t[135] = t[177] ^ x[34];
  assign t[136] = t[178] ^ x[40];
  assign t[137] = t[179] ^ x[41];
  assign t[138] = t[180] ^ x[42];
  assign t[139] = t[181] ^ x[32];
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = t[182] ^ x[51];
  assign t[141] = t[183] ^ x[46];
  assign t[142] = t[184] ^ x[47];
  assign t[143] = t[185] ^ x[48];
  assign t[144] = t[186] ^ x[52];
  assign t[145] = t[187] ^ x[49];
  assign t[146] = t[188] ^ x[50];
  assign t[147] = t[189] ^ x[63];
  assign t[148] = t[190] ^ x[58];
  assign t[149] = t[191] ^ x[59];
  assign t[14] = ~(t[61] | t[20]);
  assign t[150] = t[192] ^ x[60];
  assign t[151] = t[193] ^ x[64];
  assign t[152] = t[194] ^ x[61];
  assign t[153] = t[195] ^ x[62];
  assign t[154] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[155] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[156] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[157] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[158] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[62];
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[162] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[163] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[164] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[165] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[166] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[167] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[168] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[169] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[16] = ~(t[21] | t[22]);
  assign t[170] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[171] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[172] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[174] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[175] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[176] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[177] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[178] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[179] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[17] = ~(t[63] | t[23]);
  assign t[180] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[181] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[182] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[183] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[184] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[185] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[186] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[187] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[188] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[189] = (x[57] & ~1'b0 & ~1'b0) | (~x[57] & 1'b0 & ~1'b0) | (~x[57] & ~1'b0 & 1'b0) | (x[57] & 1'b0 & 1'b0);
  assign t[18] = ~(t[64]);
  assign t[190] = (x[57] & ~1'b0 & ~1'b0) | (~x[57] & 1'b0 & ~1'b0) | (~x[57] & ~1'b0 & 1'b0) | (x[57] & 1'b0 & 1'b0);
  assign t[191] = (x[57] & ~1'b0) | (~x[57] & 1'b0);
  assign t[192] = (x[57] & ~1'b0) | (~x[57] & 1'b0);
  assign t[193] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[194] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[195] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = ~(t[65]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[66]);
  assign t[22] = ~(t[67]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[68]);
  assign t[25] = ~(t[64] | t[65]);
  assign t[26] = ~(t[69]);
  assign t[27] = ~(t[66] | t[67]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[70];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[64] & t[19]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[68] & t[43]);
  assign t[41] = ~(t[66] & t[22]);
  assign t[42] = ~(t[69] & t[44]);
  assign t[43] = ~(t[65] & t[18]);
  assign t[44] = ~(t[67] & t[21]);
  assign t[45] = ~(t[46] ^ t[47]);
  assign t[46] = t[48];
  assign t[47] = ~(t[49] ^ t[50]);
  assign t[48] = ~(t[51] ^ t[52]);
  assign t[49] = t[8] ? x[56] : x[55];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = ~x[2] & t[71];
  assign t[51] = ~t[53];
  assign t[52] = x[2] ? x[65] : t[54];
  assign t[53] = x[2] ? x[66] : t[55];
  assign t[54] = ~(t[56] & t[57]);
  assign t[55] = ~(t[58] & t[59]);
  assign t[56] = ~(t[19] & t[24]);
  assign t[57] = t[13] | t[61];
  assign t[58] = ~(t[22] & t[26]);
  assign t[59] = t[16] | t[63];
  assign t[5] = ~(~x[2] & ~t[60]);
  assign t[60] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[61] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[62] = (t[76] & ~t[77]) | (~t[76] & t[77]);
  assign t[63] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[64] = (t[74] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[74] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[65] = (t[74] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[74] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[66] = (t[78] & ~t[85] & ~t[87]) | (~t[84] & t[85] & ~t[86]) | (~t[78] & ~t[85] & t[87]) | (t[84] & t[85] & t[86]);
  assign t[67] = (t[78] & ~t[85] & ~t[86]) | (~t[84] & t[85] & ~t[87]) | (~t[78] & ~t[85] & t[86]) | (t[84] & t[85] & t[87]);
  assign t[68] = (t[74] & ~t[82]) | (~t[74] & t[82]);
  assign t[69] = (t[78] & ~t[86]) | (~t[78] & t[86]);
  assign t[6] = ~t[9];
  assign t[70] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[71] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[72] = t[92] ^ x[9];
  assign t[73] = t[93] ^ x[10];
  assign t[74] = t[94] ^ x[18];
  assign t[75] = t[95] ^ x[19];
  assign t[76] = t[96] ^ x[26];
  assign t[77] = t[97] ^ x[27];
  assign t[78] = t[98] ^ x[33];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[35];
  assign t[81] = t[101] ^ x[36];
  assign t[82] = t[102] ^ x[37];
  assign t[83] = t[103] ^ x[38];
  assign t[84] = t[104] ^ x[39];
  assign t[85] = t[105] ^ x[40];
  assign t[86] = t[106] ^ x[41];
  assign t[87] = t[107] ^ x[42];
  assign t[88] = t[108] ^ x[51];
  assign t[89] = t[109] ^ x[52];
  assign t[8] = ~(t[11]);
  assign t[90] = t[110] ^ x[63];
  assign t[91] = t[111] ^ x[64];
  assign t[92] = (t[112] & ~t[114] & ~t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[115] & ~t[116] & ~t[118]) | (t[112] & ~t[113] & ~t[114] & ~t[117] & ~t[118]) | (~t[112] & t[113] & t[114] & t[115] & ~t[118]) | (~t[112] & t[113] & t[116] & t[117] & ~t[118]) | (t[112] & ~t[114] & ~t[116] & t[118]) | (~t[112] & t[114] & t[116] & t[118]);
  assign t[93] = (t[112] & t[113] & ~t[114] & ~t[116] & t[117] & ~t[118]) | (t[112] & t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[118]) | (~t[112] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[112] & ~t[113] & ~t[115] & t[116] & ~t[118]) | (~t[112] & ~t[114] & t[115] & t[116] & t[117]) | (t[115] & t[116] & ~t[117] & ~t[118]);
  assign t[94] = (t[119] & ~t[121] & ~t[122] & ~t[123] & ~t[124]) | (t[119] & ~t[120] & ~t[122] & ~t[123] & ~t[125]) | (t[119] & ~t[120] & ~t[121] & ~t[124] & ~t[125]) | (~t[119] & t[120] & t[121] & t[122] & ~t[125]) | (~t[119] & t[120] & t[123] & t[124] & ~t[125]) | (t[119] & ~t[121] & ~t[123] & t[125]) | (~t[119] & t[121] & t[123] & t[125]);
  assign t[95] = (t[119] & t[120] & ~t[121] & t[122] & ~t[123] & ~t[125]) | (t[119] & ~t[121] & ~t[122] & t[123] & ~t[124] & t[125]) | (~t[120] & t[121] & ~t[122] & ~t[123] & ~t[125]) | (~t[119] & t[121] & ~t[122] & ~t[123] & ~t[124]) | (~t[119] & ~t[120] & t[121] & ~t[124] & ~t[125]) | (~t[119] & t[121] & t[122] & ~t[123] & t[124]) | (t[121] & ~t[122] & t[124] & ~t[125]);
  assign t[96] = (t[126] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & ~t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[127] & ~t[128] & ~t[131] & ~t[132]) | (~t[126] & t[127] & t[128] & t[129] & ~t[132]) | (~t[126] & t[127] & t[130] & t[131] & ~t[132]) | (t[126] & ~t[128] & ~t[130] & t[132]) | (~t[126] & t[128] & t[130] & t[132]);
  assign t[97] = (t[126] & t[127] & ~t[128] & ~t[130] & t[131] & ~t[132]) | (t[126] & t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[132]) | (~t[126] & ~t[128] & ~t[129] & t[130] & ~t[131]) | (~t[126] & ~t[127] & ~t[129] & t[130] & ~t[132]) | (~t[126] & ~t[128] & t[129] & t[130] & t[131]) | (t[129] & t[130] & ~t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[135] & ~t[136] & ~t[137] & ~t[138]) | (t[133] & ~t[134] & ~t[136] & ~t[137] & ~t[139]) | (t[133] & ~t[134] & ~t[135] & ~t[138] & ~t[139]) | (~t[133] & t[134] & t[135] & t[136] & ~t[139]) | (~t[133] & t[134] & t[137] & t[138] & ~t[139]) | (t[133] & ~t[135] & ~t[137] & t[139]) | (~t[133] & t[135] & t[137] & t[139]);
  assign t[99] = (t[133] & t[134] & ~t[135] & t[136] & ~t[137] & ~t[139]) | (t[133] & ~t[135] & ~t[136] & t[137] & ~t[138] & t[139]) | (~t[134] & t[135] & ~t[136] & ~t[137] & ~t[139]) | (~t[133] & t[135] & ~t[136] & ~t[137] & ~t[138]) | (~t[133] & ~t[134] & t[135] & ~t[138] & ~t[139]) | (~t[133] & t[135] & t[136] & ~t[137] & t[138]) | (t[135] & ~t[136] & t[138] & ~t[139]);
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28] & ~t[45]) | (~t[0] & t[28] & ~t[45]) | (~t[0] & ~t[28] & t[45]) | (t[0] & t[28] & t[45]);
endmodule

module R2ind156(x, y);
 input [54:0] x;
 output y;

 wire [163:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[8];
  assign t[101] = t[136] ^ x[18];
  assign t[102] = t[137] ^ x[35];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[36];
  assign t[105] = t[140] ^ x[37];
  assign t[106] = t[141] ^ x[38];
  assign t[107] = t[142] ^ x[17];
  assign t[108] = t[143] ^ x[26];
  assign t[109] = t[144] ^ x[21];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[145] ^ x[22];
  assign t[111] = t[146] ^ x[23];
  assign t[112] = t[147] ^ x[27];
  assign t[113] = t[148] ^ x[24];
  assign t[114] = t[149] ^ x[25];
  assign t[115] = t[150] ^ x[33];
  assign t[116] = t[151] ^ x[39];
  assign t[117] = t[152] ^ x[34];
  assign t[118] = t[153] ^ x[40];
  assign t[119] = t[154] ^ x[41];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[42];
  assign t[121] = t[156] ^ x[32];
  assign t[122] = t[157] ^ x[51];
  assign t[123] = t[158] ^ x[46];
  assign t[124] = t[159] ^ x[47];
  assign t[125] = t[160] ^ x[48];
  assign t[126] = t[161] ^ x[52];
  assign t[127] = t[162] ^ x[49];
  assign t[128] = t[163] ^ x[50];
  assign t[129] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[131] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[132] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[133] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[134] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[135] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[136] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[137] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[138] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[139] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[141] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[142] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[143] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[144] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[145] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[146] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[149] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = ~(t[48] | t[20]);
  assign t[150] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[151] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[152] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[153] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[154] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[155] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[156] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[157] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[158] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[159] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[15] = ~x[2] & t[49];
  assign t[160] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[50] | t[23]);
  assign t[18] = ~(t[51]);
  assign t[19] = ~(t[52]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[53]);
  assign t[22] = ~(t[54]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[55]);
  assign t[25] = ~(t[51] | t[52]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] | t[54]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[57];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[19] & t[24]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[43] & t[48]);
  assign t[41] = ~(t[22] & t[26]);
  assign t[42] = ~(t[44] & t[50]);
  assign t[43] = ~(t[45] & t[18]);
  assign t[44] = ~(t[46] & t[21]);
  assign t[45] = ~(t[55] & t[52]);
  assign t[46] = ~(t[56] & t[54]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[49] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[60] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[60] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[52] = (t[60] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[60] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[53] = (t[64] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[64] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[54] = (t[64] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[64] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[55] = (t[60] & ~t[68]) | (~t[60] & t[68]);
  assign t[56] = (t[64] & ~t[72]) | (~t[64] & t[72]);
  assign t[57] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[58] = t[76] ^ x[9];
  assign t[59] = t[77] ^ x[10];
  assign t[5] = ~(~x[2] & ~t[47]);
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[26];
  assign t[63] = t[81] ^ x[27];
  assign t[64] = t[82] ^ x[33];
  assign t[65] = t[83] ^ x[34];
  assign t[66] = t[84] ^ x[35];
  assign t[67] = t[85] ^ x[36];
  assign t[68] = t[86] ^ x[37];
  assign t[69] = t[87] ^ x[38];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[39];
  assign t[71] = t[89] ^ x[40];
  assign t[72] = t[90] ^ x[41];
  assign t[73] = t[91] ^ x[42];
  assign t[74] = t[92] ^ x[51];
  assign t[75] = t[93] ^ x[52];
  assign t[76] = (t[94] & ~t[96] & ~t[97] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & ~t[97] & ~t[98] & ~t[100]) | (t[94] & ~t[95] & ~t[96] & ~t[99] & ~t[100]) | (~t[94] & t[95] & t[96] & t[97] & ~t[100]) | (~t[94] & t[95] & t[98] & t[99] & ~t[100]) | (t[94] & ~t[96] & ~t[98] & t[100]) | (~t[94] & t[96] & t[98] & t[100]);
  assign t[77] = (t[94] & t[95] & ~t[96] & ~t[98] & t[99] & ~t[100]) | (t[94] & t[96] & ~t[97] & ~t[98] & ~t[99] & t[100]) | (~t[95] & ~t[96] & t[98] & ~t[99] & ~t[100]) | (~t[94] & ~t[96] & ~t[97] & t[98] & ~t[99]) | (~t[94] & ~t[95] & ~t[97] & t[98] & ~t[100]) | (~t[94] & ~t[96] & t[97] & t[98] & t[99]) | (t[97] & t[98] & ~t[99] & ~t[100]);
  assign t[78] = (t[101] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & ~t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[102] & ~t[103] & ~t[106] & ~t[107]) | (~t[101] & t[102] & t[103] & t[104] & ~t[107]) | (~t[101] & t[102] & t[105] & t[106] & ~t[107]) | (t[101] & ~t[103] & ~t[105] & t[107]) | (~t[101] & t[103] & t[105] & t[107]);
  assign t[79] = (t[101] & t[102] & ~t[103] & t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[103] & ~t[104] & t[105] & ~t[106] & t[107]) | (~t[102] & t[103] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[102] & t[103] & ~t[106] & ~t[107]) | (~t[101] & t[103] & t[104] & ~t[105] & t[106]) | (t[103] & ~t[104] & t[106] & ~t[107]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[81] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[82] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[83] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[84] = (t[102] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & t[102] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[102] & ~t[103] & ~t[106] & ~t[107]) | (t[101] & ~t[102] & t[103] & t[104] & ~t[107]) | (t[101] & ~t[102] & t[105] & t[106] & ~t[107]) | (t[102] & ~t[104] & ~t[106] & t[107]) | (~t[102] & t[104] & t[106] & t[107]);
  assign t[85] = (t[101] & t[102] & t[103] & ~t[104] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & ~t[104] & ~t[105] & t[106] & t[107]) | (~t[102] & ~t[103] & t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[103] & t[104] & ~t[106] & ~t[107]) | (~t[101] & ~t[102] & t[104] & ~t[105] & ~t[107]) | (~t[102] & t[103] & t[104] & t[105] & ~t[106]) | (~t[103] & t[104] & t[105] & ~t[107]);
  assign t[86] = (t[101] & t[102] & ~t[103] & ~t[105] & t[106] & ~t[107]) | (t[101] & t[103] & ~t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & t[105] & ~t[106] & ~t[107]) | (~t[101] & ~t[103] & ~t[104] & t[105] & ~t[106]) | (~t[101] & ~t[102] & ~t[104] & t[105] & ~t[107]) | (~t[101] & ~t[103] & t[104] & t[105] & t[106]) | (t[104] & t[105] & ~t[106] & ~t[107]);
  assign t[87] = (t[101] & t[102] & ~t[104] & t[105] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[104] & ~t[105] & t[106] & ~t[107]) | (~t[101] & ~t[102] & ~t[103] & t[106] & ~t[107]) | (~t[102] & t[103] & ~t[104] & t[105] & t[106]) | (t[103] & ~t[105] & t[106] & ~t[107]);
  assign t[88] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[89] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[8] = ~(t[11]);
  assign t[90] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[91] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[93] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[94] = t[129] ^ x[9];
  assign t[95] = t[130] ^ x[4];
  assign t[96] = t[131] ^ x[5];
  assign t[97] = t[132] ^ x[6];
  assign t[98] = t[133] ^ x[10];
  assign t[99] = t[134] ^ x[7];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind157(x, y);
 input [54:0] x;
 output y;

 wire [159:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[36];
  assign t[101] = t[136] ^ x[37];
  assign t[102] = t[137] ^ x[38];
  assign t[103] = t[138] ^ x[17];
  assign t[104] = t[139] ^ x[26];
  assign t[105] = t[140] ^ x[21];
  assign t[106] = t[141] ^ x[22];
  assign t[107] = t[142] ^ x[23];
  assign t[108] = t[143] ^ x[27];
  assign t[109] = t[144] ^ x[24];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[145] ^ x[25];
  assign t[111] = t[146] ^ x[33];
  assign t[112] = t[147] ^ x[39];
  assign t[113] = t[148] ^ x[34];
  assign t[114] = t[149] ^ x[40];
  assign t[115] = t[150] ^ x[41];
  assign t[116] = t[151] ^ x[42];
  assign t[117] = t[152] ^ x[32];
  assign t[118] = t[153] ^ x[51];
  assign t[119] = t[154] ^ x[46];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[47];
  assign t[121] = t[156] ^ x[48];
  assign t[122] = t[157] ^ x[52];
  assign t[123] = t[158] ^ x[49];
  assign t[124] = t[159] ^ x[50];
  assign t[125] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[126] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[127] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[128] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[133] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[134] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[135] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[136] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[137] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[138] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[139] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[141] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[142] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[147] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[148] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[149] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[14] = ~(t[44] | t[20]);
  assign t[150] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[151] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[152] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[153] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[154] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[155] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[156] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[157] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[158] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[45];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[46] | t[23]);
  assign t[18] = ~(t[47]);
  assign t[19] = ~(t[48]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[49]);
  assign t[22] = ~(t[50]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[51]);
  assign t[25] = ~(t[47] | t[48]);
  assign t[26] = ~(t[52]);
  assign t[27] = ~(t[49] | t[50]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[53];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[19] & t[24]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[13] | t[44];
  assign t[41] = ~(t[22] & t[26]);
  assign t[42] = t[16] | t[46];
  assign t[43] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[44] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[45] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[46] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[47] = (t[56] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[56] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[48] = (t[56] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[56] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[49] = (t[60] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[60] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[60] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[60] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[51] = (t[56] & ~t[64]) | (~t[56] & t[64]);
  assign t[52] = (t[60] & ~t[68]) | (~t[60] & t[68]);
  assign t[53] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[18];
  assign t[57] = t[75] ^ x[19];
  assign t[58] = t[76] ^ x[26];
  assign t[59] = t[77] ^ x[27];
  assign t[5] = ~(~x[2] & ~t[43]);
  assign t[60] = t[78] ^ x[33];
  assign t[61] = t[79] ^ x[34];
  assign t[62] = t[80] ^ x[35];
  assign t[63] = t[81] ^ x[36];
  assign t[64] = t[82] ^ x[37];
  assign t[65] = t[83] ^ x[38];
  assign t[66] = t[84] ^ x[39];
  assign t[67] = t[85] ^ x[40];
  assign t[68] = t[86] ^ x[41];
  assign t[69] = t[87] ^ x[42];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[51];
  assign t[71] = t[89] ^ x[52];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[76] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[77] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[78] = (t[111] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (t[111] & ~t[112] & ~t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[112] & ~t[113] & ~t[116] & ~t[117]) | (~t[111] & t[112] & t[113] & t[114] & ~t[117]) | (~t[111] & t[112] & t[115] & t[116] & ~t[117]) | (t[111] & ~t[113] & ~t[115] & t[117]) | (~t[111] & t[113] & t[115] & t[117]);
  assign t[79] = (t[111] & t[112] & ~t[113] & t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[113] & ~t[114] & t[115] & ~t[116] & t[117]) | (~t[112] & t[113] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[112] & t[113] & ~t[116] & ~t[117]) | (~t[111] & t[113] & t[114] & ~t[115] & t[116]) | (t[113] & ~t[114] & t[116] & ~t[117]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[81] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[82] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[83] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[84] = (t[112] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & t[112] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[112] & ~t[113] & ~t[116] & ~t[117]) | (t[111] & ~t[112] & t[113] & t[114] & ~t[117]) | (t[111] & ~t[112] & t[115] & t[116] & ~t[117]) | (t[112] & ~t[114] & ~t[116] & t[117]) | (~t[112] & t[114] & t[116] & t[117]);
  assign t[85] = (t[111] & t[112] & t[113] & ~t[114] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[114] & ~t[115] & t[116] & t[117]) | (~t[112] & ~t[113] & t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[113] & t[114] & ~t[116] & ~t[117]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[117]) | (~t[112] & t[113] & t[114] & t[115] & ~t[116]) | (~t[113] & t[114] & t[115] & ~t[117]);
  assign t[86] = (t[111] & t[112] & ~t[113] & ~t[115] & t[116] & ~t[117]) | (t[111] & t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[117]) | (~t[111] & ~t[113] & ~t[114] & t[115] & ~t[116]) | (~t[111] & ~t[112] & ~t[114] & t[115] & ~t[117]) | (~t[111] & ~t[113] & t[114] & t[115] & t[116]) | (t[114] & t[115] & ~t[116] & ~t[117]);
  assign t[87] = (t[111] & t[112] & ~t[114] & t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[111] & ~t[112] & ~t[113] & t[116] & ~t[117]) | (~t[112] & t[113] & ~t[114] & t[115] & t[116]) | (t[113] & ~t[115] & t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[120] & ~t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[121] & ~t[122] & ~t[124]) | (t[118] & ~t[119] & ~t[120] & ~t[123] & ~t[124]) | (~t[118] & t[119] & t[120] & t[121] & ~t[124]) | (~t[118] & t[119] & t[122] & t[123] & ~t[124]) | (t[118] & ~t[120] & ~t[122] & t[124]) | (~t[118] & t[120] & t[122] & t[124]);
  assign t[89] = (t[118] & t[119] & ~t[120] & ~t[122] & t[123] & ~t[124]) | (t[118] & t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[124]) | (~t[118] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[118] & ~t[119] & ~t[121] & t[122] & ~t[124]) | (~t[118] & ~t[120] & t[121] & t[122] & t[123]) | (t[121] & t[122] & ~t[123] & ~t[124]);
  assign t[8] = ~(t[11]);
  assign t[90] = t[125] ^ x[9];
  assign t[91] = t[126] ^ x[4];
  assign t[92] = t[127] ^ x[5];
  assign t[93] = t[128] ^ x[6];
  assign t[94] = t[129] ^ x[10];
  assign t[95] = t[130] ^ x[7];
  assign t[96] = t[131] ^ x[8];
  assign t[97] = t[132] ^ x[18];
  assign t[98] = t[133] ^ x[35];
  assign t[99] = t[134] ^ x[19];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind158(x, y);
 input [54:0] x;
 output y;

 wire [161:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[19];
  assign t[101] = t[136] ^ x[53];
  assign t[102] = t[137] ^ x[20];
  assign t[103] = t[138] ^ x[21];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[17];
  assign t[106] = t[141] ^ x[29];
  assign t[107] = t[142] ^ x[24];
  assign t[108] = t[143] ^ x[25];
  assign t[109] = t[144] ^ x[26];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[145] ^ x[30];
  assign t[111] = t[146] ^ x[27];
  assign t[112] = t[147] ^ x[28];
  assign t[113] = t[148] ^ x[36];
  assign t[114] = t[149] ^ x[37];
  assign t[115] = t[150] ^ x[54];
  assign t[116] = t[151] ^ x[38];
  assign t[117] = t[152] ^ x[39];
  assign t[118] = t[153] ^ x[40];
  assign t[119] = t[154] ^ x[35];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[49];
  assign t[121] = t[156] ^ x[44];
  assign t[122] = t[157] ^ x[45];
  assign t[123] = t[158] ^ x[46];
  assign t[124] = t[159] ^ x[50];
  assign t[125] = t[160] ^ x[47];
  assign t[126] = t[161] ^ x[48];
  assign t[127] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[128] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[129] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[12] = ~(t[16] & t[17]);
  assign t[130] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[133] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[134] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[135] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[136] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[137] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[138] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[139] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[13] = ~(t[46] & t[18]);
  assign t[140] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[141] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[142] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[143] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[144] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[31] & ~x[32] & ~x[33]) | (~x[31] & x[32] & ~x[33]) | (~x[31] & ~x[32] & x[33]) | (x[31] & x[32] & x[33]);
  assign t[149] = (x[31] & ~x[32] & ~x[34]) | (~x[31] & x[32] & ~x[34]) | (~x[31] & ~x[32] & x[34]) | (x[31] & x[32] & x[34]);
  assign t[14] = ~(t[47] & t[19]);
  assign t[150] = (x[31] & ~x[33]) | (~x[31] & x[33]);
  assign t[151] = (x[31] & ~x[34]) | (~x[31] & x[34]);
  assign t[152] = (x[32] & ~x[33]) | (~x[32] & x[33]);
  assign t[153] = (x[32] & ~x[34]) | (~x[32] & x[34]);
  assign t[154] = (x[33] & ~x[34]) | (~x[33] & x[34]);
  assign t[155] = (x[43] & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0);
  assign t[156] = (x[43] & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0);
  assign t[157] = (x[43] & ~1'b0) | (~x[43] & 1'b0);
  assign t[158] = (x[43] & ~1'b0) | (~x[43] & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[48];
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[16] = ~(t[49] & t[20]);
  assign t[17] = ~(t[50] & t[21]);
  assign t[18] = ~(t[51]);
  assign t[19] = ~(t[51] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[52]);
  assign t[21] = ~(t[52] & t[23]);
  assign t[22] = ~(t[46]);
  assign t[23] = ~(t[49]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27];
  assign t[26] = ~(t[28] ^ t[29]);
  assign t[27] = ~(t[30] ^ t[31]);
  assign t[28] = t[8] ? x[42] : x[41];
  assign t[29] = ~x[2] & t[53];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[51] : t[33];
  assign t[32] = x[2] ? x[52] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[18] & t[39]);
  assign t[36] = ~(t[40] & t[54]);
  assign t[37] = ~(t[20] & t[41]);
  assign t[38] = ~(t[42] & t[55]);
  assign t[39] = ~(t[47]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[43] & t[22]);
  assign t[41] = ~(t[50]);
  assign t[42] = ~(t[44] & t[23]);
  assign t[43] = ~(t[47] & t[51]);
  assign t[44] = ~(t[50] & t[52]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[58] & ~t[60] & ~t[62]) | (~t[59] & t[60] & ~t[61]) | (~t[58] & ~t[60] & t[62]) | (t[59] & t[60] & t[61]);
  assign t[47] = (t[58] & ~t[61]) | (~t[58] & t[61]);
  assign t[48] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[49] = (t[65] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[65] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[65] & ~t[68]) | (~t[65] & t[68]);
  assign t[51] = (t[58] & ~t[60] & ~t[61]) | (~t[59] & t[60] & ~t[62]) | (~t[58] & ~t[60] & t[61]) | (t[59] & t[60] & t[62]);
  assign t[52] = (t[65] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[65] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[53] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[54] = (t[58] & ~t[72]) | (~t[58] & t[72]);
  assign t[55] = (t[65] & ~t[73]) | (~t[65] & t[73]);
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[10];
  assign t[58] = t[76] ^ x[18];
  assign t[59] = t[77] ^ x[19];
  assign t[5] = ~x[2] & t[45];
  assign t[60] = t[78] ^ x[20];
  assign t[61] = t[79] ^ x[21];
  assign t[62] = t[80] ^ x[22];
  assign t[63] = t[81] ^ x[29];
  assign t[64] = t[82] ^ x[30];
  assign t[65] = t[83] ^ x[36];
  assign t[66] = t[84] ^ x[37];
  assign t[67] = t[85] ^ x[38];
  assign t[68] = t[86] ^ x[39];
  assign t[69] = t[87] ^ x[40];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[49];
  assign t[71] = t[89] ^ x[50];
  assign t[72] = t[90] ^ x[53];
  assign t[73] = t[91] ^ x[54];
  assign t[74] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[78] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[79] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[82] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[83] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[84] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[85] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[86] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[87] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[89] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[8] = ~(t[11]);
  assign t[90] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = t[127] ^ x[9];
  assign t[93] = t[128] ^ x[4];
  assign t[94] = t[129] ^ x[5];
  assign t[95] = t[130] ^ x[6];
  assign t[96] = t[131] ^ x[10];
  assign t[97] = t[132] ^ x[7];
  assign t[98] = t[133] ^ x[8];
  assign t[99] = t[134] ^ x[18];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[24]) | (~t[0] & t[24]);
endmodule

module R2ind159(x, y);
 input [54:0] x;
 output y;

 wire [159:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[20];
  assign t[101] = t[136] ^ x[21];
  assign t[102] = t[137] ^ x[22];
  assign t[103] = t[138] ^ x[17];
  assign t[104] = t[139] ^ x[29];
  assign t[105] = t[140] ^ x[24];
  assign t[106] = t[141] ^ x[25];
  assign t[107] = t[142] ^ x[26];
  assign t[108] = t[143] ^ x[30];
  assign t[109] = t[144] ^ x[27];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[145] ^ x[28];
  assign t[111] = t[146] ^ x[36];
  assign t[112] = t[147] ^ x[37];
  assign t[113] = t[148] ^ x[54];
  assign t[114] = t[149] ^ x[38];
  assign t[115] = t[150] ^ x[39];
  assign t[116] = t[151] ^ x[40];
  assign t[117] = t[152] ^ x[35];
  assign t[118] = t[153] ^ x[49];
  assign t[119] = t[154] ^ x[44];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[45];
  assign t[121] = t[156] ^ x[46];
  assign t[122] = t[157] ^ x[50];
  assign t[123] = t[158] ^ x[47];
  assign t[124] = t[159] ^ x[48];
  assign t[125] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[126] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[127] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[128] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~(t[16] & t[17]);
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[133] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[134] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[135] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[136] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[137] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[138] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[139] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[13] = ~(t[44] & t[18]);
  assign t[140] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[141] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[142] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (x[31] & ~x[32] & ~x[33]) | (~x[31] & x[32] & ~x[33]) | (~x[31] & ~x[32] & x[33]) | (x[31] & x[32] & x[33]);
  assign t[147] = (x[31] & ~x[32] & ~x[34]) | (~x[31] & x[32] & ~x[34]) | (~x[31] & ~x[32] & x[34]) | (x[31] & x[32] & x[34]);
  assign t[148] = (x[31] & ~x[33]) | (~x[31] & x[33]);
  assign t[149] = (x[31] & ~x[34]) | (~x[31] & x[34]);
  assign t[14] = ~(t[45] & t[19]);
  assign t[150] = (x[32] & ~x[33]) | (~x[32] & x[33]);
  assign t[151] = (x[32] & ~x[34]) | (~x[32] & x[34]);
  assign t[152] = (x[33] & ~x[34]) | (~x[33] & x[34]);
  assign t[153] = (x[43] & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0);
  assign t[154] = (x[43] & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0);
  assign t[155] = (x[43] & ~1'b0) | (~x[43] & 1'b0);
  assign t[156] = (x[43] & ~1'b0) | (~x[43] & 1'b0);
  assign t[157] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[158] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[46];
  assign t[16] = ~(t[47] & t[20]);
  assign t[17] = ~(t[48] & t[21]);
  assign t[18] = ~(t[49]);
  assign t[19] = ~(t[49] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[50]);
  assign t[21] = ~(t[50] & t[23]);
  assign t[22] = ~(t[44]);
  assign t[23] = ~(t[47]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27];
  assign t[26] = ~(t[28] ^ t[29]);
  assign t[27] = ~(t[30] ^ t[31]);
  assign t[28] = t[8] ? x[42] : x[41];
  assign t[29] = ~x[2] & t[51];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[51] : t[33];
  assign t[32] = x[2] ? x[52] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[18] & t[39]);
  assign t[36] = t[40] | t[52];
  assign t[37] = ~(t[20] & t[41]);
  assign t[38] = t[42] | t[53];
  assign t[39] = ~(t[45]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[22] | t[18]);
  assign t[41] = ~(t[48]);
  assign t[42] = ~(t[23] | t[20]);
  assign t[43] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[44] = (t[56] & ~t[58] & ~t[60]) | (~t[57] & t[58] & ~t[59]) | (~t[56] & ~t[58] & t[60]) | (t[57] & t[58] & t[59]);
  assign t[45] = (t[56] & ~t[59]) | (~t[56] & t[59]);
  assign t[46] = (t[61] & ~t[62]) | (~t[61] & t[62]);
  assign t[47] = (t[63] & ~t[65] & ~t[67]) | (~t[64] & t[65] & ~t[66]) | (~t[63] & ~t[65] & t[67]) | (t[64] & t[65] & t[66]);
  assign t[48] = (t[63] & ~t[66]) | (~t[63] & t[66]);
  assign t[49] = (t[56] & ~t[58] & ~t[59]) | (~t[57] & t[58] & ~t[60]) | (~t[56] & ~t[58] & t[59]) | (t[57] & t[58] & t[60]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[63] & ~t[65] & ~t[66]) | (~t[64] & t[65] & ~t[67]) | (~t[63] & ~t[65] & t[66]) | (t[64] & t[65] & t[67]);
  assign t[51] = (t[68] & ~t[69]) | (~t[68] & t[69]);
  assign t[52] = (t[56] & ~t[70]) | (~t[56] & t[70]);
  assign t[53] = (t[63] & ~t[71]) | (~t[63] & t[71]);
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[18];
  assign t[57] = t[75] ^ x[19];
  assign t[58] = t[76] ^ x[20];
  assign t[59] = t[77] ^ x[21];
  assign t[5] = ~x[2] & t[43];
  assign t[60] = t[78] ^ x[22];
  assign t[61] = t[79] ^ x[29];
  assign t[62] = t[80] ^ x[30];
  assign t[63] = t[81] ^ x[36];
  assign t[64] = t[82] ^ x[37];
  assign t[65] = t[83] ^ x[38];
  assign t[66] = t[84] ^ x[39];
  assign t[67] = t[85] ^ x[40];
  assign t[68] = t[86] ^ x[49];
  assign t[69] = t[87] ^ x[50];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[53];
  assign t[71] = t[89] ^ x[54];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[76] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[77] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[78] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[79] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[81] = (t[111] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (t[111] & ~t[112] & ~t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[112] & ~t[113] & ~t[116] & ~t[117]) | (~t[111] & t[112] & t[113] & t[114] & ~t[117]) | (~t[111] & t[112] & t[115] & t[116] & ~t[117]) | (t[111] & ~t[113] & ~t[115] & t[117]) | (~t[111] & t[113] & t[115] & t[117]);
  assign t[82] = (t[112] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & t[112] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[112] & ~t[113] & ~t[116] & ~t[117]) | (t[111] & ~t[112] & t[113] & t[114] & ~t[117]) | (t[111] & ~t[112] & t[115] & t[116] & ~t[117]) | (t[112] & ~t[114] & ~t[116] & t[117]) | (~t[112] & t[114] & t[116] & t[117]);
  assign t[83] = (t[111] & t[112] & t[113] & ~t[114] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[114] & ~t[115] & t[116] & t[117]) | (~t[112] & ~t[113] & t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[113] & t[114] & ~t[116] & ~t[117]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[117]) | (~t[112] & t[113] & t[114] & t[115] & ~t[116]) | (~t[113] & t[114] & t[115] & ~t[117]);
  assign t[84] = (t[111] & t[112] & ~t[113] & ~t[115] & t[116] & ~t[117]) | (t[111] & t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[117]) | (~t[111] & ~t[113] & ~t[114] & t[115] & ~t[116]) | (~t[111] & ~t[112] & ~t[114] & t[115] & ~t[117]) | (~t[111] & ~t[113] & t[114] & t[115] & t[116]) | (t[114] & t[115] & ~t[116] & ~t[117]);
  assign t[85] = (t[111] & t[112] & ~t[114] & t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[111] & ~t[112] & ~t[113] & t[116] & ~t[117]) | (~t[112] & t[113] & ~t[114] & t[115] & t[116]) | (t[113] & ~t[115] & t[116] & ~t[117]);
  assign t[86] = (t[118] & ~t[120] & ~t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[121] & ~t[122] & ~t[124]) | (t[118] & ~t[119] & ~t[120] & ~t[123] & ~t[124]) | (~t[118] & t[119] & t[120] & t[121] & ~t[124]) | (~t[118] & t[119] & t[122] & t[123] & ~t[124]) | (t[118] & ~t[120] & ~t[122] & t[124]) | (~t[118] & t[120] & t[122] & t[124]);
  assign t[87] = (t[118] & t[119] & ~t[120] & ~t[122] & t[123] & ~t[124]) | (t[118] & t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[124]) | (~t[118] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[118] & ~t[119] & ~t[121] & t[122] & ~t[124]) | (~t[118] & ~t[120] & t[121] & t[122] & t[123]) | (t[121] & t[122] & ~t[123] & ~t[124]);
  assign t[88] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[89] = (t[111] & t[112] & ~t[113] & t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[113] & ~t[114] & t[115] & ~t[116] & t[117]) | (~t[112] & t[113] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[112] & t[113] & ~t[116] & ~t[117]) | (~t[111] & t[113] & t[114] & ~t[115] & t[116]) | (t[113] & ~t[114] & t[116] & ~t[117]);
  assign t[8] = ~(t[11]);
  assign t[90] = t[125] ^ x[9];
  assign t[91] = t[126] ^ x[4];
  assign t[92] = t[127] ^ x[5];
  assign t[93] = t[128] ^ x[6];
  assign t[94] = t[129] ^ x[10];
  assign t[95] = t[130] ^ x[7];
  assign t[96] = t[131] ^ x[8];
  assign t[97] = t[132] ^ x[18];
  assign t[98] = t[133] ^ x[19];
  assign t[99] = t[134] ^ x[53];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[24]) | (~t[0] & t[24]);
endmodule

module R2ind160(x, y);
 input [54:0] x;
 output y;

 wire [159:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[135] ^ x[36];
  assign t[101] = t[136] ^ x[37];
  assign t[102] = t[137] ^ x[38];
  assign t[103] = t[138] ^ x[17];
  assign t[104] = t[139] ^ x[26];
  assign t[105] = t[140] ^ x[21];
  assign t[106] = t[141] ^ x[22];
  assign t[107] = t[142] ^ x[23];
  assign t[108] = t[143] ^ x[27];
  assign t[109] = t[144] ^ x[24];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[145] ^ x[25];
  assign t[111] = t[146] ^ x[33];
  assign t[112] = t[147] ^ x[39];
  assign t[113] = t[148] ^ x[34];
  assign t[114] = t[149] ^ x[40];
  assign t[115] = t[150] ^ x[41];
  assign t[116] = t[151] ^ x[42];
  assign t[117] = t[152] ^ x[32];
  assign t[118] = t[153] ^ x[51];
  assign t[119] = t[154] ^ x[46];
  assign t[11] = ~(t[15]);
  assign t[120] = t[155] ^ x[47];
  assign t[121] = t[156] ^ x[48];
  assign t[122] = t[157] ^ x[52];
  assign t[123] = t[158] ^ x[49];
  assign t[124] = t[159] ^ x[50];
  assign t[125] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[126] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[127] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[128] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = ~(t[16] & t[17]);
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[133] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[134] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[135] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[136] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[137] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[138] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[139] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[13] = ~(t[18] & t[19]);
  assign t[140] = (x[20] & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0);
  assign t[141] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[142] = (x[20] & ~1'b0) | (~x[20] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[147] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[148] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[149] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[14] = ~(t[20] & t[44]);
  assign t[150] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[151] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[152] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[153] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[154] = (x[45] & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0);
  assign t[155] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[156] = (x[45] & ~1'b0) | (~x[45] & 1'b0);
  assign t[157] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[158] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~x[2] & t[45];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[46]);
  assign t[18] = ~(t[47]);
  assign t[19] = ~(t[48]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[49]);
  assign t[22] = ~(t[50]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[48] & t[47]);
  assign t[25] = ~(t[51]);
  assign t[26] = ~(t[50] & t[49]);
  assign t[27] = ~(t[52]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[44] : x[43];
  assign t[33] = ~x[2] & t[53];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[53] : t[37];
  assign t[36] = x[2] ? x[54] : t[38];
  assign t[37] = ~(t[13] & t[39]);
  assign t[38] = ~(t[16] & t[40]);
  assign t[39] = t[41] | t[44];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[42] | t[46];
  assign t[41] = ~(t[25] | t[18]);
  assign t[42] = ~(t[27] | t[21]);
  assign t[43] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[44] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[45] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[46] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[47] = (t[56] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[56] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[48] = (t[56] & ~t[64]) | (~t[56] & t[64]);
  assign t[49] = (t[60] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[60] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[60] & ~t[68]) | (~t[60] & t[68]);
  assign t[51] = (t[56] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[56] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[52] = (t[60] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[60] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[18];
  assign t[57] = t[75] ^ x[19];
  assign t[58] = t[76] ^ x[26];
  assign t[59] = t[77] ^ x[27];
  assign t[5] = ~x[2] & t[43];
  assign t[60] = t[78] ^ x[33];
  assign t[61] = t[79] ^ x[34];
  assign t[62] = t[80] ^ x[35];
  assign t[63] = t[81] ^ x[36];
  assign t[64] = t[82] ^ x[37];
  assign t[65] = t[83] ^ x[38];
  assign t[66] = t[84] ^ x[39];
  assign t[67] = t[85] ^ x[40];
  assign t[68] = t[86] ^ x[41];
  assign t[69] = t[87] ^ x[42];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[51];
  assign t[71] = t[89] ^ x[52];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[76] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[77] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[78] = (t[111] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (t[111] & ~t[112] & ~t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[112] & ~t[113] & ~t[116] & ~t[117]) | (~t[111] & t[112] & t[113] & t[114] & ~t[117]) | (~t[111] & t[112] & t[115] & t[116] & ~t[117]) | (t[111] & ~t[113] & ~t[115] & t[117]) | (~t[111] & t[113] & t[115] & t[117]);
  assign t[79] = (t[111] & t[112] & ~t[113] & t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[113] & ~t[114] & t[115] & ~t[116] & t[117]) | (~t[112] & t[113] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[112] & t[113] & ~t[116] & ~t[117]) | (~t[111] & t[113] & t[114] & ~t[115] & t[116]) | (t[113] & ~t[114] & t[116] & ~t[117]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[81] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[82] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[83] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[84] = (t[112] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & t[112] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[112] & ~t[113] & ~t[116] & ~t[117]) | (t[111] & ~t[112] & t[113] & t[114] & ~t[117]) | (t[111] & ~t[112] & t[115] & t[116] & ~t[117]) | (t[112] & ~t[114] & ~t[116] & t[117]) | (~t[112] & t[114] & t[116] & t[117]);
  assign t[85] = (t[111] & t[112] & t[113] & ~t[114] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[114] & ~t[115] & t[116] & t[117]) | (~t[112] & ~t[113] & t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[113] & t[114] & ~t[116] & ~t[117]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[117]) | (~t[112] & t[113] & t[114] & t[115] & ~t[116]) | (~t[113] & t[114] & t[115] & ~t[117]);
  assign t[86] = (t[111] & t[112] & ~t[113] & ~t[115] & t[116] & ~t[117]) | (t[111] & t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[117]) | (~t[111] & ~t[113] & ~t[114] & t[115] & ~t[116]) | (~t[111] & ~t[112] & ~t[114] & t[115] & ~t[117]) | (~t[111] & ~t[113] & t[114] & t[115] & t[116]) | (t[114] & t[115] & ~t[116] & ~t[117]);
  assign t[87] = (t[111] & t[112] & ~t[114] & t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[111] & ~t[112] & ~t[113] & t[116] & ~t[117]) | (~t[112] & t[113] & ~t[114] & t[115] & t[116]) | (t[113] & ~t[115] & t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[120] & ~t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[121] & ~t[122] & ~t[124]) | (t[118] & ~t[119] & ~t[120] & ~t[123] & ~t[124]) | (~t[118] & t[119] & t[120] & t[121] & ~t[124]) | (~t[118] & t[119] & t[122] & t[123] & ~t[124]) | (t[118] & ~t[120] & ~t[122] & t[124]) | (~t[118] & t[120] & t[122] & t[124]);
  assign t[89] = (t[118] & t[119] & ~t[120] & ~t[122] & t[123] & ~t[124]) | (t[118] & t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[124]) | (~t[118] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[118] & ~t[119] & ~t[121] & t[122] & ~t[124]) | (~t[118] & ~t[120] & t[121] & t[122] & t[123]) | (t[121] & t[122] & ~t[123] & ~t[124]);
  assign t[8] = ~(t[11]);
  assign t[90] = t[125] ^ x[9];
  assign t[91] = t[126] ^ x[4];
  assign t[92] = t[127] ^ x[5];
  assign t[93] = t[128] ^ x[6];
  assign t[94] = t[129] ^ x[10];
  assign t[95] = t[130] ^ x[7];
  assign t[96] = t[131] ^ x[8];
  assign t[97] = t[132] ^ x[18];
  assign t[98] = t[133] ^ x[35];
  assign t[99] = t[134] ^ x[19];
  assign t[9] = x[2] ? x[12] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind161(x, y);
 input [56:0] x;
 output y;

 wire [189:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[33];
  assign t[101] = t[121] ^ x[34];
  assign t[102] = t[122] ^ x[35];
  assign t[103] = t[123] ^ x[36];
  assign t[104] = t[124] ^ x[37];
  assign t[105] = t[125] ^ x[38];
  assign t[106] = t[126] ^ x[39];
  assign t[107] = t[127] ^ x[40];
  assign t[108] = t[128] ^ x[41];
  assign t[109] = t[129] ^ x[42];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[130] ^ x[43];
  assign t[111] = t[131] ^ x[44];
  assign t[112] = t[132] ^ x[45];
  assign t[113] = t[133] ^ x[46];
  assign t[114] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[115] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[116] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[117] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[118] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[119] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[11] = ~x[2] & t[81];
  assign t[120] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[121] = (t[155] & t[156] & ~t[157] & t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[157] & ~t[158] & t[159] & ~t[160] & t[161]) | (~t[156] & t[157] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[156] & t[157] & ~t[160] & ~t[161]) | (~t[155] & t[157] & t[158] & ~t[159] & t[160]) | (t[157] & ~t[158] & t[160] & ~t[161]);
  assign t[122] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[123] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[124] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[125] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[126] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[127] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[128] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[129] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (t[156] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & t[156] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[156] & ~t[157] & ~t[160] & ~t[161]) | (t[155] & ~t[156] & t[157] & t[158] & ~t[161]) | (t[155] & ~t[156] & t[159] & t[160] & ~t[161]) | (t[156] & ~t[158] & ~t[160] & t[161]) | (~t[156] & t[158] & t[160] & t[161]);
  assign t[131] = (t[155] & t[156] & t[157] & ~t[158] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & ~t[158] & ~t[159] & t[160] & t[161]) | (~t[156] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[157] & t[158] & ~t[160] & ~t[161]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[161]) | (~t[156] & t[157] & t[158] & t[159] & ~t[160]) | (~t[157] & t[158] & t[159] & ~t[161]);
  assign t[132] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[133] = (t[155] & t[156] & ~t[158] & t[159] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[158] & ~t[159] & t[160] & ~t[161]) | (~t[155] & ~t[156] & ~t[157] & t[160] & ~t[161]) | (~t[156] & t[157] & ~t[158] & t[159] & t[160]) | (t[157] & ~t[159] & t[160] & ~t[161]);
  assign t[134] = t[162] ^ x[12];
  assign t[135] = t[163] ^ x[7];
  assign t[136] = t[164] ^ x[8];
  assign t[137] = t[165] ^ x[9];
  assign t[138] = t[166] ^ x[13];
  assign t[139] = t[167] ^ x[10];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[11];
  assign t[141] = t[169] ^ x[19];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[20];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[18];
  assign t[148] = t[176] ^ x[26];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[178] ^ x[27];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[25];
  assign t[155] = t[183] ^ x[33];
  assign t[156] = t[184] ^ x[43];
  assign t[157] = t[185] ^ x[34];
  assign t[158] = t[186] ^ x[44];
  assign t[159] = t[187] ^ x[45];
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = t[188] ^ x[46];
  assign t[161] = t[189] ^ x[32];
  assign t[162] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[163] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[164] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[165] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[166] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[167] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[168] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[169] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[16] = ~(t[82] | t[23]);
  assign t[170] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[171] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[172] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[173] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[174] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[175] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[176] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[177] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[178] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[179] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[180] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[181] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[182] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[183] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[184] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[185] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[186] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[187] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[188] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[189] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[83] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[84] | t[29]);
  assign t[21] = ~(t[85]);
  assign t[22] = ~(t[86]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[87]);
  assign t[25] = ~(t[88]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[89]);
  assign t[28] = ~(t[90]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[91]);
  assign t[31] = ~(t[85] | t[86]);
  assign t[32] = ~(t[92]);
  assign t[33] = ~(t[87] | t[88]);
  assign t[34] = ~(t[93]);
  assign t[35] = ~(t[89] | t[90]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[85] & t[22]);
  assign t[49] = ~(t[91] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[87] & t[25]);
  assign t[51] = ~(t[92] & t[55]);
  assign t[52] = ~(t[89] & t[28]);
  assign t[53] = ~(t[93] & t[56]);
  assign t[54] = ~(t[86] & t[21]);
  assign t[55] = ~(t[88] & t[24]);
  assign t[56] = ~(t[90] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[4] ? x[53] : x[52];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = ~(t[75] & t[82]);
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = ~(t[76] & t[83]);
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = ~(t[77] & t[84]);
  assign t[75] = ~(t[78] & t[21]);
  assign t[76] = ~(t[79] & t[24]);
  assign t[77] = ~(t[80] & t[27]);
  assign t[78] = ~(t[91] & t[86]);
  assign t[79] = ~(t[92] & t[88]);
  assign t[7] = ~(t[11]);
  assign t[80] = ~(t[93] & t[90]);
  assign t[81] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[82] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[83] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[84] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[85] = (t[96] & ~t[103] & ~t[105]) | (~t[102] & t[103] & ~t[104]) | (~t[96] & ~t[103] & t[105]) | (t[102] & t[103] & t[104]);
  assign t[86] = (t[96] & ~t[103] & ~t[104]) | (~t[102] & t[103] & ~t[105]) | (~t[96] & ~t[103] & t[104]) | (t[102] & t[103] & t[105]);
  assign t[87] = (t[98] & ~t[107] & ~t[109]) | (~t[106] & t[107] & ~t[108]) | (~t[98] & ~t[107] & t[109]) | (t[106] & t[107] & t[108]);
  assign t[88] = (t[98] & ~t[107] & ~t[108]) | (~t[106] & t[107] & ~t[109]) | (~t[98] & ~t[107] & t[108]) | (t[106] & t[107] & t[109]);
  assign t[89] = (t[100] & ~t[111] & ~t[113]) | (~t[110] & t[111] & ~t[112]) | (~t[100] & ~t[111] & t[113]) | (t[110] & t[111] & t[112]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[100] & ~t[111] & ~t[112]) | (~t[110] & t[111] & ~t[113]) | (~t[100] & ~t[111] & t[112]) | (t[110] & t[111] & t[113]);
  assign t[91] = (t[96] & ~t[104]) | (~t[96] & t[104]);
  assign t[92] = (t[98] & ~t[108]) | (~t[98] & t[108]);
  assign t[93] = (t[100] & ~t[112]) | (~t[100] & t[112]);
  assign t[94] = t[114] ^ x[12];
  assign t[95] = t[115] ^ x[13];
  assign t[96] = t[116] ^ x[19];
  assign t[97] = t[117] ^ x[20];
  assign t[98] = t[118] ^ x[26];
  assign t[99] = t[119] ^ x[27];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57]) | (~t[0] & t[36] & ~t[57]) | (~t[0] & ~t[36] & t[57]) | (t[0] & t[36] & t[57]);
endmodule

module R2ind162(x, y);
 input [56:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[39];
  assign t[101] = t[121] ^ x[40];
  assign t[102] = t[122] ^ x[41];
  assign t[103] = t[123] ^ x[42];
  assign t[104] = t[124] ^ x[43];
  assign t[105] = t[125] ^ x[44];
  assign t[106] = t[126] ^ x[45];
  assign t[107] = t[127] ^ x[46];
  assign t[108] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[109] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (t[135] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[136] & ~t[137] & ~t[140] & ~t[141]) | (~t[135] & t[136] & t[137] & t[138] & ~t[141]) | (~t[135] & t[136] & t[139] & t[140] & ~t[141]) | (t[135] & ~t[137] & ~t[139] & t[141]) | (~t[135] & t[137] & t[139] & t[141]);
  assign t[111] = (t[135] & t[136] & ~t[137] & t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[137] & ~t[138] & t[139] & ~t[140] & t[141]) | (~t[136] & t[137] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[136] & t[137] & ~t[140] & ~t[141]) | (~t[135] & t[137] & t[138] & ~t[139] & t[140]) | (t[137] & ~t[138] & t[140] & ~t[141]);
  assign t[112] = (t[142] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[143] & ~t[144] & ~t[147] & ~t[148]) | (~t[142] & t[143] & t[144] & t[145] & ~t[148]) | (~t[142] & t[143] & t[146] & t[147] & ~t[148]) | (t[142] & ~t[144] & ~t[146] & t[148]) | (~t[142] & t[144] & t[146] & t[148]);
  assign t[113] = (t[142] & t[143] & ~t[144] & t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[144] & ~t[145] & t[146] & ~t[147] & t[148]) | (~t[143] & t[144] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[143] & t[144] & ~t[147] & ~t[148]) | (~t[142] & t[144] & t[145] & ~t[146] & t[147]) | (t[144] & ~t[145] & t[147] & ~t[148]);
  assign t[114] = (t[149] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[150] & ~t[151] & ~t[154] & ~t[155]) | (~t[149] & t[150] & t[151] & t[152] & ~t[155]) | (~t[149] & t[150] & t[153] & t[154] & ~t[155]) | (t[149] & ~t[151] & ~t[153] & t[155]) | (~t[149] & t[151] & t[153] & t[155]);
  assign t[115] = (t[149] & t[150] & ~t[151] & t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[151] & ~t[152] & t[153] & ~t[154] & t[155]) | (~t[150] & t[151] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[150] & t[151] & ~t[154] & ~t[155]) | (~t[149] & t[151] & t[152] & ~t[153] & t[154]) | (t[151] & ~t[152] & t[154] & ~t[155]);
  assign t[116] = (t[136] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & t[136] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[136] & ~t[137] & ~t[140] & ~t[141]) | (t[135] & ~t[136] & t[137] & t[138] & ~t[141]) | (t[135] & ~t[136] & t[139] & t[140] & ~t[141]) | (t[136] & ~t[138] & ~t[140] & t[141]) | (~t[136] & t[138] & t[140] & t[141]);
  assign t[117] = (t[135] & t[136] & t[137] & ~t[138] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & ~t[138] & ~t[139] & t[140] & t[141]) | (~t[136] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[137] & t[138] & ~t[140] & ~t[141]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[141]) | (~t[136] & t[137] & t[138] & t[139] & ~t[140]) | (~t[137] & t[138] & t[139] & ~t[141]);
  assign t[118] = (t[135] & t[136] & ~t[137] & ~t[139] & t[140] & ~t[141]) | (t[135] & t[137] & ~t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & t[139] & ~t[140] & ~t[141]) | (~t[135] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[135] & ~t[136] & ~t[138] & t[139] & ~t[141]) | (~t[135] & ~t[137] & t[138] & t[139] & t[140]) | (t[138] & t[139] & ~t[140] & ~t[141]);
  assign t[119] = (t[135] & t[136] & ~t[138] & t[139] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[138] & ~t[139] & t[140] & ~t[141]) | (~t[135] & ~t[136] & ~t[137] & t[140] & ~t[141]) | (~t[136] & t[137] & ~t[138] & t[139] & t[140]) | (t[137] & ~t[139] & t[140] & ~t[141]);
  assign t[11] = ~x[2] & t[75];
  assign t[120] = (t[143] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & t[143] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[143] & ~t[144] & ~t[147] & ~t[148]) | (t[142] & ~t[143] & t[144] & t[145] & ~t[148]) | (t[142] & ~t[143] & t[146] & t[147] & ~t[148]) | (t[143] & ~t[145] & ~t[147] & t[148]) | (~t[143] & t[145] & t[147] & t[148]);
  assign t[121] = (t[142] & t[143] & t[144] & ~t[145] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & ~t[145] & ~t[146] & t[147] & t[148]) | (~t[143] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[144] & t[145] & ~t[147] & ~t[148]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[148]) | (~t[143] & t[144] & t[145] & t[146] & ~t[147]) | (~t[144] & t[145] & t[146] & ~t[148]);
  assign t[122] = (t[142] & t[143] & ~t[144] & ~t[146] & t[147] & ~t[148]) | (t[142] & t[144] & ~t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & t[146] & ~t[147] & ~t[148]) | (~t[142] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[142] & ~t[143] & ~t[145] & t[146] & ~t[148]) | (~t[142] & ~t[144] & t[145] & t[146] & t[147]) | (t[145] & t[146] & ~t[147] & ~t[148]);
  assign t[123] = (t[142] & t[143] & ~t[145] & t[146] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[145] & ~t[146] & t[147] & ~t[148]) | (~t[142] & ~t[143] & ~t[144] & t[147] & ~t[148]) | (~t[143] & t[144] & ~t[145] & t[146] & t[147]) | (t[144] & ~t[146] & t[147] & ~t[148]);
  assign t[124] = (t[150] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & t[150] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[150] & ~t[151] & ~t[154] & ~t[155]) | (t[149] & ~t[150] & t[151] & t[152] & ~t[155]) | (t[149] & ~t[150] & t[153] & t[154] & ~t[155]) | (t[150] & ~t[152] & ~t[154] & t[155]) | (~t[150] & t[152] & t[154] & t[155]);
  assign t[125] = (t[149] & t[150] & t[151] & ~t[152] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & ~t[152] & ~t[153] & t[154] & t[155]) | (~t[150] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[151] & t[152] & ~t[154] & ~t[155]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[155]) | (~t[150] & t[151] & t[152] & t[153] & ~t[154]) | (~t[151] & t[152] & t[153] & ~t[155]);
  assign t[126] = (t[149] & t[150] & ~t[151] & ~t[153] & t[154] & ~t[155]) | (t[149] & t[151] & ~t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & t[153] & ~t[154] & ~t[155]) | (~t[149] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[149] & ~t[150] & ~t[152] & t[153] & ~t[155]) | (~t[149] & ~t[151] & t[152] & t[153] & t[154]) | (t[152] & t[153] & ~t[154] & ~t[155]);
  assign t[127] = (t[149] & t[150] & ~t[152] & t[153] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[152] & ~t[153] & t[154] & ~t[155]) | (~t[149] & ~t[150] & ~t[151] & t[154] & ~t[155]) | (~t[150] & t[151] & ~t[152] & t[153] & t[154]) | (t[151] & ~t[153] & t[154] & ~t[155]);
  assign t[128] = t[156] ^ x[12];
  assign t[129] = t[157] ^ x[7];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[8];
  assign t[131] = t[159] ^ x[9];
  assign t[132] = t[160] ^ x[13];
  assign t[133] = t[161] ^ x[10];
  assign t[134] = t[162] ^ x[11];
  assign t[135] = t[163] ^ x[19];
  assign t[136] = t[164] ^ x[35];
  assign t[137] = t[165] ^ x[20];
  assign t[138] = t[166] ^ x[36];
  assign t[139] = t[167] ^ x[37];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[38];
  assign t[141] = t[169] ^ x[18];
  assign t[142] = t[170] ^ x[26];
  assign t[143] = t[171] ^ x[39];
  assign t[144] = t[172] ^ x[27];
  assign t[145] = t[173] ^ x[40];
  assign t[146] = t[174] ^ x[41];
  assign t[147] = t[175] ^ x[42];
  assign t[148] = t[176] ^ x[25];
  assign t[149] = t[177] ^ x[33];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[178] ^ x[43];
  assign t[151] = t[179] ^ x[34];
  assign t[152] = t[180] ^ x[44];
  assign t[153] = t[181] ^ x[45];
  assign t[154] = t[182] ^ x[46];
  assign t[155] = t[183] ^ x[32];
  assign t[156] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[157] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[158] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[159] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[164] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[165] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[166] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[167] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[168] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[169] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[16] = ~(t[76] | t[23]);
  assign t[170] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[171] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[172] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[173] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[174] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[175] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[176] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[177] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[178] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[179] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[180] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[181] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[182] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[183] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[77] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[78] | t[29]);
  assign t[21] = ~(t[79]);
  assign t[22] = ~(t[80]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[81]);
  assign t[25] = ~(t[82]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[83]);
  assign t[28] = ~(t[84]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[85]);
  assign t[31] = ~(t[79] | t[80]);
  assign t[32] = ~(t[86]);
  assign t[33] = ~(t[81] | t[82]);
  assign t[34] = ~(t[87]);
  assign t[35] = ~(t[83] | t[84]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[79] & t[22]);
  assign t[49] = ~(t[85] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[81] & t[25]);
  assign t[51] = ~(t[86] & t[55]);
  assign t[52] = ~(t[83] & t[28]);
  assign t[53] = ~(t[87] & t[56]);
  assign t[54] = ~(t[80] & t[21]);
  assign t[55] = ~(t[82] & t[24]);
  assign t[56] = ~(t[84] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[4] ? x[53] : x[52];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[15] | t[76];
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = t[17] | t[77];
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = t[19] | t[78];
  assign t[75] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[76] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[77] = (t[92] & ~t[93]) | (~t[92] & t[93]);
  assign t[78] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[79] = (t[90] & ~t[97] & ~t[99]) | (~t[96] & t[97] & ~t[98]) | (~t[90] & ~t[97] & t[99]) | (t[96] & t[97] & t[98]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[90] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[99]) | (~t[90] & ~t[97] & t[98]) | (t[96] & t[97] & t[99]);
  assign t[81] = (t[92] & ~t[101] & ~t[103]) | (~t[100] & t[101] & ~t[102]) | (~t[92] & ~t[101] & t[103]) | (t[100] & t[101] & t[102]);
  assign t[82] = (t[92] & ~t[101] & ~t[102]) | (~t[100] & t[101] & ~t[103]) | (~t[92] & ~t[101] & t[102]) | (t[100] & t[101] & t[103]);
  assign t[83] = (t[94] & ~t[105] & ~t[107]) | (~t[104] & t[105] & ~t[106]) | (~t[94] & ~t[105] & t[107]) | (t[104] & t[105] & t[106]);
  assign t[84] = (t[94] & ~t[105] & ~t[106]) | (~t[104] & t[105] & ~t[107]) | (~t[94] & ~t[105] & t[106]) | (t[104] & t[105] & t[107]);
  assign t[85] = (t[90] & ~t[98]) | (~t[90] & t[98]);
  assign t[86] = (t[92] & ~t[102]) | (~t[92] & t[102]);
  assign t[87] = (t[94] & ~t[106]) | (~t[94] & t[106]);
  assign t[88] = t[108] ^ x[12];
  assign t[89] = t[109] ^ x[13];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[110] ^ x[19];
  assign t[91] = t[111] ^ x[20];
  assign t[92] = t[112] ^ x[26];
  assign t[93] = t[113] ^ x[27];
  assign t[94] = t[114] ^ x[33];
  assign t[95] = t[115] ^ x[34];
  assign t[96] = t[116] ^ x[35];
  assign t[97] = t[117] ^ x[36];
  assign t[98] = t[118] ^ x[37];
  assign t[99] = t[119] ^ x[38];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57]) | (~t[0] & t[36] & ~t[57]) | (~t[0] & ~t[36] & t[57]) | (t[0] & t[36] & t[57]);
endmodule

module R2ind163(x, y);
 input [51:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[101] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[102] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[103] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[104] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[105] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[106] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[107] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[108] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[109] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[111] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[112] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[113] = t[141] ^ x[12];
  assign t[114] = t[142] ^ x[7];
  assign t[115] = t[143] ^ x[8];
  assign t[116] = t[144] ^ x[9];
  assign t[117] = t[145] ^ x[13];
  assign t[118] = t[146] ^ x[10];
  assign t[119] = t[147] ^ x[11];
  assign t[11] = ~x[2] & t[60];
  assign t[120] = t[148] ^ x[19];
  assign t[121] = t[149] ^ x[35];
  assign t[122] = t[150] ^ x[20];
  assign t[123] = t[151] ^ x[36];
  assign t[124] = t[152] ^ x[37];
  assign t[125] = t[153] ^ x[38];
  assign t[126] = t[154] ^ x[18];
  assign t[127] = t[155] ^ x[26];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[27];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[25];
  assign t[134] = t[162] ^ x[33];
  assign t[135] = t[163] ^ x[43];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[44];
  assign t[138] = t[166] ^ x[45];
  assign t[139] = t[167] ^ x[46];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[32];
  assign t[141] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[142] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[143] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[144] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[149] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[151] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[152] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[153] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[154] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[155] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[156] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[157] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[158] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[159] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[161] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[162] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[163] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[164] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[165] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[166] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[167] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[168] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[61] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[62] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[63] | t[29]);
  assign t[21] = ~(t[64]);
  assign t[22] = ~(t[65]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[66]);
  assign t[25] = ~(t[67]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[69]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[70]);
  assign t[31] = ~(t[64] | t[65]);
  assign t[32] = ~(t[71]);
  assign t[33] = ~(t[66] | t[67]);
  assign t[34] = ~(t[72]);
  assign t[35] = ~(t[68] | t[69]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[22] & t[30]);
  assign t[49] = ~(t[54] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[25] & t[32]);
  assign t[51] = ~(t[55] & t[62]);
  assign t[52] = ~(t[28] & t[34]);
  assign t[53] = ~(t[56] & t[63]);
  assign t[54] = ~(t[57] & t[21]);
  assign t[55] = ~(t[58] & t[24]);
  assign t[56] = ~(t[59] & t[27]);
  assign t[57] = ~(t[70] & t[65]);
  assign t[58] = ~(t[71] & t[67]);
  assign t[59] = ~(t[72] & t[69]);
  assign t[5] = t[8];
  assign t[60] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[61] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[62] = (t[77] & ~t[78]) | (~t[77] & t[78]);
  assign t[63] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[64] = (t[75] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[75] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[65] = (t[75] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[75] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[66] = (t[77] & ~t[86] & ~t[88]) | (~t[85] & t[86] & ~t[87]) | (~t[77] & ~t[86] & t[88]) | (t[85] & t[86] & t[87]);
  assign t[67] = (t[77] & ~t[86] & ~t[87]) | (~t[85] & t[86] & ~t[88]) | (~t[77] & ~t[86] & t[87]) | (t[85] & t[86] & t[88]);
  assign t[68] = (t[79] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[79] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[69] = (t[79] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[79] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[75] & ~t[83]) | (~t[75] & t[83]);
  assign t[71] = (t[77] & ~t[87]) | (~t[77] & t[87]);
  assign t[72] = (t[79] & ~t[91]) | (~t[79] & t[91]);
  assign t[73] = t[93] ^ x[12];
  assign t[74] = t[94] ^ x[13];
  assign t[75] = t[95] ^ x[19];
  assign t[76] = t[96] ^ x[20];
  assign t[77] = t[97] ^ x[26];
  assign t[78] = t[98] ^ x[27];
  assign t[79] = t[99] ^ x[33];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[34];
  assign t[81] = t[101] ^ x[35];
  assign t[82] = t[102] ^ x[36];
  assign t[83] = t[103] ^ x[37];
  assign t[84] = t[104] ^ x[38];
  assign t[85] = t[105] ^ x[39];
  assign t[86] = t[106] ^ x[40];
  assign t[87] = t[107] ^ x[41];
  assign t[88] = t[108] ^ x[42];
  assign t[89] = t[109] ^ x[43];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[110] ^ x[44];
  assign t[91] = t[111] ^ x[45];
  assign t[92] = t[112] ^ x[46];
  assign t[93] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[97] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[98] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[99] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind164(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[55] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[56] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[57] | t[29]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[61]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[62]);
  assign t[28] = ~(t[63]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[64]);
  assign t[31] = ~(t[58] | t[59]);
  assign t[32] = ~(t[65]);
  assign t[33] = ~(t[60] | t[61]);
  assign t[34] = ~(t[66]);
  assign t[35] = ~(t[62] | t[63]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[22] & t[30]);
  assign t[49] = t[15] | t[55];
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[25] & t[32]);
  assign t[51] = t[17] | t[56];
  assign t[52] = ~(t[28] & t[34]);
  assign t[53] = t[19] | t[57];
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[59] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[5] = t[8];
  assign t[60] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[61] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[62] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[63] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[64] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[65] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[66] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind165(x, y);
 input [51:0] x;
 output y;

 wire [165:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[101] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[102] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[103] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[104] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[105] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[106] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[107] = (t[117] & t[118] & ~t[119] & t[120] & ~t[121] & ~t[123]) | (t[117] & ~t[119] & ~t[120] & t[121] & ~t[122] & t[123]) | (~t[118] & t[119] & ~t[120] & ~t[121] & ~t[123]) | (~t[117] & t[119] & ~t[120] & ~t[121] & ~t[122]) | (~t[117] & ~t[118] & t[119] & ~t[122] & ~t[123]) | (~t[117] & t[119] & t[120] & ~t[121] & t[122]) | (t[119] & ~t[120] & t[122] & ~t[123]);
  assign t[108] = (t[124] & t[125] & ~t[126] & t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[126] & ~t[127] & t[128] & ~t[129] & t[130]) | (~t[125] & t[126] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[125] & t[126] & ~t[129] & ~t[130]) | (~t[124] & t[126] & t[127] & ~t[128] & t[129]) | (t[126] & ~t[127] & t[129] & ~t[130]);
  assign t[109] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[12];
  assign t[111] = t[139] ^ x[7];
  assign t[112] = t[140] ^ x[8];
  assign t[113] = t[141] ^ x[9];
  assign t[114] = t[142] ^ x[13];
  assign t[115] = t[143] ^ x[10];
  assign t[116] = t[144] ^ x[11];
  assign t[117] = t[145] ^ x[19];
  assign t[118] = t[146] ^ x[20];
  assign t[119] = t[147] ^ x[49];
  assign t[11] = ~x[2] & t[57];
  assign t[120] = t[148] ^ x[21];
  assign t[121] = t[149] ^ x[22];
  assign t[122] = t[150] ^ x[23];
  assign t[123] = t[151] ^ x[18];
  assign t[124] = t[152] ^ x[29];
  assign t[125] = t[153] ^ x[30];
  assign t[126] = t[154] ^ x[50];
  assign t[127] = t[155] ^ x[31];
  assign t[128] = t[156] ^ x[32];
  assign t[129] = t[157] ^ x[33];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[28];
  assign t[131] = t[159] ^ x[39];
  assign t[132] = t[160] ^ x[40];
  assign t[133] = t[161] ^ x[51];
  assign t[134] = t[162] ^ x[41];
  assign t[135] = t[163] ^ x[42];
  assign t[136] = t[164] ^ x[43];
  assign t[137] = t[165] ^ x[38];
  assign t[138] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[139] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[141] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[142] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[146] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[147] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[148] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[149] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[151] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[152] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[153] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[154] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[155] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[156] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[157] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[158] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[159] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[15] = ~(t[58] & t[21]);
  assign t[160] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[161] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[162] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[163] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[164] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[165] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[59] & t[22]);
  assign t[17] = ~(t[60] & t[23]);
  assign t[18] = ~(t[61] & t[24]);
  assign t[19] = ~(t[62] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[63] & t[26]);
  assign t[21] = ~(t[64]);
  assign t[22] = ~(t[64] & t[27]);
  assign t[23] = ~(t[65]);
  assign t[24] = ~(t[65] & t[28]);
  assign t[25] = ~(t[66]);
  assign t[26] = ~(t[66] & t[29]);
  assign t[27] = ~(t[58]);
  assign t[28] = ~(t[60]);
  assign t[29] = ~(t[62]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[4] ? x[45] : x[44];
  assign t[33] = ~(t[34] ^ t[35]);
  assign t[34] = t[36];
  assign t[35] = ~(t[37] ^ t[38]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = ~(t[49] & t[67]);
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = ~(t[51] & t[68]);
  assign t[46] = ~(t[25] & t[52]);
  assign t[47] = ~(t[53] & t[69]);
  assign t[48] = ~(t[59]);
  assign t[49] = ~(t[54] & t[27]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[61]);
  assign t[51] = ~(t[55] & t[28]);
  assign t[52] = ~(t[63]);
  assign t[53] = ~(t[56] & t[29]);
  assign t[54] = ~(t[59] & t[64]);
  assign t[55] = ~(t[61] & t[65]);
  assign t[56] = ~(t[63] & t[66]);
  assign t[57] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[58] = (t[72] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[72] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[59] = (t[72] & ~t[75]) | (~t[72] & t[75]);
  assign t[5] = t[8];
  assign t[60] = (t[77] & ~t[79] & ~t[81]) | (~t[78] & t[79] & ~t[80]) | (~t[77] & ~t[79] & t[81]) | (t[78] & t[79] & t[80]);
  assign t[61] = (t[77] & ~t[80]) | (~t[77] & t[80]);
  assign t[62] = (t[82] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[82] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[63] = (t[82] & ~t[85]) | (~t[82] & t[85]);
  assign t[64] = (t[72] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[72] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[65] = (t[77] & ~t[79] & ~t[80]) | (~t[78] & t[79] & ~t[81]) | (~t[77] & ~t[79] & t[80]) | (t[78] & t[79] & t[81]);
  assign t[66] = (t[82] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[82] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[67] = (t[72] & ~t[87]) | (~t[72] & t[87]);
  assign t[68] = (t[77] & ~t[88]) | (~t[77] & t[88]);
  assign t[69] = (t[82] & ~t[89]) | (~t[82] & t[89]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[12];
  assign t[71] = t[91] ^ x[13];
  assign t[72] = t[92] ^ x[19];
  assign t[73] = t[93] ^ x[20];
  assign t[74] = t[94] ^ x[21];
  assign t[75] = t[95] ^ x[22];
  assign t[76] = t[96] ^ x[23];
  assign t[77] = t[97] ^ x[29];
  assign t[78] = t[98] ^ x[30];
  assign t[79] = t[99] ^ x[31];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[32];
  assign t[81] = t[101] ^ x[33];
  assign t[82] = t[102] ^ x[39];
  assign t[83] = t[103] ^ x[40];
  assign t[84] = t[104] ^ x[41];
  assign t[85] = t[105] ^ x[42];
  assign t[86] = t[106] ^ x[43];
  assign t[87] = t[107] ^ x[49];
  assign t[88] = t[108] ^ x[50];
  assign t[89] = t[109] ^ x[51];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[110] & ~t[112] & ~t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[113] & ~t[114] & ~t[116]) | (t[110] & ~t[111] & ~t[112] & ~t[115] & ~t[116]) | (~t[110] & t[111] & t[112] & t[113] & ~t[116]) | (~t[110] & t[111] & t[114] & t[115] & ~t[116]) | (t[110] & ~t[112] & ~t[114] & t[116]) | (~t[110] & t[112] & t[114] & t[116]);
  assign t[91] = (t[110] & t[111] & ~t[112] & ~t[114] & t[115] & ~t[116]) | (t[110] & t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[116]) | (~t[110] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[110] & ~t[111] & ~t[113] & t[114] & ~t[116]) | (~t[110] & ~t[112] & t[113] & t[114] & t[115]) | (t[113] & t[114] & ~t[115] & ~t[116]);
  assign t[92] = (t[117] & ~t[119] & ~t[120] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & ~t[120] & ~t[121] & ~t[123]) | (t[117] & ~t[118] & ~t[119] & ~t[122] & ~t[123]) | (~t[117] & t[118] & t[119] & t[120] & ~t[123]) | (~t[117] & t[118] & t[121] & t[122] & ~t[123]) | (t[117] & ~t[119] & ~t[121] & t[123]) | (~t[117] & t[119] & t[121] & t[123]);
  assign t[93] = (t[118] & ~t[119] & ~t[120] & ~t[121] & ~t[122]) | (~t[117] & t[118] & ~t[120] & ~t[121] & ~t[123]) | (~t[117] & t[118] & ~t[119] & ~t[122] & ~t[123]) | (t[117] & ~t[118] & t[119] & t[120] & ~t[123]) | (t[117] & ~t[118] & t[121] & t[122] & ~t[123]) | (t[118] & ~t[120] & ~t[122] & t[123]) | (~t[118] & t[120] & t[122] & t[123]);
  assign t[94] = (t[117] & t[118] & t[119] & ~t[120] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[120] & ~t[121] & t[122] & t[123]) | (~t[118] & ~t[119] & t[120] & ~t[121] & ~t[122]) | (~t[117] & ~t[119] & t[120] & ~t[122] & ~t[123]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[123]) | (~t[118] & t[119] & t[120] & t[121] & ~t[122]) | (~t[119] & t[120] & t[121] & ~t[123]);
  assign t[95] = (t[117] & t[118] & ~t[119] & ~t[121] & t[122] & ~t[123]) | (t[117] & t[119] & ~t[120] & ~t[121] & ~t[122] & t[123]) | (~t[118] & ~t[119] & t[121] & ~t[122] & ~t[123]) | (~t[117] & ~t[119] & ~t[120] & t[121] & ~t[122]) | (~t[117] & ~t[118] & ~t[120] & t[121] & ~t[123]) | (~t[117] & ~t[119] & t[120] & t[121] & t[122]) | (t[120] & t[121] & ~t[122] & ~t[123]);
  assign t[96] = (t[117] & t[118] & ~t[120] & t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & t[120] & ~t[121] & ~t[122] & t[123]) | (~t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[117] & ~t[118] & ~t[119] & t[122] & ~t[123]) | (~t[118] & t[119] & ~t[120] & t[121] & t[122]) | (t[119] & ~t[121] & t[122] & ~t[123]);
  assign t[97] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[98] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[99] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[30]) | (~t[0] & t[30]);
endmodule

module R2ind166(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[101] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[102] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[103] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[104] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[105] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[106] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[20];
  assign t[116] = t[144] ^ x[49];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[23];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[30];
  assign t[123] = t[151] ^ x[50];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[33];
  assign t[127] = t[155] ^ x[28];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[40];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[51];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[43];
  assign t[134] = t[162] ^ x[38];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[151] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[152] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[153] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[154] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[155] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[156] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[157] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[158] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[159] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[15] = ~(t[55] & t[21]);
  assign t[160] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[161] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[162] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[56] & t[22]);
  assign t[17] = ~(t[57] & t[23]);
  assign t[18] = ~(t[58] & t[24]);
  assign t[19] = ~(t[59] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[60] & t[26]);
  assign t[21] = ~(t[61]);
  assign t[22] = ~(t[61] & t[27]);
  assign t[23] = ~(t[62]);
  assign t[24] = ~(t[62] & t[28]);
  assign t[25] = ~(t[63]);
  assign t[26] = ~(t[63] & t[29]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[59]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[4] ? x[45] : x[44];
  assign t[33] = ~(t[34] ^ t[35]);
  assign t[34] = t[36];
  assign t[35] = ~(t[37] ^ t[38]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = t[49] | t[64];
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = t[51] | t[65];
  assign t[46] = ~(t[25] & t[52]);
  assign t[47] = t[53] | t[66];
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[27] | t[21]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[58]);
  assign t[51] = ~(t[28] | t[23]);
  assign t[52] = ~(t[60]);
  assign t[53] = ~(t[29] | t[25]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[69] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = (t[69] & ~t[72]) | (~t[69] & t[72]);
  assign t[57] = (t[74] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[74] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[58] = (t[74] & ~t[77]) | (~t[74] & t[77]);
  assign t[59] = (t[79] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[79] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[5] = t[8];
  assign t[60] = (t[79] & ~t[82]) | (~t[79] & t[82]);
  assign t[61] = (t[69] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[69] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[62] = (t[74] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[74] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[63] = (t[79] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[79] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[64] = (t[69] & ~t[84]) | (~t[69] & t[84]);
  assign t[65] = (t[74] & ~t[85]) | (~t[74] & t[85]);
  assign t[66] = (t[79] & ~t[86]) | (~t[79] & t[86]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[21];
  assign t[72] = t[92] ^ x[22];
  assign t[73] = t[93] ^ x[23];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[31];
  assign t[77] = t[97] ^ x[32];
  assign t[78] = t[98] ^ x[33];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[49];
  assign t[85] = t[105] ^ x[50];
  assign t[86] = t[106] ^ x[51];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[91] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[92] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[93] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[94] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[95] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[96] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[97] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[98] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[99] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[30]) | (~t[0] & t[30]);
endmodule

module R2ind167(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[23] & t[55]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[56]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[57]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[61]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[62]);
  assign t[28] = ~(t[63]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[59] & t[58]);
  assign t[31] = ~(t[64]);
  assign t[32] = ~(t[61] & t[60]);
  assign t[33] = ~(t[65]);
  assign t[34] = ~(t[63] & t[62]);
  assign t[35] = ~(t[66]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[15] & t[48]);
  assign t[46] = ~(t[17] & t[49]);
  assign t[47] = ~(t[19] & t[50]);
  assign t[48] = t[51] | t[55];
  assign t[49] = t[52] | t[56];
  assign t[4] = ~(t[7]);
  assign t[50] = t[53] | t[57];
  assign t[51] = ~(t[31] | t[21]);
  assign t[52] = ~(t[33] | t[24]);
  assign t[53] = ~(t[35] | t[27]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[59] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[5] = t[8];
  assign t[60] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[61] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[62] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[63] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[64] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[65] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[66] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind168(x, y);
 input [56:0] x;
 output y;

 wire [189:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[33];
  assign t[101] = t[121] ^ x[34];
  assign t[102] = t[122] ^ x[35];
  assign t[103] = t[123] ^ x[36];
  assign t[104] = t[124] ^ x[37];
  assign t[105] = t[125] ^ x[38];
  assign t[106] = t[126] ^ x[39];
  assign t[107] = t[127] ^ x[40];
  assign t[108] = t[128] ^ x[41];
  assign t[109] = t[129] ^ x[42];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[130] ^ x[43];
  assign t[111] = t[131] ^ x[44];
  assign t[112] = t[132] ^ x[45];
  assign t[113] = t[133] ^ x[46];
  assign t[114] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[115] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[116] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[117] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[118] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[119] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[11] = ~x[2] & t[81];
  assign t[120] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[121] = (t[155] & t[156] & ~t[157] & t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[157] & ~t[158] & t[159] & ~t[160] & t[161]) | (~t[156] & t[157] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[156] & t[157] & ~t[160] & ~t[161]) | (~t[155] & t[157] & t[158] & ~t[159] & t[160]) | (t[157] & ~t[158] & t[160] & ~t[161]);
  assign t[122] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[123] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[124] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[125] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[126] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[127] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[128] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[129] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (t[156] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & t[156] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[156] & ~t[157] & ~t[160] & ~t[161]) | (t[155] & ~t[156] & t[157] & t[158] & ~t[161]) | (t[155] & ~t[156] & t[159] & t[160] & ~t[161]) | (t[156] & ~t[158] & ~t[160] & t[161]) | (~t[156] & t[158] & t[160] & t[161]);
  assign t[131] = (t[155] & t[156] & t[157] & ~t[158] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & ~t[158] & ~t[159] & t[160] & t[161]) | (~t[156] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[157] & t[158] & ~t[160] & ~t[161]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[161]) | (~t[156] & t[157] & t[158] & t[159] & ~t[160]) | (~t[157] & t[158] & t[159] & ~t[161]);
  assign t[132] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[133] = (t[155] & t[156] & ~t[158] & t[159] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[158] & ~t[159] & t[160] & ~t[161]) | (~t[155] & ~t[156] & ~t[157] & t[160] & ~t[161]) | (~t[156] & t[157] & ~t[158] & t[159] & t[160]) | (t[157] & ~t[159] & t[160] & ~t[161]);
  assign t[134] = t[162] ^ x[12];
  assign t[135] = t[163] ^ x[7];
  assign t[136] = t[164] ^ x[8];
  assign t[137] = t[165] ^ x[9];
  assign t[138] = t[166] ^ x[13];
  assign t[139] = t[167] ^ x[10];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[11];
  assign t[141] = t[169] ^ x[19];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[20];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[18];
  assign t[148] = t[176] ^ x[26];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[178] ^ x[27];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[25];
  assign t[155] = t[183] ^ x[33];
  assign t[156] = t[184] ^ x[43];
  assign t[157] = t[185] ^ x[34];
  assign t[158] = t[186] ^ x[44];
  assign t[159] = t[187] ^ x[45];
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = t[188] ^ x[46];
  assign t[161] = t[189] ^ x[32];
  assign t[162] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[163] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[164] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[165] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[166] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[167] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[168] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[169] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[16] = ~(t[82] | t[23]);
  assign t[170] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[171] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[172] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[173] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[174] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[175] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[176] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[177] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[178] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[179] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[180] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[181] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[182] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[183] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[184] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[185] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[186] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[187] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[188] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[189] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[83] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[84] | t[29]);
  assign t[21] = ~(t[85]);
  assign t[22] = ~(t[86]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[87]);
  assign t[25] = ~(t[88]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[89]);
  assign t[28] = ~(t[90]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[91]);
  assign t[31] = ~(t[85] | t[86]);
  assign t[32] = ~(t[92]);
  assign t[33] = ~(t[87] | t[88]);
  assign t[34] = ~(t[93]);
  assign t[35] = ~(t[89] | t[90]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[11] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[85] & t[22]);
  assign t[49] = ~(t[91] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[87] & t[25]);
  assign t[51] = ~(t[92] & t[55]);
  assign t[52] = ~(t[89] & t[28]);
  assign t[53] = ~(t[93] & t[56]);
  assign t[54] = ~(t[86] & t[21]);
  assign t[55] = ~(t[88] & t[24]);
  assign t[56] = ~(t[90] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[11] ? x[53] : x[52];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = ~(t[75] & t[82]);
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = ~(t[76] & t[83]);
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = ~(t[77] & t[84]);
  assign t[75] = ~(t[78] & t[21]);
  assign t[76] = ~(t[79] & t[24]);
  assign t[77] = ~(t[80] & t[27]);
  assign t[78] = ~(t[91] & t[86]);
  assign t[79] = ~(t[92] & t[88]);
  assign t[7] = ~(t[11]);
  assign t[80] = ~(t[93] & t[90]);
  assign t[81] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[82] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[83] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[84] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[85] = (t[96] & ~t[103] & ~t[105]) | (~t[102] & t[103] & ~t[104]) | (~t[96] & ~t[103] & t[105]) | (t[102] & t[103] & t[104]);
  assign t[86] = (t[96] & ~t[103] & ~t[104]) | (~t[102] & t[103] & ~t[105]) | (~t[96] & ~t[103] & t[104]) | (t[102] & t[103] & t[105]);
  assign t[87] = (t[98] & ~t[107] & ~t[109]) | (~t[106] & t[107] & ~t[108]) | (~t[98] & ~t[107] & t[109]) | (t[106] & t[107] & t[108]);
  assign t[88] = (t[98] & ~t[107] & ~t[108]) | (~t[106] & t[107] & ~t[109]) | (~t[98] & ~t[107] & t[108]) | (t[106] & t[107] & t[109]);
  assign t[89] = (t[100] & ~t[111] & ~t[113]) | (~t[110] & t[111] & ~t[112]) | (~t[100] & ~t[111] & t[113]) | (t[110] & t[111] & t[112]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[100] & ~t[111] & ~t[112]) | (~t[110] & t[111] & ~t[113]) | (~t[100] & ~t[111] & t[112]) | (t[110] & t[111] & t[113]);
  assign t[91] = (t[96] & ~t[104]) | (~t[96] & t[104]);
  assign t[92] = (t[98] & ~t[108]) | (~t[98] & t[108]);
  assign t[93] = (t[100] & ~t[112]) | (~t[100] & t[112]);
  assign t[94] = t[114] ^ x[12];
  assign t[95] = t[115] ^ x[13];
  assign t[96] = t[116] ^ x[19];
  assign t[97] = t[117] ^ x[20];
  assign t[98] = t[118] ^ x[26];
  assign t[99] = t[119] ^ x[27];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57]) | (~t[0] & t[36] & ~t[57]) | (~t[0] & ~t[36] & t[57]) | (t[0] & t[36] & t[57]);
endmodule

module R2ind169(x, y);
 input [56:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[39];
  assign t[101] = t[121] ^ x[40];
  assign t[102] = t[122] ^ x[41];
  assign t[103] = t[123] ^ x[42];
  assign t[104] = t[124] ^ x[43];
  assign t[105] = t[125] ^ x[44];
  assign t[106] = t[126] ^ x[45];
  assign t[107] = t[127] ^ x[46];
  assign t[108] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[109] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (t[135] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[136] & ~t[137] & ~t[140] & ~t[141]) | (~t[135] & t[136] & t[137] & t[138] & ~t[141]) | (~t[135] & t[136] & t[139] & t[140] & ~t[141]) | (t[135] & ~t[137] & ~t[139] & t[141]) | (~t[135] & t[137] & t[139] & t[141]);
  assign t[111] = (t[135] & t[136] & ~t[137] & t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[137] & ~t[138] & t[139] & ~t[140] & t[141]) | (~t[136] & t[137] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[136] & t[137] & ~t[140] & ~t[141]) | (~t[135] & t[137] & t[138] & ~t[139] & t[140]) | (t[137] & ~t[138] & t[140] & ~t[141]);
  assign t[112] = (t[142] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[143] & ~t[144] & ~t[147] & ~t[148]) | (~t[142] & t[143] & t[144] & t[145] & ~t[148]) | (~t[142] & t[143] & t[146] & t[147] & ~t[148]) | (t[142] & ~t[144] & ~t[146] & t[148]) | (~t[142] & t[144] & t[146] & t[148]);
  assign t[113] = (t[142] & t[143] & ~t[144] & t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[144] & ~t[145] & t[146] & ~t[147] & t[148]) | (~t[143] & t[144] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[143] & t[144] & ~t[147] & ~t[148]) | (~t[142] & t[144] & t[145] & ~t[146] & t[147]) | (t[144] & ~t[145] & t[147] & ~t[148]);
  assign t[114] = (t[149] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[150] & ~t[151] & ~t[154] & ~t[155]) | (~t[149] & t[150] & t[151] & t[152] & ~t[155]) | (~t[149] & t[150] & t[153] & t[154] & ~t[155]) | (t[149] & ~t[151] & ~t[153] & t[155]) | (~t[149] & t[151] & t[153] & t[155]);
  assign t[115] = (t[149] & t[150] & ~t[151] & t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[151] & ~t[152] & t[153] & ~t[154] & t[155]) | (~t[150] & t[151] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[150] & t[151] & ~t[154] & ~t[155]) | (~t[149] & t[151] & t[152] & ~t[153] & t[154]) | (t[151] & ~t[152] & t[154] & ~t[155]);
  assign t[116] = (t[136] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & t[136] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[136] & ~t[137] & ~t[140] & ~t[141]) | (t[135] & ~t[136] & t[137] & t[138] & ~t[141]) | (t[135] & ~t[136] & t[139] & t[140] & ~t[141]) | (t[136] & ~t[138] & ~t[140] & t[141]) | (~t[136] & t[138] & t[140] & t[141]);
  assign t[117] = (t[135] & t[136] & t[137] & ~t[138] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & ~t[138] & ~t[139] & t[140] & t[141]) | (~t[136] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[137] & t[138] & ~t[140] & ~t[141]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[141]) | (~t[136] & t[137] & t[138] & t[139] & ~t[140]) | (~t[137] & t[138] & t[139] & ~t[141]);
  assign t[118] = (t[135] & t[136] & ~t[137] & ~t[139] & t[140] & ~t[141]) | (t[135] & t[137] & ~t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & t[139] & ~t[140] & ~t[141]) | (~t[135] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[135] & ~t[136] & ~t[138] & t[139] & ~t[141]) | (~t[135] & ~t[137] & t[138] & t[139] & t[140]) | (t[138] & t[139] & ~t[140] & ~t[141]);
  assign t[119] = (t[135] & t[136] & ~t[138] & t[139] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[138] & ~t[139] & t[140] & ~t[141]) | (~t[135] & ~t[136] & ~t[137] & t[140] & ~t[141]) | (~t[136] & t[137] & ~t[138] & t[139] & t[140]) | (t[137] & ~t[139] & t[140] & ~t[141]);
  assign t[11] = ~x[2] & t[75];
  assign t[120] = (t[143] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & t[143] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[143] & ~t[144] & ~t[147] & ~t[148]) | (t[142] & ~t[143] & t[144] & t[145] & ~t[148]) | (t[142] & ~t[143] & t[146] & t[147] & ~t[148]) | (t[143] & ~t[145] & ~t[147] & t[148]) | (~t[143] & t[145] & t[147] & t[148]);
  assign t[121] = (t[142] & t[143] & t[144] & ~t[145] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & ~t[145] & ~t[146] & t[147] & t[148]) | (~t[143] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[144] & t[145] & ~t[147] & ~t[148]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[148]) | (~t[143] & t[144] & t[145] & t[146] & ~t[147]) | (~t[144] & t[145] & t[146] & ~t[148]);
  assign t[122] = (t[142] & t[143] & ~t[144] & ~t[146] & t[147] & ~t[148]) | (t[142] & t[144] & ~t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & t[146] & ~t[147] & ~t[148]) | (~t[142] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[142] & ~t[143] & ~t[145] & t[146] & ~t[148]) | (~t[142] & ~t[144] & t[145] & t[146] & t[147]) | (t[145] & t[146] & ~t[147] & ~t[148]);
  assign t[123] = (t[142] & t[143] & ~t[145] & t[146] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[145] & ~t[146] & t[147] & ~t[148]) | (~t[142] & ~t[143] & ~t[144] & t[147] & ~t[148]) | (~t[143] & t[144] & ~t[145] & t[146] & t[147]) | (t[144] & ~t[146] & t[147] & ~t[148]);
  assign t[124] = (t[150] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & t[150] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[150] & ~t[151] & ~t[154] & ~t[155]) | (t[149] & ~t[150] & t[151] & t[152] & ~t[155]) | (t[149] & ~t[150] & t[153] & t[154] & ~t[155]) | (t[150] & ~t[152] & ~t[154] & t[155]) | (~t[150] & t[152] & t[154] & t[155]);
  assign t[125] = (t[149] & t[150] & t[151] & ~t[152] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & ~t[152] & ~t[153] & t[154] & t[155]) | (~t[150] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[151] & t[152] & ~t[154] & ~t[155]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[155]) | (~t[150] & t[151] & t[152] & t[153] & ~t[154]) | (~t[151] & t[152] & t[153] & ~t[155]);
  assign t[126] = (t[149] & t[150] & ~t[151] & ~t[153] & t[154] & ~t[155]) | (t[149] & t[151] & ~t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & t[153] & ~t[154] & ~t[155]) | (~t[149] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[149] & ~t[150] & ~t[152] & t[153] & ~t[155]) | (~t[149] & ~t[151] & t[152] & t[153] & t[154]) | (t[152] & t[153] & ~t[154] & ~t[155]);
  assign t[127] = (t[149] & t[150] & ~t[152] & t[153] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[152] & ~t[153] & t[154] & ~t[155]) | (~t[149] & ~t[150] & ~t[151] & t[154] & ~t[155]) | (~t[150] & t[151] & ~t[152] & t[153] & t[154]) | (t[151] & ~t[153] & t[154] & ~t[155]);
  assign t[128] = t[156] ^ x[12];
  assign t[129] = t[157] ^ x[7];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[8];
  assign t[131] = t[159] ^ x[9];
  assign t[132] = t[160] ^ x[13];
  assign t[133] = t[161] ^ x[10];
  assign t[134] = t[162] ^ x[11];
  assign t[135] = t[163] ^ x[19];
  assign t[136] = t[164] ^ x[35];
  assign t[137] = t[165] ^ x[20];
  assign t[138] = t[166] ^ x[36];
  assign t[139] = t[167] ^ x[37];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[38];
  assign t[141] = t[169] ^ x[18];
  assign t[142] = t[170] ^ x[26];
  assign t[143] = t[171] ^ x[39];
  assign t[144] = t[172] ^ x[27];
  assign t[145] = t[173] ^ x[40];
  assign t[146] = t[174] ^ x[41];
  assign t[147] = t[175] ^ x[42];
  assign t[148] = t[176] ^ x[25];
  assign t[149] = t[177] ^ x[33];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[178] ^ x[43];
  assign t[151] = t[179] ^ x[34];
  assign t[152] = t[180] ^ x[44];
  assign t[153] = t[181] ^ x[45];
  assign t[154] = t[182] ^ x[46];
  assign t[155] = t[183] ^ x[32];
  assign t[156] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[157] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[158] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[159] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[164] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[165] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[166] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[167] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[168] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[169] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[16] = ~(t[76] | t[23]);
  assign t[170] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[171] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[172] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[173] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[174] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[175] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[176] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[177] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[178] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[179] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[180] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[181] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[182] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[183] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[77] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[78] | t[29]);
  assign t[21] = ~(t[79]);
  assign t[22] = ~(t[80]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[81]);
  assign t[25] = ~(t[82]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[83]);
  assign t[28] = ~(t[84]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[85]);
  assign t[31] = ~(t[79] | t[80]);
  assign t[32] = ~(t[86]);
  assign t[33] = ~(t[81] | t[82]);
  assign t[34] = ~(t[87]);
  assign t[35] = ~(t[83] | t[84]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[11] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[79] & t[22]);
  assign t[49] = ~(t[85] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[81] & t[25]);
  assign t[51] = ~(t[86] & t[55]);
  assign t[52] = ~(t[83] & t[28]);
  assign t[53] = ~(t[87] & t[56]);
  assign t[54] = ~(t[80] & t[21]);
  assign t[55] = ~(t[82] & t[24]);
  assign t[56] = ~(t[84] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[4] ? x[53] : x[52];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[15] | t[76];
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = t[17] | t[77];
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = t[19] | t[78];
  assign t[75] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[76] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[77] = (t[92] & ~t[93]) | (~t[92] & t[93]);
  assign t[78] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[79] = (t[90] & ~t[97] & ~t[99]) | (~t[96] & t[97] & ~t[98]) | (~t[90] & ~t[97] & t[99]) | (t[96] & t[97] & t[98]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[90] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[99]) | (~t[90] & ~t[97] & t[98]) | (t[96] & t[97] & t[99]);
  assign t[81] = (t[92] & ~t[101] & ~t[103]) | (~t[100] & t[101] & ~t[102]) | (~t[92] & ~t[101] & t[103]) | (t[100] & t[101] & t[102]);
  assign t[82] = (t[92] & ~t[101] & ~t[102]) | (~t[100] & t[101] & ~t[103]) | (~t[92] & ~t[101] & t[102]) | (t[100] & t[101] & t[103]);
  assign t[83] = (t[94] & ~t[105] & ~t[107]) | (~t[104] & t[105] & ~t[106]) | (~t[94] & ~t[105] & t[107]) | (t[104] & t[105] & t[106]);
  assign t[84] = (t[94] & ~t[105] & ~t[106]) | (~t[104] & t[105] & ~t[107]) | (~t[94] & ~t[105] & t[106]) | (t[104] & t[105] & t[107]);
  assign t[85] = (t[90] & ~t[98]) | (~t[90] & t[98]);
  assign t[86] = (t[92] & ~t[102]) | (~t[92] & t[102]);
  assign t[87] = (t[94] & ~t[106]) | (~t[94] & t[106]);
  assign t[88] = t[108] ^ x[12];
  assign t[89] = t[109] ^ x[13];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[110] ^ x[19];
  assign t[91] = t[111] ^ x[20];
  assign t[92] = t[112] ^ x[26];
  assign t[93] = t[113] ^ x[27];
  assign t[94] = t[114] ^ x[33];
  assign t[95] = t[115] ^ x[34];
  assign t[96] = t[116] ^ x[35];
  assign t[97] = t[117] ^ x[36];
  assign t[98] = t[118] ^ x[37];
  assign t[99] = t[119] ^ x[38];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57]) | (~t[0] & t[36] & ~t[57]) | (~t[0] & ~t[36] & t[57]) | (t[0] & t[36] & t[57]);
endmodule

module R2ind170(x, y);
 input [51:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[101] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[102] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[103] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[104] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[105] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[106] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[107] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[108] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[109] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[111] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[112] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[113] = t[141] ^ x[12];
  assign t[114] = t[142] ^ x[7];
  assign t[115] = t[143] ^ x[8];
  assign t[116] = t[144] ^ x[9];
  assign t[117] = t[145] ^ x[13];
  assign t[118] = t[146] ^ x[10];
  assign t[119] = t[147] ^ x[11];
  assign t[11] = ~x[2] & t[60];
  assign t[120] = t[148] ^ x[19];
  assign t[121] = t[149] ^ x[35];
  assign t[122] = t[150] ^ x[20];
  assign t[123] = t[151] ^ x[36];
  assign t[124] = t[152] ^ x[37];
  assign t[125] = t[153] ^ x[38];
  assign t[126] = t[154] ^ x[18];
  assign t[127] = t[155] ^ x[26];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[27];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[25];
  assign t[134] = t[162] ^ x[33];
  assign t[135] = t[163] ^ x[43];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[44];
  assign t[138] = t[166] ^ x[45];
  assign t[139] = t[167] ^ x[46];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[32];
  assign t[141] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[142] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[143] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[144] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[149] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[151] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[152] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[153] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[154] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[155] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[156] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[157] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[158] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[159] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[161] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[162] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[163] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[164] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[165] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[166] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[167] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[168] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[61] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[62] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[63] | t[29]);
  assign t[21] = ~(t[64]);
  assign t[22] = ~(t[65]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[66]);
  assign t[25] = ~(t[67]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[69]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[70]);
  assign t[31] = ~(t[64] | t[65]);
  assign t[32] = ~(t[71]);
  assign t[33] = ~(t[66] | t[67]);
  assign t[34] = ~(t[72]);
  assign t[35] = ~(t[68] | t[69]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[11] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[22] & t[30]);
  assign t[49] = ~(t[54] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[25] & t[32]);
  assign t[51] = ~(t[55] & t[62]);
  assign t[52] = ~(t[28] & t[34]);
  assign t[53] = ~(t[56] & t[63]);
  assign t[54] = ~(t[57] & t[21]);
  assign t[55] = ~(t[58] & t[24]);
  assign t[56] = ~(t[59] & t[27]);
  assign t[57] = ~(t[70] & t[65]);
  assign t[58] = ~(t[71] & t[67]);
  assign t[59] = ~(t[72] & t[69]);
  assign t[5] = t[8];
  assign t[60] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[61] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[62] = (t[77] & ~t[78]) | (~t[77] & t[78]);
  assign t[63] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[64] = (t[75] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[75] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[65] = (t[75] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[75] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[66] = (t[77] & ~t[86] & ~t[88]) | (~t[85] & t[86] & ~t[87]) | (~t[77] & ~t[86] & t[88]) | (t[85] & t[86] & t[87]);
  assign t[67] = (t[77] & ~t[86] & ~t[87]) | (~t[85] & t[86] & ~t[88]) | (~t[77] & ~t[86] & t[87]) | (t[85] & t[86] & t[88]);
  assign t[68] = (t[79] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[79] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[69] = (t[79] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[79] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[75] & ~t[83]) | (~t[75] & t[83]);
  assign t[71] = (t[77] & ~t[87]) | (~t[77] & t[87]);
  assign t[72] = (t[79] & ~t[91]) | (~t[79] & t[91]);
  assign t[73] = t[93] ^ x[12];
  assign t[74] = t[94] ^ x[13];
  assign t[75] = t[95] ^ x[19];
  assign t[76] = t[96] ^ x[20];
  assign t[77] = t[97] ^ x[26];
  assign t[78] = t[98] ^ x[27];
  assign t[79] = t[99] ^ x[33];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[34];
  assign t[81] = t[101] ^ x[35];
  assign t[82] = t[102] ^ x[36];
  assign t[83] = t[103] ^ x[37];
  assign t[84] = t[104] ^ x[38];
  assign t[85] = t[105] ^ x[39];
  assign t[86] = t[106] ^ x[40];
  assign t[87] = t[107] ^ x[41];
  assign t[88] = t[108] ^ x[42];
  assign t[89] = t[109] ^ x[43];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[110] ^ x[44];
  assign t[91] = t[111] ^ x[45];
  assign t[92] = t[112] ^ x[46];
  assign t[93] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[97] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[98] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[99] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind171(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[55] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[56] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[57] | t[29]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[61]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[62]);
  assign t[28] = ~(t[63]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[64]);
  assign t[31] = ~(t[58] | t[59]);
  assign t[32] = ~(t[65]);
  assign t[33] = ~(t[60] | t[61]);
  assign t[34] = ~(t[66]);
  assign t[35] = ~(t[62] | t[63]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[22] & t[30]);
  assign t[49] = t[15] | t[55];
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[25] & t[32]);
  assign t[51] = t[17] | t[56];
  assign t[52] = ~(t[28] & t[34]);
  assign t[53] = t[19] | t[57];
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[59] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[5] = t[8];
  assign t[60] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[61] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[62] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[63] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[64] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[65] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[66] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind172(x, y);
 input [51:0] x;
 output y;

 wire [163:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[129] & ~t[131] & ~t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[132] & ~t[133] & ~t[135]) | (t[129] & ~t[130] & ~t[131] & ~t[134] & ~t[135]) | (~t[129] & t[130] & t[131] & t[132] & ~t[135]) | (~t[129] & t[130] & t[133] & t[134] & ~t[135]) | (t[129] & ~t[131] & ~t[133] & t[135]) | (~t[129] & t[131] & t[133] & t[135]);
  assign t[101] = (t[130] & ~t[131] & ~t[132] & ~t[133] & ~t[134]) | (~t[129] & t[130] & ~t[132] & ~t[133] & ~t[135]) | (~t[129] & t[130] & ~t[131] & ~t[134] & ~t[135]) | (t[129] & ~t[130] & t[131] & t[132] & ~t[135]) | (t[129] & ~t[130] & t[133] & t[134] & ~t[135]) | (t[130] & ~t[132] & ~t[134] & t[135]) | (~t[130] & t[132] & t[134] & t[135]);
  assign t[102] = (t[129] & t[130] & t[131] & ~t[132] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[132] & ~t[133] & t[134] & t[135]) | (~t[130] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (~t[129] & ~t[131] & t[132] & ~t[134] & ~t[135]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[135]) | (~t[130] & t[131] & t[132] & t[133] & ~t[134]) | (~t[131] & t[132] & t[133] & ~t[135]);
  assign t[103] = (t[129] & t[130] & ~t[131] & ~t[133] & t[134] & ~t[135]) | (t[129] & t[131] & ~t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[131] & t[133] & ~t[134] & ~t[135]) | (~t[129] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[129] & ~t[130] & ~t[132] & t[133] & ~t[135]) | (~t[129] & ~t[131] & t[132] & t[133] & t[134]) | (t[132] & t[133] & ~t[134] & ~t[135]);
  assign t[104] = (t[129] & t[130] & ~t[132] & t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[129] & ~t[130] & ~t[131] & t[134] & ~t[135]) | (~t[130] & t[131] & ~t[132] & t[133] & t[134]) | (t[131] & ~t[133] & t[134] & ~t[135]);
  assign t[105] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[106] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[107] = (t[129] & t[130] & ~t[131] & t[132] & ~t[133] & ~t[135]) | (t[129] & ~t[131] & ~t[132] & t[133] & ~t[134] & t[135]) | (~t[130] & t[131] & ~t[132] & ~t[133] & ~t[135]) | (~t[129] & t[131] & ~t[132] & ~t[133] & ~t[134]) | (~t[129] & ~t[130] & t[131] & ~t[134] & ~t[135]) | (~t[129] & t[131] & t[132] & ~t[133] & t[134]) | (t[131] & ~t[132] & t[134] & ~t[135]);
  assign t[108] = t[136] ^ x[9];
  assign t[109] = t[137] ^ x[4];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[138] ^ x[5];
  assign t[111] = t[139] ^ x[6];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[7];
  assign t[114] = t[142] ^ x[8];
  assign t[115] = t[143] ^ x[19];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[49];
  assign t[118] = t[146] ^ x[21];
  assign t[119] = t[147] ^ x[22];
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = t[148] ^ x[23];
  assign t[121] = t[149] ^ x[18];
  assign t[122] = t[150] ^ x[29];
  assign t[123] = t[151] ^ x[30];
  assign t[124] = t[152] ^ x[50];
  assign t[125] = t[153] ^ x[31];
  assign t[126] = t[154] ^ x[32];
  assign t[127] = t[155] ^ x[33];
  assign t[128] = t[156] ^ x[28];
  assign t[129] = t[157] ^ x[39];
  assign t[12] = ~(t[17] & t[18]);
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[51];
  assign t[132] = t[160] ^ x[41];
  assign t[133] = t[161] ^ x[42];
  assign t[134] = t[162] ^ x[43];
  assign t[135] = t[163] ^ x[38];
  assign t[136] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[137] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[138] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[139] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[13] = ~(t[56] & t[19]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[143] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[144] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[145] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[146] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[147] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[148] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[149] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[14] = ~(t[57] & t[20]);
  assign t[150] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[151] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[152] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[153] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[154] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[155] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[156] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[157] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[158] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[159] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[15] = ~(t[58] & t[21]);
  assign t[160] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[161] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[162] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[163] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[59] & t[22]);
  assign t[17] = ~(t[60] & t[23]);
  assign t[18] = ~(t[61] & t[24]);
  assign t[19] = ~(t[62]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[62] & t[25]);
  assign t[21] = ~(t[63]);
  assign t[22] = ~(t[63] & t[26]);
  assign t[23] = ~(t[64]);
  assign t[24] = ~(t[64] & t[27]);
  assign t[25] = ~(t[56]);
  assign t[26] = ~(t[58]);
  assign t[27] = ~(t[60]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = ~t[31];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[4] ? x[45] : x[44];
  assign t[31] = ~(t[32] ^ t[33]);
  assign t[32] = t[34];
  assign t[33] = ~(t[35] ^ t[36]);
  assign t[34] = x[2] ? x[46] : t[37];
  assign t[35] = x[2] ? x[47] : t[38];
  assign t[36] = x[2] ? x[48] : t[39];
  assign t[37] = ~(t[40] & t[41]);
  assign t[38] = ~(t[42] & t[43]);
  assign t[39] = ~(t[44] & t[45]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[19] & t[46]);
  assign t[41] = ~(t[47] & t[65]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = ~(t[49] & t[66]);
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = ~(t[51] & t[67]);
  assign t[46] = ~(t[57]);
  assign t[47] = ~(t[52] & t[25]);
  assign t[48] = ~(t[59]);
  assign t[49] = ~(t[53] & t[26]);
  assign t[4] = ~x[2] & t[55];
  assign t[50] = ~(t[61]);
  assign t[51] = ~(t[54] & t[27]);
  assign t[52] = ~(t[57] & t[62]);
  assign t[53] = ~(t[59] & t[63]);
  assign t[54] = ~(t[61] & t[64]);
  assign t[55] = (t[68] & ~t[69]) | (~t[68] & t[69]);
  assign t[56] = (t[70] & ~t[72] & ~t[74]) | (~t[71] & t[72] & ~t[73]) | (~t[70] & ~t[72] & t[74]) | (t[71] & t[72] & t[73]);
  assign t[57] = (t[70] & ~t[73]) | (~t[70] & t[73]);
  assign t[58] = (t[75] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[75] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[59] = (t[75] & ~t[78]) | (~t[75] & t[78]);
  assign t[5] = t[7];
  assign t[60] = (t[80] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[80] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[61] = (t[80] & ~t[83]) | (~t[80] & t[83]);
  assign t[62] = (t[70] & ~t[72] & ~t[73]) | (~t[71] & t[72] & ~t[74]) | (~t[70] & ~t[72] & t[73]) | (t[71] & t[72] & t[74]);
  assign t[63] = (t[75] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[75] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[64] = (t[80] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[80] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[65] = (t[70] & ~t[85]) | (~t[70] & t[85]);
  assign t[66] = (t[75] & ~t[86]) | (~t[75] & t[86]);
  assign t[67] = (t[80] & ~t[87]) | (~t[80] & t[87]);
  assign t[68] = t[88] ^ x[9];
  assign t[69] = t[89] ^ x[10];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[19];
  assign t[71] = t[91] ^ x[20];
  assign t[72] = t[92] ^ x[21];
  assign t[73] = t[93] ^ x[22];
  assign t[74] = t[94] ^ x[23];
  assign t[75] = t[95] ^ x[29];
  assign t[76] = t[96] ^ x[30];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[32];
  assign t[79] = t[99] ^ x[33];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[39];
  assign t[81] = t[101] ^ x[40];
  assign t[82] = t[102] ^ x[41];
  assign t[83] = t[103] ^ x[42];
  assign t[84] = t[104] ^ x[43];
  assign t[85] = t[105] ^ x[49];
  assign t[86] = t[106] ^ x[50];
  assign t[87] = t[107] ^ x[51];
  assign t[88] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[89] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[91] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[92] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[93] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[94] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[95] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[96] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[97] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[98] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[99] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind173(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[101] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[102] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[103] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[104] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[105] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[106] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[9];
  assign t[108] = t[136] ^ x[4];
  assign t[109] = t[137] ^ x[5];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[138] ^ x[6];
  assign t[111] = t[139] ^ x[10];
  assign t[112] = t[140] ^ x[7];
  assign t[113] = t[141] ^ x[8];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[20];
  assign t[116] = t[144] ^ x[49];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[23];
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[30];
  assign t[123] = t[151] ^ x[50];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[33];
  assign t[127] = t[155] ^ x[28];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[40];
  assign t[12] = ~(t[17] & t[18]);
  assign t[130] = t[158] ^ x[51];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[43];
  assign t[134] = t[162] ^ x[38];
  assign t[135] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[136] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[137] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[138] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[55] & t[19]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[14] = ~(t[56] & t[20]);
  assign t[150] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[151] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[152] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[153] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[154] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[155] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[156] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[157] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[158] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[159] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[15] = ~(t[57] & t[21]);
  assign t[160] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[161] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[162] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[58] & t[22]);
  assign t[17] = ~(t[59] & t[23]);
  assign t[18] = ~(t[60] & t[24]);
  assign t[19] = ~(t[61]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[61] & t[25]);
  assign t[21] = ~(t[62]);
  assign t[22] = ~(t[62] & t[26]);
  assign t[23] = ~(t[63]);
  assign t[24] = ~(t[63] & t[27]);
  assign t[25] = ~(t[55]);
  assign t[26] = ~(t[57]);
  assign t[27] = ~(t[59]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = ~t[31];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[32] ? x[45] : x[44];
  assign t[31] = ~(t[33] ^ t[34]);
  assign t[32] = ~(t[35]);
  assign t[33] = t[36];
  assign t[34] = ~(t[37] ^ t[38]);
  assign t[35] = ~(t[4]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[19] & t[48]);
  assign t[43] = t[49] | t[64];
  assign t[44] = ~(t[21] & t[50]);
  assign t[45] = t[51] | t[65];
  assign t[46] = ~(t[23] & t[52]);
  assign t[47] = t[53] | t[66];
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[25] | t[19]);
  assign t[4] = ~x[2] & t[54];
  assign t[50] = ~(t[58]);
  assign t[51] = ~(t[26] | t[21]);
  assign t[52] = ~(t[60]);
  assign t[53] = ~(t[27] | t[23]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[69] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = (t[69] & ~t[72]) | (~t[69] & t[72]);
  assign t[57] = (t[74] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[74] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[58] = (t[74] & ~t[77]) | (~t[74] & t[77]);
  assign t[59] = (t[79] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[79] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[5] = t[7];
  assign t[60] = (t[79] & ~t[82]) | (~t[79] & t[82]);
  assign t[61] = (t[69] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[69] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[62] = (t[74] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[74] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[63] = (t[79] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[79] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[64] = (t[69] & ~t[84]) | (~t[69] & t[84]);
  assign t[65] = (t[74] & ~t[85]) | (~t[74] & t[85]);
  assign t[66] = (t[79] & ~t[86]) | (~t[79] & t[86]);
  assign t[67] = t[87] ^ x[9];
  assign t[68] = t[88] ^ x[10];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[21];
  assign t[72] = t[92] ^ x[22];
  assign t[73] = t[93] ^ x[23];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[31];
  assign t[77] = t[97] ^ x[32];
  assign t[78] = t[98] ^ x[33];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[49];
  assign t[85] = t[105] ^ x[50];
  assign t[86] = t[106] ^ x[51];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[91] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[92] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[93] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[94] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[95] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[96] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[97] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[98] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[99] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[28]) | (~t[0] & t[28]);
endmodule

module R2ind174(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[9];
  assign t[108] = t[136] ^ x[4];
  assign t[109] = t[137] ^ x[5];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[138] ^ x[6];
  assign t[111] = t[139] ^ x[10];
  assign t[112] = t[140] ^ x[7];
  assign t[113] = t[141] ^ x[8];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[17] & t[18]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[136] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[137] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[138] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[19] & t[20]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[21] & t[55]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[24] & t[56]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[57]);
  assign t[19] = ~(t[58]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[59]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[60]);
  assign t[23] = ~(t[61]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[62]);
  assign t[26] = ~(t[63]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[59] & t[58]);
  assign t[29] = ~(t[64]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[61] & t[60]);
  assign t[31] = ~(t[65]);
  assign t[32] = ~(t[63] & t[62]);
  assign t[33] = ~(t[66]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[38] ? x[48] : x[47];
  assign t[37] = ~(t[39] ^ t[40]);
  assign t[38] = ~(t[41]);
  assign t[39] = t[42];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[43] ^ t[44]);
  assign t[41] = ~(t[4]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[13] & t[48]);
  assign t[46] = ~(t[15] & t[49]);
  assign t[47] = ~(t[17] & t[50]);
  assign t[48] = t[51] | t[55];
  assign t[49] = t[52] | t[56];
  assign t[4] = ~x[2] & t[54];
  assign t[50] = t[53] | t[57];
  assign t[51] = ~(t[29] | t[19]);
  assign t[52] = ~(t[31] | t[22]);
  assign t[53] = ~(t[33] | t[25]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[59] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[5] = t[7];
  assign t[60] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[61] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[62] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[63] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[64] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[65] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[66] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[67] = t[87] ^ x[9];
  assign t[68] = t[88] ^ x[10];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[34]) | (~t[0] & t[34]);
endmodule

module R2ind175(x, y);
 input [56:0] x;
 output y;

 wire [189:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[33];
  assign t[101] = t[121] ^ x[34];
  assign t[102] = t[122] ^ x[35];
  assign t[103] = t[123] ^ x[36];
  assign t[104] = t[124] ^ x[37];
  assign t[105] = t[125] ^ x[38];
  assign t[106] = t[126] ^ x[39];
  assign t[107] = t[127] ^ x[40];
  assign t[108] = t[128] ^ x[41];
  assign t[109] = t[129] ^ x[42];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[130] ^ x[43];
  assign t[111] = t[131] ^ x[44];
  assign t[112] = t[132] ^ x[45];
  assign t[113] = t[133] ^ x[46];
  assign t[114] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[115] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[116] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[117] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[118] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[119] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[121] = (t[155] & t[156] & ~t[157] & t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[157] & ~t[158] & t[159] & ~t[160] & t[161]) | (~t[156] & t[157] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[156] & t[157] & ~t[160] & ~t[161]) | (~t[155] & t[157] & t[158] & ~t[159] & t[160]) | (t[157] & ~t[158] & t[160] & ~t[161]);
  assign t[122] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[123] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[124] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[125] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[126] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[127] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[128] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[129] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = (t[156] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & t[156] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[156] & ~t[157] & ~t[160] & ~t[161]) | (t[155] & ~t[156] & t[157] & t[158] & ~t[161]) | (t[155] & ~t[156] & t[159] & t[160] & ~t[161]) | (t[156] & ~t[158] & ~t[160] & t[161]) | (~t[156] & t[158] & t[160] & t[161]);
  assign t[131] = (t[155] & t[156] & t[157] & ~t[158] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & ~t[158] & ~t[159] & t[160] & t[161]) | (~t[156] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[157] & t[158] & ~t[160] & ~t[161]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[161]) | (~t[156] & t[157] & t[158] & t[159] & ~t[160]) | (~t[157] & t[158] & t[159] & ~t[161]);
  assign t[132] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[133] = (t[155] & t[156] & ~t[158] & t[159] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[158] & ~t[159] & t[160] & ~t[161]) | (~t[155] & ~t[156] & ~t[157] & t[160] & ~t[161]) | (~t[156] & t[157] & ~t[158] & t[159] & t[160]) | (t[157] & ~t[159] & t[160] & ~t[161]);
  assign t[134] = t[162] ^ x[9];
  assign t[135] = t[163] ^ x[4];
  assign t[136] = t[164] ^ x[5];
  assign t[137] = t[165] ^ x[6];
  assign t[138] = t[166] ^ x[10];
  assign t[139] = t[167] ^ x[7];
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = t[168] ^ x[8];
  assign t[141] = t[169] ^ x[19];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[20];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[18];
  assign t[148] = t[176] ^ x[26];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = ~(t[82] | t[21]);
  assign t[150] = t[178] ^ x[27];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[25];
  assign t[155] = t[183] ^ x[33];
  assign t[156] = t[184] ^ x[43];
  assign t[157] = t[185] ^ x[34];
  assign t[158] = t[186] ^ x[44];
  assign t[159] = t[187] ^ x[45];
  assign t[15] = ~(t[22] | t[23]);
  assign t[160] = t[188] ^ x[46];
  assign t[161] = t[189] ^ x[32];
  assign t[162] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[163] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[164] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[165] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[166] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[167] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[168] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[169] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[16] = ~(t[83] | t[24]);
  assign t[170] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[171] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[172] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[173] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[174] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[175] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[176] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[177] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[178] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[179] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[180] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[181] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[182] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[183] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[184] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[185] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[186] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[187] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[188] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[189] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[84] | t[27]);
  assign t[19] = ~(t[85]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[86]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[87]);
  assign t[23] = ~(t[88]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[89]);
  assign t[26] = ~(t[90]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[91]);
  assign t[29] = ~(t[85] | t[86]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[92]);
  assign t[31] = ~(t[87] | t[88]);
  assign t[32] = ~(t[93]);
  assign t[33] = ~(t[89] | t[90]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[38] ? x[48] : x[47];
  assign t[37] = ~(t[39] ^ t[40]);
  assign t[38] = ~(t[41]);
  assign t[39] = t[42];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[43] ^ t[44]);
  assign t[41] = ~(t[4]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[85] & t[20]);
  assign t[49] = ~(t[91] & t[54]);
  assign t[4] = ~x[2] & t[81];
  assign t[50] = ~(t[87] & t[23]);
  assign t[51] = ~(t[92] & t[55]);
  assign t[52] = ~(t[89] & t[26]);
  assign t[53] = ~(t[93] & t[56]);
  assign t[54] = ~(t[86] & t[19]);
  assign t[55] = ~(t[88] & t[22]);
  assign t[56] = ~(t[90] & t[25]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[38] ? x[53] : x[52];
  assign t[5] = t[7];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[20] & t[28]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = ~(t[75] & t[82]);
  assign t[71] = ~(t[23] & t[30]);
  assign t[72] = ~(t[76] & t[83]);
  assign t[73] = ~(t[26] & t[32]);
  assign t[74] = ~(t[77] & t[84]);
  assign t[75] = ~(t[78] & t[19]);
  assign t[76] = ~(t[79] & t[22]);
  assign t[77] = ~(t[80] & t[25]);
  assign t[78] = ~(t[91] & t[86]);
  assign t[79] = ~(t[92] & t[88]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = ~(t[93] & t[90]);
  assign t[81] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[82] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[83] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[84] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[85] = (t[96] & ~t[103] & ~t[105]) | (~t[102] & t[103] & ~t[104]) | (~t[96] & ~t[103] & t[105]) | (t[102] & t[103] & t[104]);
  assign t[86] = (t[96] & ~t[103] & ~t[104]) | (~t[102] & t[103] & ~t[105]) | (~t[96] & ~t[103] & t[104]) | (t[102] & t[103] & t[105]);
  assign t[87] = (t[98] & ~t[107] & ~t[109]) | (~t[106] & t[107] & ~t[108]) | (~t[98] & ~t[107] & t[109]) | (t[106] & t[107] & t[108]);
  assign t[88] = (t[98] & ~t[107] & ~t[108]) | (~t[106] & t[107] & ~t[109]) | (~t[98] & ~t[107] & t[108]) | (t[106] & t[107] & t[109]);
  assign t[89] = (t[100] & ~t[111] & ~t[113]) | (~t[110] & t[111] & ~t[112]) | (~t[100] & ~t[111] & t[113]) | (t[110] & t[111] & t[112]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = (t[100] & ~t[111] & ~t[112]) | (~t[110] & t[111] & ~t[113]) | (~t[100] & ~t[111] & t[112]) | (t[110] & t[111] & t[113]);
  assign t[91] = (t[96] & ~t[104]) | (~t[96] & t[104]);
  assign t[92] = (t[98] & ~t[108]) | (~t[98] & t[108]);
  assign t[93] = (t[100] & ~t[112]) | (~t[100] & t[112]);
  assign t[94] = t[114] ^ x[9];
  assign t[95] = t[115] ^ x[10];
  assign t[96] = t[116] ^ x[19];
  assign t[97] = t[117] ^ x[20];
  assign t[98] = t[118] ^ x[26];
  assign t[99] = t[119] ^ x[27];
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[34] & ~t[57]) | (~t[0] & t[34] & ~t[57]) | (~t[0] & ~t[34] & t[57]) | (t[0] & t[34] & t[57]);
endmodule

module R2ind176(x, y);
 input [56:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[39];
  assign t[101] = t[121] ^ x[40];
  assign t[102] = t[122] ^ x[41];
  assign t[103] = t[123] ^ x[42];
  assign t[104] = t[124] ^ x[43];
  assign t[105] = t[125] ^ x[44];
  assign t[106] = t[126] ^ x[45];
  assign t[107] = t[127] ^ x[46];
  assign t[108] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[109] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (t[135] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[136] & ~t[137] & ~t[140] & ~t[141]) | (~t[135] & t[136] & t[137] & t[138] & ~t[141]) | (~t[135] & t[136] & t[139] & t[140] & ~t[141]) | (t[135] & ~t[137] & ~t[139] & t[141]) | (~t[135] & t[137] & t[139] & t[141]);
  assign t[111] = (t[135] & t[136] & ~t[137] & t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[137] & ~t[138] & t[139] & ~t[140] & t[141]) | (~t[136] & t[137] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[136] & t[137] & ~t[140] & ~t[141]) | (~t[135] & t[137] & t[138] & ~t[139] & t[140]) | (t[137] & ~t[138] & t[140] & ~t[141]);
  assign t[112] = (t[142] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[143] & ~t[144] & ~t[147] & ~t[148]) | (~t[142] & t[143] & t[144] & t[145] & ~t[148]) | (~t[142] & t[143] & t[146] & t[147] & ~t[148]) | (t[142] & ~t[144] & ~t[146] & t[148]) | (~t[142] & t[144] & t[146] & t[148]);
  assign t[113] = (t[142] & t[143] & ~t[144] & t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[144] & ~t[145] & t[146] & ~t[147] & t[148]) | (~t[143] & t[144] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[143] & t[144] & ~t[147] & ~t[148]) | (~t[142] & t[144] & t[145] & ~t[146] & t[147]) | (t[144] & ~t[145] & t[147] & ~t[148]);
  assign t[114] = (t[149] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[150] & ~t[151] & ~t[154] & ~t[155]) | (~t[149] & t[150] & t[151] & t[152] & ~t[155]) | (~t[149] & t[150] & t[153] & t[154] & ~t[155]) | (t[149] & ~t[151] & ~t[153] & t[155]) | (~t[149] & t[151] & t[153] & t[155]);
  assign t[115] = (t[149] & t[150] & ~t[151] & t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[151] & ~t[152] & t[153] & ~t[154] & t[155]) | (~t[150] & t[151] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[150] & t[151] & ~t[154] & ~t[155]) | (~t[149] & t[151] & t[152] & ~t[153] & t[154]) | (t[151] & ~t[152] & t[154] & ~t[155]);
  assign t[116] = (t[136] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & t[136] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[136] & ~t[137] & ~t[140] & ~t[141]) | (t[135] & ~t[136] & t[137] & t[138] & ~t[141]) | (t[135] & ~t[136] & t[139] & t[140] & ~t[141]) | (t[136] & ~t[138] & ~t[140] & t[141]) | (~t[136] & t[138] & t[140] & t[141]);
  assign t[117] = (t[135] & t[136] & t[137] & ~t[138] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & ~t[138] & ~t[139] & t[140] & t[141]) | (~t[136] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[137] & t[138] & ~t[140] & ~t[141]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[141]) | (~t[136] & t[137] & t[138] & t[139] & ~t[140]) | (~t[137] & t[138] & t[139] & ~t[141]);
  assign t[118] = (t[135] & t[136] & ~t[137] & ~t[139] & t[140] & ~t[141]) | (t[135] & t[137] & ~t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & t[139] & ~t[140] & ~t[141]) | (~t[135] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[135] & ~t[136] & ~t[138] & t[139] & ~t[141]) | (~t[135] & ~t[137] & t[138] & t[139] & t[140]) | (t[138] & t[139] & ~t[140] & ~t[141]);
  assign t[119] = (t[135] & t[136] & ~t[138] & t[139] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[138] & ~t[139] & t[140] & ~t[141]) | (~t[135] & ~t[136] & ~t[137] & t[140] & ~t[141]) | (~t[136] & t[137] & ~t[138] & t[139] & t[140]) | (t[137] & ~t[139] & t[140] & ~t[141]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (t[143] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & t[143] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[143] & ~t[144] & ~t[147] & ~t[148]) | (t[142] & ~t[143] & t[144] & t[145] & ~t[148]) | (t[142] & ~t[143] & t[146] & t[147] & ~t[148]) | (t[143] & ~t[145] & ~t[147] & t[148]) | (~t[143] & t[145] & t[147] & t[148]);
  assign t[121] = (t[142] & t[143] & t[144] & ~t[145] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & ~t[145] & ~t[146] & t[147] & t[148]) | (~t[143] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[144] & t[145] & ~t[147] & ~t[148]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[148]) | (~t[143] & t[144] & t[145] & t[146] & ~t[147]) | (~t[144] & t[145] & t[146] & ~t[148]);
  assign t[122] = (t[142] & t[143] & ~t[144] & ~t[146] & t[147] & ~t[148]) | (t[142] & t[144] & ~t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & t[146] & ~t[147] & ~t[148]) | (~t[142] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[142] & ~t[143] & ~t[145] & t[146] & ~t[148]) | (~t[142] & ~t[144] & t[145] & t[146] & t[147]) | (t[145] & t[146] & ~t[147] & ~t[148]);
  assign t[123] = (t[142] & t[143] & ~t[145] & t[146] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[145] & ~t[146] & t[147] & ~t[148]) | (~t[142] & ~t[143] & ~t[144] & t[147] & ~t[148]) | (~t[143] & t[144] & ~t[145] & t[146] & t[147]) | (t[144] & ~t[146] & t[147] & ~t[148]);
  assign t[124] = (t[150] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & t[150] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[150] & ~t[151] & ~t[154] & ~t[155]) | (t[149] & ~t[150] & t[151] & t[152] & ~t[155]) | (t[149] & ~t[150] & t[153] & t[154] & ~t[155]) | (t[150] & ~t[152] & ~t[154] & t[155]) | (~t[150] & t[152] & t[154] & t[155]);
  assign t[125] = (t[149] & t[150] & t[151] & ~t[152] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & ~t[152] & ~t[153] & t[154] & t[155]) | (~t[150] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[151] & t[152] & ~t[154] & ~t[155]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[155]) | (~t[150] & t[151] & t[152] & t[153] & ~t[154]) | (~t[151] & t[152] & t[153] & ~t[155]);
  assign t[126] = (t[149] & t[150] & ~t[151] & ~t[153] & t[154] & ~t[155]) | (t[149] & t[151] & ~t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & t[153] & ~t[154] & ~t[155]) | (~t[149] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[149] & ~t[150] & ~t[152] & t[153] & ~t[155]) | (~t[149] & ~t[151] & t[152] & t[153] & t[154]) | (t[152] & t[153] & ~t[154] & ~t[155]);
  assign t[127] = (t[149] & t[150] & ~t[152] & t[153] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[152] & ~t[153] & t[154] & ~t[155]) | (~t[149] & ~t[150] & ~t[151] & t[154] & ~t[155]) | (~t[150] & t[151] & ~t[152] & t[153] & t[154]) | (t[151] & ~t[153] & t[154] & ~t[155]);
  assign t[128] = t[156] ^ x[9];
  assign t[129] = t[157] ^ x[4];
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = t[158] ^ x[5];
  assign t[131] = t[159] ^ x[6];
  assign t[132] = t[160] ^ x[10];
  assign t[133] = t[161] ^ x[7];
  assign t[134] = t[162] ^ x[8];
  assign t[135] = t[163] ^ x[19];
  assign t[136] = t[164] ^ x[35];
  assign t[137] = t[165] ^ x[20];
  assign t[138] = t[166] ^ x[36];
  assign t[139] = t[167] ^ x[37];
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = t[168] ^ x[38];
  assign t[141] = t[169] ^ x[18];
  assign t[142] = t[170] ^ x[26];
  assign t[143] = t[171] ^ x[39];
  assign t[144] = t[172] ^ x[27];
  assign t[145] = t[173] ^ x[40];
  assign t[146] = t[174] ^ x[41];
  assign t[147] = t[175] ^ x[42];
  assign t[148] = t[176] ^ x[25];
  assign t[149] = t[177] ^ x[33];
  assign t[14] = ~(t[76] | t[21]);
  assign t[150] = t[178] ^ x[43];
  assign t[151] = t[179] ^ x[34];
  assign t[152] = t[180] ^ x[44];
  assign t[153] = t[181] ^ x[45];
  assign t[154] = t[182] ^ x[46];
  assign t[155] = t[183] ^ x[32];
  assign t[156] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[157] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[158] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[159] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[15] = ~(t[22] | t[23]);
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[164] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[165] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[166] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[167] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[168] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[169] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[16] = ~(t[77] | t[24]);
  assign t[170] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[171] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[172] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[173] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[174] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[175] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[176] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[177] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[178] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[179] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[180] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[181] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[182] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[183] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[78] | t[27]);
  assign t[19] = ~(t[79]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[80]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[81]);
  assign t[23] = ~(t[82]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[83]);
  assign t[26] = ~(t[84]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[85]);
  assign t[29] = ~(t[79] | t[80]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[86]);
  assign t[31] = ~(t[81] | t[82]);
  assign t[32] = ~(t[87]);
  assign t[33] = ~(t[83] | t[84]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[38] ? x[48] : x[47];
  assign t[37] = ~(t[39] ^ t[40]);
  assign t[38] = ~(t[41]);
  assign t[39] = t[42];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[43] ^ t[44]);
  assign t[41] = ~(t[4]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[79] & t[20]);
  assign t[49] = ~(t[85] & t[54]);
  assign t[4] = ~x[2] & t[75];
  assign t[50] = ~(t[81] & t[23]);
  assign t[51] = ~(t[86] & t[55]);
  assign t[52] = ~(t[83] & t[26]);
  assign t[53] = ~(t[87] & t[56]);
  assign t[54] = ~(t[80] & t[19]);
  assign t[55] = ~(t[82] & t[22]);
  assign t[56] = ~(t[84] & t[25]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[4] ? x[53] : x[52];
  assign t[5] = t[7];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[20] & t[28]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[13] | t[76];
  assign t[71] = ~(t[23] & t[30]);
  assign t[72] = t[15] | t[77];
  assign t[73] = ~(t[26] & t[32]);
  assign t[74] = t[17] | t[78];
  assign t[75] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[76] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[77] = (t[92] & ~t[93]) | (~t[92] & t[93]);
  assign t[78] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[79] = (t[90] & ~t[97] & ~t[99]) | (~t[96] & t[97] & ~t[98]) | (~t[90] & ~t[97] & t[99]) | (t[96] & t[97] & t[98]);
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = (t[90] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[99]) | (~t[90] & ~t[97] & t[98]) | (t[96] & t[97] & t[99]);
  assign t[81] = (t[92] & ~t[101] & ~t[103]) | (~t[100] & t[101] & ~t[102]) | (~t[92] & ~t[101] & t[103]) | (t[100] & t[101] & t[102]);
  assign t[82] = (t[92] & ~t[101] & ~t[102]) | (~t[100] & t[101] & ~t[103]) | (~t[92] & ~t[101] & t[102]) | (t[100] & t[101] & t[103]);
  assign t[83] = (t[94] & ~t[105] & ~t[107]) | (~t[104] & t[105] & ~t[106]) | (~t[94] & ~t[105] & t[107]) | (t[104] & t[105] & t[106]);
  assign t[84] = (t[94] & ~t[105] & ~t[106]) | (~t[104] & t[105] & ~t[107]) | (~t[94] & ~t[105] & t[106]) | (t[104] & t[105] & t[107]);
  assign t[85] = (t[90] & ~t[98]) | (~t[90] & t[98]);
  assign t[86] = (t[92] & ~t[102]) | (~t[92] & t[102]);
  assign t[87] = (t[94] & ~t[106]) | (~t[94] & t[106]);
  assign t[88] = t[108] ^ x[9];
  assign t[89] = t[109] ^ x[10];
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = t[110] ^ x[19];
  assign t[91] = t[111] ^ x[20];
  assign t[92] = t[112] ^ x[26];
  assign t[93] = t[113] ^ x[27];
  assign t[94] = t[114] ^ x[33];
  assign t[95] = t[115] ^ x[34];
  assign t[96] = t[116] ^ x[35];
  assign t[97] = t[117] ^ x[36];
  assign t[98] = t[118] ^ x[37];
  assign t[99] = t[119] ^ x[38];
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[34] & ~t[57]) | (~t[0] & t[34] & ~t[57]) | (~t[0] & ~t[34] & t[57]) | (t[0] & t[34] & t[57]);
endmodule

module R2ind177(x, y);
 input [51:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[101] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[102] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[103] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[104] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[105] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[106] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[107] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[108] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[109] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[111] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[112] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[113] = t[141] ^ x[9];
  assign t[114] = t[142] ^ x[4];
  assign t[115] = t[143] ^ x[5];
  assign t[116] = t[144] ^ x[6];
  assign t[117] = t[145] ^ x[10];
  assign t[118] = t[146] ^ x[7];
  assign t[119] = t[147] ^ x[8];
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = t[148] ^ x[19];
  assign t[121] = t[149] ^ x[35];
  assign t[122] = t[150] ^ x[20];
  assign t[123] = t[151] ^ x[36];
  assign t[124] = t[152] ^ x[37];
  assign t[125] = t[153] ^ x[38];
  assign t[126] = t[154] ^ x[18];
  assign t[127] = t[155] ^ x[26];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[27];
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[25];
  assign t[134] = t[162] ^ x[33];
  assign t[135] = t[163] ^ x[43];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[44];
  assign t[138] = t[166] ^ x[45];
  assign t[139] = t[167] ^ x[46];
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = t[168] ^ x[32];
  assign t[141] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[142] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[143] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[144] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[149] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[14] = ~(t[61] | t[21]);
  assign t[150] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[151] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[152] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[153] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[154] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[155] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[156] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[157] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[158] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[159] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[15] = ~(t[22] | t[23]);
  assign t[160] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[161] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[162] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[163] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[164] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[165] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[166] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[167] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[168] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[62] | t[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[18] = ~(t[63] | t[27]);
  assign t[19] = ~(t[64]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[65]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[66]);
  assign t[23] = ~(t[67]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[68]);
  assign t[26] = ~(t[69]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[70]);
  assign t[29] = ~(t[64] | t[65]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[71]);
  assign t[31] = ~(t[66] | t[67]);
  assign t[32] = ~(t[72]);
  assign t[33] = ~(t[68] | t[69]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[38] ? x[48] : x[47];
  assign t[37] = ~(t[39] ^ t[40]);
  assign t[38] = ~(t[41]);
  assign t[39] = t[42];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[43] ^ t[44]);
  assign t[41] = ~(t[4]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[20] & t[28]);
  assign t[49] = ~(t[54] & t[61]);
  assign t[4] = ~x[2] & t[60];
  assign t[50] = ~(t[23] & t[30]);
  assign t[51] = ~(t[55] & t[62]);
  assign t[52] = ~(t[26] & t[32]);
  assign t[53] = ~(t[56] & t[63]);
  assign t[54] = ~(t[57] & t[19]);
  assign t[55] = ~(t[58] & t[22]);
  assign t[56] = ~(t[59] & t[25]);
  assign t[57] = ~(t[70] & t[65]);
  assign t[58] = ~(t[71] & t[67]);
  assign t[59] = ~(t[72] & t[69]);
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[61] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[62] = (t[77] & ~t[78]) | (~t[77] & t[78]);
  assign t[63] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[64] = (t[75] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[75] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[65] = (t[75] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[75] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[66] = (t[77] & ~t[86] & ~t[88]) | (~t[85] & t[86] & ~t[87]) | (~t[77] & ~t[86] & t[88]) | (t[85] & t[86] & t[87]);
  assign t[67] = (t[77] & ~t[86] & ~t[87]) | (~t[85] & t[86] & ~t[88]) | (~t[77] & ~t[86] & t[87]) | (t[85] & t[86] & t[88]);
  assign t[68] = (t[79] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[79] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[69] = (t[79] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[79] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[75] & ~t[83]) | (~t[75] & t[83]);
  assign t[71] = (t[77] & ~t[87]) | (~t[77] & t[87]);
  assign t[72] = (t[79] & ~t[91]) | (~t[79] & t[91]);
  assign t[73] = t[93] ^ x[9];
  assign t[74] = t[94] ^ x[10];
  assign t[75] = t[95] ^ x[19];
  assign t[76] = t[96] ^ x[20];
  assign t[77] = t[97] ^ x[26];
  assign t[78] = t[98] ^ x[27];
  assign t[79] = t[99] ^ x[33];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[34];
  assign t[81] = t[101] ^ x[35];
  assign t[82] = t[102] ^ x[36];
  assign t[83] = t[103] ^ x[37];
  assign t[84] = t[104] ^ x[38];
  assign t[85] = t[105] ^ x[39];
  assign t[86] = t[106] ^ x[40];
  assign t[87] = t[107] ^ x[41];
  assign t[88] = t[108] ^ x[42];
  assign t[89] = t[109] ^ x[43];
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = t[110] ^ x[44];
  assign t[91] = t[111] ^ x[45];
  assign t[92] = t[112] ^ x[46];
  assign t[93] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[97] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[98] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[99] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[34]) | (~t[0] & t[34]);
endmodule

module R2ind178(x, y);
 input [51:0] x;
 output y;

 wire [160:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[119] & t[120] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[119] & ~t[120] & ~t[121] & t[124] & ~t[125]) | (~t[120] & t[121] & ~t[122] & t[123] & t[124]) | (t[121] & ~t[123] & t[124] & ~t[125]);
  assign t[101] = (t[127] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (~t[126] & t[127] & ~t[129] & ~t[130] & ~t[132]) | (~t[126] & t[127] & ~t[128] & ~t[131] & ~t[132]) | (t[126] & ~t[127] & t[128] & t[129] & ~t[132]) | (t[126] & ~t[127] & t[130] & t[131] & ~t[132]) | (t[127] & ~t[129] & ~t[131] & t[132]) | (~t[127] & t[129] & t[131] & t[132]);
  assign t[102] = (t[126] & t[127] & t[128] & ~t[129] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[129] & ~t[130] & t[131] & t[132]) | (~t[127] & ~t[128] & t[129] & ~t[130] & ~t[131]) | (~t[126] & ~t[128] & t[129] & ~t[131] & ~t[132]) | (~t[126] & ~t[127] & t[129] & ~t[130] & ~t[132]) | (~t[127] & t[128] & t[129] & t[130] & ~t[131]) | (~t[128] & t[129] & t[130] & ~t[132]);
  assign t[103] = (t[126] & t[127] & ~t[128] & ~t[130] & t[131] & ~t[132]) | (t[126] & t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[132]) | (~t[126] & ~t[128] & ~t[129] & t[130] & ~t[131]) | (~t[126] & ~t[127] & ~t[129] & t[130] & ~t[132]) | (~t[126] & ~t[128] & t[129] & t[130] & t[131]) | (t[129] & t[130] & ~t[131] & ~t[132]);
  assign t[104] = (t[126] & t[127] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[126] & ~t[127] & ~t[128] & t[131] & ~t[132]) | (~t[127] & t[128] & ~t[129] & t[130] & t[131]) | (t[128] & ~t[130] & t[131] & ~t[132]);
  assign t[105] = t[133] ^ x[9];
  assign t[106] = t[134] ^ x[4];
  assign t[107] = t[135] ^ x[5];
  assign t[108] = t[136] ^ x[6];
  assign t[109] = t[137] ^ x[10];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[138] ^ x[7];
  assign t[111] = t[139] ^ x[8];
  assign t[112] = t[140] ^ x[19];
  assign t[113] = t[141] ^ x[35];
  assign t[114] = t[142] ^ x[20];
  assign t[115] = t[143] ^ x[36];
  assign t[116] = t[144] ^ x[37];
  assign t[117] = t[145] ^ x[38];
  assign t[118] = t[146] ^ x[18];
  assign t[119] = t[147] ^ x[26];
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = t[148] ^ x[39];
  assign t[121] = t[149] ^ x[27];
  assign t[122] = t[150] ^ x[40];
  assign t[123] = t[151] ^ x[41];
  assign t[124] = t[152] ^ x[42];
  assign t[125] = t[153] ^ x[25];
  assign t[126] = t[154] ^ x[33];
  assign t[127] = t[155] ^ x[43];
  assign t[128] = t[156] ^ x[34];
  assign t[129] = t[157] ^ x[44];
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = t[158] ^ x[45];
  assign t[131] = t[159] ^ x[46];
  assign t[132] = t[160] ^ x[32];
  assign t[133] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[134] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[135] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[136] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[137] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[138] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[141] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[142] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[143] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[144] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[145] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[146] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[147] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[148] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[149] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[14] = ~(t[53] | t[21]);
  assign t[150] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[151] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[152] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[153] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[154] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[155] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[156] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[157] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[158] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[159] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[15] = ~(t[22] | t[23]);
  assign t[160] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[54] | t[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[18] = ~(t[55] | t[27]);
  assign t[19] = ~(t[56]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[57]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[58]);
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[60]);
  assign t[26] = ~(t[61]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[62]);
  assign t[29] = ~(t[56] | t[57]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[63]);
  assign t[31] = ~(t[58] | t[59]);
  assign t[32] = ~(t[64]);
  assign t[33] = ~(t[60] | t[61]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[4] ? x[48] : x[47];
  assign t[37] = ~(t[38] ^ t[39]);
  assign t[38] = t[40];
  assign t[39] = ~(t[41] ^ t[42]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = x[2] ? x[49] : t[43];
  assign t[41] = x[2] ? x[50] : t[44];
  assign t[42] = x[2] ? x[51] : t[45];
  assign t[43] = ~(t[46] & t[47]);
  assign t[44] = ~(t[48] & t[49]);
  assign t[45] = ~(t[50] & t[51]);
  assign t[46] = ~(t[20] & t[28]);
  assign t[47] = t[13] | t[53];
  assign t[48] = ~(t[23] & t[30]);
  assign t[49] = t[15] | t[54];
  assign t[4] = ~x[2] & t[52];
  assign t[50] = ~(t[26] & t[32]);
  assign t[51] = t[17] | t[55];
  assign t[52] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[53] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[54] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[55] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[56] = (t[67] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[67] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[57] = (t[67] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[67] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[58] = (t[69] & ~t[78] & ~t[80]) | (~t[77] & t[78] & ~t[79]) | (~t[69] & ~t[78] & t[80]) | (t[77] & t[78] & t[79]);
  assign t[59] = (t[69] & ~t[78] & ~t[79]) | (~t[77] & t[78] & ~t[80]) | (~t[69] & ~t[78] & t[79]) | (t[77] & t[78] & t[80]);
  assign t[5] = t[7];
  assign t[60] = (t[71] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[71] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[61] = (t[71] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[71] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[62] = (t[67] & ~t[75]) | (~t[67] & t[75]);
  assign t[63] = (t[69] & ~t[79]) | (~t[69] & t[79]);
  assign t[64] = (t[71] & ~t[83]) | (~t[71] & t[83]);
  assign t[65] = t[85] ^ x[9];
  assign t[66] = t[86] ^ x[10];
  assign t[67] = t[87] ^ x[19];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[26];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[33];
  assign t[72] = t[92] ^ x[34];
  assign t[73] = t[93] ^ x[35];
  assign t[74] = t[94] ^ x[36];
  assign t[75] = t[95] ^ x[37];
  assign t[76] = t[96] ^ x[38];
  assign t[77] = t[97] ^ x[39];
  assign t[78] = t[98] ^ x[40];
  assign t[79] = t[99] ^ x[41];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[42];
  assign t[81] = t[101] ^ x[43];
  assign t[82] = t[102] ^ x[44];
  assign t[83] = t[103] ^ x[45];
  assign t[84] = t[104] ^ x[46];
  assign t[85] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[86] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[114] & ~t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[115] & ~t[116] & ~t[118]) | (t[112] & ~t[113] & ~t[114] & ~t[117] & ~t[118]) | (~t[112] & t[113] & t[114] & t[115] & ~t[118]) | (~t[112] & t[113] & t[116] & t[117] & ~t[118]) | (t[112] & ~t[114] & ~t[116] & t[118]) | (~t[112] & t[114] & t[116] & t[118]);
  assign t[88] = (t[112] & t[113] & ~t[114] & t[115] & ~t[116] & ~t[118]) | (t[112] & ~t[114] & ~t[115] & t[116] & ~t[117] & t[118]) | (~t[113] & t[114] & ~t[115] & ~t[116] & ~t[118]) | (~t[112] & t[114] & ~t[115] & ~t[116] & ~t[117]) | (~t[112] & ~t[113] & t[114] & ~t[117] & ~t[118]) | (~t[112] & t[114] & t[115] & ~t[116] & t[117]) | (t[114] & ~t[115] & t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[121] & ~t[122] & ~t[123] & ~t[124]) | (t[119] & ~t[120] & ~t[122] & ~t[123] & ~t[125]) | (t[119] & ~t[120] & ~t[121] & ~t[124] & ~t[125]) | (~t[119] & t[120] & t[121] & t[122] & ~t[125]) | (~t[119] & t[120] & t[123] & t[124] & ~t[125]) | (t[119] & ~t[121] & ~t[123] & t[125]) | (~t[119] & t[121] & t[123] & t[125]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = (t[119] & t[120] & ~t[121] & t[122] & ~t[123] & ~t[125]) | (t[119] & ~t[121] & ~t[122] & t[123] & ~t[124] & t[125]) | (~t[120] & t[121] & ~t[122] & ~t[123] & ~t[125]) | (~t[119] & t[121] & ~t[122] & ~t[123] & ~t[124]) | (~t[119] & ~t[120] & t[121] & ~t[124] & ~t[125]) | (~t[119] & t[121] & t[122] & ~t[123] & t[124]) | (t[121] & ~t[122] & t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & ~t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[127] & ~t[128] & ~t[131] & ~t[132]) | (~t[126] & t[127] & t[128] & t[129] & ~t[132]) | (~t[126] & t[127] & t[130] & t[131] & ~t[132]) | (t[126] & ~t[128] & ~t[130] & t[132]) | (~t[126] & t[128] & t[130] & t[132]);
  assign t[92] = (t[126] & t[127] & ~t[128] & t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[128] & ~t[129] & t[130] & ~t[131] & t[132]) | (~t[127] & t[128] & ~t[129] & ~t[130] & ~t[132]) | (~t[126] & t[128] & ~t[129] & ~t[130] & ~t[131]) | (~t[126] & ~t[127] & t[128] & ~t[131] & ~t[132]) | (~t[126] & t[128] & t[129] & ~t[130] & t[131]) | (t[128] & ~t[129] & t[131] & ~t[132]);
  assign t[93] = (t[113] & ~t[114] & ~t[115] & ~t[116] & ~t[117]) | (~t[112] & t[113] & ~t[115] & ~t[116] & ~t[118]) | (~t[112] & t[113] & ~t[114] & ~t[117] & ~t[118]) | (t[112] & ~t[113] & t[114] & t[115] & ~t[118]) | (t[112] & ~t[113] & t[116] & t[117] & ~t[118]) | (t[113] & ~t[115] & ~t[117] & t[118]) | (~t[113] & t[115] & t[117] & t[118]);
  assign t[94] = (t[112] & t[113] & t[114] & ~t[115] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[115] & ~t[116] & t[117] & t[118]) | (~t[113] & ~t[114] & t[115] & ~t[116] & ~t[117]) | (~t[112] & ~t[114] & t[115] & ~t[117] & ~t[118]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[118]) | (~t[113] & t[114] & t[115] & t[116] & ~t[117]) | (~t[114] & t[115] & t[116] & ~t[118]);
  assign t[95] = (t[112] & t[113] & ~t[114] & ~t[116] & t[117] & ~t[118]) | (t[112] & t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[118]) | (~t[112] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[112] & ~t[113] & ~t[115] & t[116] & ~t[118]) | (~t[112] & ~t[114] & t[115] & t[116] & t[117]) | (t[115] & t[116] & ~t[117] & ~t[118]);
  assign t[96] = (t[112] & t[113] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[112] & ~t[113] & ~t[114] & t[117] & ~t[118]) | (~t[113] & t[114] & ~t[115] & t[116] & t[117]) | (t[114] & ~t[116] & t[117] & ~t[118]);
  assign t[97] = (t[120] & ~t[121] & ~t[122] & ~t[123] & ~t[124]) | (~t[119] & t[120] & ~t[122] & ~t[123] & ~t[125]) | (~t[119] & t[120] & ~t[121] & ~t[124] & ~t[125]) | (t[119] & ~t[120] & t[121] & t[122] & ~t[125]) | (t[119] & ~t[120] & t[123] & t[124] & ~t[125]) | (t[120] & ~t[122] & ~t[124] & t[125]) | (~t[120] & t[122] & t[124] & t[125]);
  assign t[98] = (t[119] & t[120] & t[121] & ~t[122] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[122] & ~t[123] & t[124] & t[125]) | (~t[120] & ~t[121] & t[122] & ~t[123] & ~t[124]) | (~t[119] & ~t[121] & t[122] & ~t[124] & ~t[125]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[125]) | (~t[120] & t[121] & t[122] & t[123] & ~t[124]) | (~t[121] & t[122] & t[123] & ~t[125]);
  assign t[99] = (t[119] & t[120] & ~t[121] & ~t[123] & t[124] & ~t[125]) | (t[119] & t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[125]) | (~t[119] & ~t[121] & ~t[122] & t[123] & ~t[124]) | (~t[119] & ~t[120] & ~t[122] & t[123] & ~t[125]) | (~t[119] & ~t[121] & t[122] & t[123] & t[124]) | (t[122] & t[123] & ~t[124] & ~t[125]);
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[34]) | (~t[0] & t[34]);
endmodule

module R2ind179(x, y);
 input [51:0] x;
 output y;

 wire [165:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[101] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[102] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[103] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[104] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[105] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[106] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[107] = (t[117] & t[118] & ~t[119] & t[120] & ~t[121] & ~t[123]) | (t[117] & ~t[119] & ~t[120] & t[121] & ~t[122] & t[123]) | (~t[118] & t[119] & ~t[120] & ~t[121] & ~t[123]) | (~t[117] & t[119] & ~t[120] & ~t[121] & ~t[122]) | (~t[117] & ~t[118] & t[119] & ~t[122] & ~t[123]) | (~t[117] & t[119] & t[120] & ~t[121] & t[122]) | (t[119] & ~t[120] & t[122] & ~t[123]);
  assign t[108] = (t[124] & t[125] & ~t[126] & t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[126] & ~t[127] & t[128] & ~t[129] & t[130]) | (~t[125] & t[126] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[125] & t[126] & ~t[129] & ~t[130]) | (~t[124] & t[126] & t[127] & ~t[128] & t[129]) | (t[126] & ~t[127] & t[129] & ~t[130]);
  assign t[109] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[12];
  assign t[111] = t[139] ^ x[7];
  assign t[112] = t[140] ^ x[8];
  assign t[113] = t[141] ^ x[9];
  assign t[114] = t[142] ^ x[13];
  assign t[115] = t[143] ^ x[10];
  assign t[116] = t[144] ^ x[11];
  assign t[117] = t[145] ^ x[19];
  assign t[118] = t[146] ^ x[20];
  assign t[119] = t[147] ^ x[49];
  assign t[11] = ~x[2] & t[57];
  assign t[120] = t[148] ^ x[21];
  assign t[121] = t[149] ^ x[22];
  assign t[122] = t[150] ^ x[23];
  assign t[123] = t[151] ^ x[18];
  assign t[124] = t[152] ^ x[29];
  assign t[125] = t[153] ^ x[30];
  assign t[126] = t[154] ^ x[50];
  assign t[127] = t[155] ^ x[31];
  assign t[128] = t[156] ^ x[32];
  assign t[129] = t[157] ^ x[33];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[28];
  assign t[131] = t[159] ^ x[39];
  assign t[132] = t[160] ^ x[40];
  assign t[133] = t[161] ^ x[51];
  assign t[134] = t[162] ^ x[41];
  assign t[135] = t[163] ^ x[42];
  assign t[136] = t[164] ^ x[43];
  assign t[137] = t[165] ^ x[38];
  assign t[138] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[139] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[141] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[142] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[146] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[147] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[148] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[149] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[151] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[152] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[153] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[154] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[155] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[156] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[157] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[158] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[159] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[15] = ~(t[58] & t[21]);
  assign t[160] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[161] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[162] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[163] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[164] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[165] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[59] & t[22]);
  assign t[17] = ~(t[60] & t[23]);
  assign t[18] = ~(t[61] & t[24]);
  assign t[19] = ~(t[62] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[63] & t[26]);
  assign t[21] = ~(t[64]);
  assign t[22] = ~(t[64] & t[27]);
  assign t[23] = ~(t[65]);
  assign t[24] = ~(t[65] & t[28]);
  assign t[25] = ~(t[66]);
  assign t[26] = ~(t[66] & t[29]);
  assign t[27] = ~(t[58]);
  assign t[28] = ~(t[60]);
  assign t[29] = ~(t[62]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[4] ? x[45] : x[44];
  assign t[33] = ~(t[34] ^ t[35]);
  assign t[34] = t[36];
  assign t[35] = ~(t[37] ^ t[38]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = ~(t[49] & t[67]);
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = ~(t[51] & t[68]);
  assign t[46] = ~(t[25] & t[52]);
  assign t[47] = ~(t[53] & t[69]);
  assign t[48] = ~(t[59]);
  assign t[49] = ~(t[54] & t[27]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[61]);
  assign t[51] = ~(t[55] & t[28]);
  assign t[52] = ~(t[63]);
  assign t[53] = ~(t[56] & t[29]);
  assign t[54] = ~(t[59] & t[64]);
  assign t[55] = ~(t[61] & t[65]);
  assign t[56] = ~(t[63] & t[66]);
  assign t[57] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[58] = (t[72] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[72] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[59] = (t[72] & ~t[75]) | (~t[72] & t[75]);
  assign t[5] = t[8];
  assign t[60] = (t[77] & ~t[79] & ~t[81]) | (~t[78] & t[79] & ~t[80]) | (~t[77] & ~t[79] & t[81]) | (t[78] & t[79] & t[80]);
  assign t[61] = (t[77] & ~t[80]) | (~t[77] & t[80]);
  assign t[62] = (t[82] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[82] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[63] = (t[82] & ~t[85]) | (~t[82] & t[85]);
  assign t[64] = (t[72] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[72] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[65] = (t[77] & ~t[79] & ~t[80]) | (~t[78] & t[79] & ~t[81]) | (~t[77] & ~t[79] & t[80]) | (t[78] & t[79] & t[81]);
  assign t[66] = (t[82] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[82] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[67] = (t[72] & ~t[87]) | (~t[72] & t[87]);
  assign t[68] = (t[77] & ~t[88]) | (~t[77] & t[88]);
  assign t[69] = (t[82] & ~t[89]) | (~t[82] & t[89]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[12];
  assign t[71] = t[91] ^ x[13];
  assign t[72] = t[92] ^ x[19];
  assign t[73] = t[93] ^ x[20];
  assign t[74] = t[94] ^ x[21];
  assign t[75] = t[95] ^ x[22];
  assign t[76] = t[96] ^ x[23];
  assign t[77] = t[97] ^ x[29];
  assign t[78] = t[98] ^ x[30];
  assign t[79] = t[99] ^ x[31];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[32];
  assign t[81] = t[101] ^ x[33];
  assign t[82] = t[102] ^ x[39];
  assign t[83] = t[103] ^ x[40];
  assign t[84] = t[104] ^ x[41];
  assign t[85] = t[105] ^ x[42];
  assign t[86] = t[106] ^ x[43];
  assign t[87] = t[107] ^ x[49];
  assign t[88] = t[108] ^ x[50];
  assign t[89] = t[109] ^ x[51];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[110] & ~t[112] & ~t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[113] & ~t[114] & ~t[116]) | (t[110] & ~t[111] & ~t[112] & ~t[115] & ~t[116]) | (~t[110] & t[111] & t[112] & t[113] & ~t[116]) | (~t[110] & t[111] & t[114] & t[115] & ~t[116]) | (t[110] & ~t[112] & ~t[114] & t[116]) | (~t[110] & t[112] & t[114] & t[116]);
  assign t[91] = (t[110] & t[111] & ~t[112] & ~t[114] & t[115] & ~t[116]) | (t[110] & t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[116]) | (~t[110] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[110] & ~t[111] & ~t[113] & t[114] & ~t[116]) | (~t[110] & ~t[112] & t[113] & t[114] & t[115]) | (t[113] & t[114] & ~t[115] & ~t[116]);
  assign t[92] = (t[117] & ~t[119] & ~t[120] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & ~t[120] & ~t[121] & ~t[123]) | (t[117] & ~t[118] & ~t[119] & ~t[122] & ~t[123]) | (~t[117] & t[118] & t[119] & t[120] & ~t[123]) | (~t[117] & t[118] & t[121] & t[122] & ~t[123]) | (t[117] & ~t[119] & ~t[121] & t[123]) | (~t[117] & t[119] & t[121] & t[123]);
  assign t[93] = (t[118] & ~t[119] & ~t[120] & ~t[121] & ~t[122]) | (~t[117] & t[118] & ~t[120] & ~t[121] & ~t[123]) | (~t[117] & t[118] & ~t[119] & ~t[122] & ~t[123]) | (t[117] & ~t[118] & t[119] & t[120] & ~t[123]) | (t[117] & ~t[118] & t[121] & t[122] & ~t[123]) | (t[118] & ~t[120] & ~t[122] & t[123]) | (~t[118] & t[120] & t[122] & t[123]);
  assign t[94] = (t[117] & t[118] & t[119] & ~t[120] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[120] & ~t[121] & t[122] & t[123]) | (~t[118] & ~t[119] & t[120] & ~t[121] & ~t[122]) | (~t[117] & ~t[119] & t[120] & ~t[122] & ~t[123]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[123]) | (~t[118] & t[119] & t[120] & t[121] & ~t[122]) | (~t[119] & t[120] & t[121] & ~t[123]);
  assign t[95] = (t[117] & t[118] & ~t[119] & ~t[121] & t[122] & ~t[123]) | (t[117] & t[119] & ~t[120] & ~t[121] & ~t[122] & t[123]) | (~t[118] & ~t[119] & t[121] & ~t[122] & ~t[123]) | (~t[117] & ~t[119] & ~t[120] & t[121] & ~t[122]) | (~t[117] & ~t[118] & ~t[120] & t[121] & ~t[123]) | (~t[117] & ~t[119] & t[120] & t[121] & t[122]) | (t[120] & t[121] & ~t[122] & ~t[123]);
  assign t[96] = (t[117] & t[118] & ~t[120] & t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & t[120] & ~t[121] & ~t[122] & t[123]) | (~t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[117] & ~t[118] & ~t[119] & t[122] & ~t[123]) | (~t[118] & t[119] & ~t[120] & t[121] & t[122]) | (t[119] & ~t[121] & t[122] & ~t[123]);
  assign t[97] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[98] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[99] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[30]) | (~t[0] & t[30]);
endmodule

module R2ind180(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[101] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[102] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[103] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[104] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[105] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[106] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[20];
  assign t[116] = t[144] ^ x[49];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[23];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[30];
  assign t[123] = t[151] ^ x[50];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[33];
  assign t[127] = t[155] ^ x[28];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[40];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[51];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[43];
  assign t[134] = t[162] ^ x[38];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[151] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[152] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[153] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[154] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[155] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[156] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[157] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[158] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[159] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[15] = ~(t[55] & t[21]);
  assign t[160] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[161] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[162] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[56] & t[22]);
  assign t[17] = ~(t[57] & t[23]);
  assign t[18] = ~(t[58] & t[24]);
  assign t[19] = ~(t[59] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[60] & t[26]);
  assign t[21] = ~(t[61]);
  assign t[22] = ~(t[61] & t[27]);
  assign t[23] = ~(t[62]);
  assign t[24] = ~(t[62] & t[28]);
  assign t[25] = ~(t[63]);
  assign t[26] = ~(t[63] & t[29]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[59]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[11] ? x[45] : x[44];
  assign t[33] = ~(t[34] ^ t[35]);
  assign t[34] = t[36];
  assign t[35] = ~(t[37] ^ t[38]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = t[49] | t[64];
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = t[51] | t[65];
  assign t[46] = ~(t[25] & t[52]);
  assign t[47] = t[53] | t[66];
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[27] | t[21]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[58]);
  assign t[51] = ~(t[28] | t[23]);
  assign t[52] = ~(t[60]);
  assign t[53] = ~(t[29] | t[25]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[69] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = (t[69] & ~t[72]) | (~t[69] & t[72]);
  assign t[57] = (t[74] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[74] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[58] = (t[74] & ~t[77]) | (~t[74] & t[77]);
  assign t[59] = (t[79] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[79] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[5] = t[8];
  assign t[60] = (t[79] & ~t[82]) | (~t[79] & t[82]);
  assign t[61] = (t[69] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[69] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[62] = (t[74] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[74] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[63] = (t[79] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[79] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[64] = (t[69] & ~t[84]) | (~t[69] & t[84]);
  assign t[65] = (t[74] & ~t[85]) | (~t[74] & t[85]);
  assign t[66] = (t[79] & ~t[86]) | (~t[79] & t[86]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[21];
  assign t[72] = t[92] ^ x[22];
  assign t[73] = t[93] ^ x[23];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[31];
  assign t[77] = t[97] ^ x[32];
  assign t[78] = t[98] ^ x[33];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[49];
  assign t[85] = t[105] ^ x[50];
  assign t[86] = t[106] ^ x[51];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[91] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[92] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[93] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[94] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[95] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[96] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[97] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[98] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[99] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[30]) | (~t[0] & t[30]);
endmodule

module R2ind181(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[23] & t[55]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[56]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[57]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[61]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[62]);
  assign t[28] = ~(t[63]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[59] & t[58]);
  assign t[31] = ~(t[64]);
  assign t[32] = ~(t[61] & t[60]);
  assign t[33] = ~(t[65]);
  assign t[34] = ~(t[63] & t[62]);
  assign t[35] = ~(t[66]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[11] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[15] & t[48]);
  assign t[46] = ~(t[17] & t[49]);
  assign t[47] = ~(t[19] & t[50]);
  assign t[48] = t[51] | t[55];
  assign t[49] = t[52] | t[56];
  assign t[4] = ~(t[7]);
  assign t[50] = t[53] | t[57];
  assign t[51] = ~(t[31] | t[21]);
  assign t[52] = ~(t[33] | t[24]);
  assign t[53] = ~(t[35] | t[27]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[59] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[5] = t[8];
  assign t[60] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[61] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[62] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[63] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[64] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[65] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[66] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind182(x, y);
 input [56:0] x;
 output y;

 wire [189:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[33];
  assign t[101] = t[121] ^ x[34];
  assign t[102] = t[122] ^ x[35];
  assign t[103] = t[123] ^ x[36];
  assign t[104] = t[124] ^ x[37];
  assign t[105] = t[125] ^ x[38];
  assign t[106] = t[126] ^ x[39];
  assign t[107] = t[127] ^ x[40];
  assign t[108] = t[128] ^ x[41];
  assign t[109] = t[129] ^ x[42];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[130] ^ x[43];
  assign t[111] = t[131] ^ x[44];
  assign t[112] = t[132] ^ x[45];
  assign t[113] = t[133] ^ x[46];
  assign t[114] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[115] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[116] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[117] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[118] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[119] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[11] = ~x[2] & t[81];
  assign t[120] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[121] = (t[155] & t[156] & ~t[157] & t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[157] & ~t[158] & t[159] & ~t[160] & t[161]) | (~t[156] & t[157] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[156] & t[157] & ~t[160] & ~t[161]) | (~t[155] & t[157] & t[158] & ~t[159] & t[160]) | (t[157] & ~t[158] & t[160] & ~t[161]);
  assign t[122] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[123] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[124] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[125] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[126] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[127] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[128] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[129] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (t[156] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & t[156] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[156] & ~t[157] & ~t[160] & ~t[161]) | (t[155] & ~t[156] & t[157] & t[158] & ~t[161]) | (t[155] & ~t[156] & t[159] & t[160] & ~t[161]) | (t[156] & ~t[158] & ~t[160] & t[161]) | (~t[156] & t[158] & t[160] & t[161]);
  assign t[131] = (t[155] & t[156] & t[157] & ~t[158] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & ~t[158] & ~t[159] & t[160] & t[161]) | (~t[156] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[157] & t[158] & ~t[160] & ~t[161]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[161]) | (~t[156] & t[157] & t[158] & t[159] & ~t[160]) | (~t[157] & t[158] & t[159] & ~t[161]);
  assign t[132] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[133] = (t[155] & t[156] & ~t[158] & t[159] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[158] & ~t[159] & t[160] & ~t[161]) | (~t[155] & ~t[156] & ~t[157] & t[160] & ~t[161]) | (~t[156] & t[157] & ~t[158] & t[159] & t[160]) | (t[157] & ~t[159] & t[160] & ~t[161]);
  assign t[134] = t[162] ^ x[12];
  assign t[135] = t[163] ^ x[7];
  assign t[136] = t[164] ^ x[8];
  assign t[137] = t[165] ^ x[9];
  assign t[138] = t[166] ^ x[13];
  assign t[139] = t[167] ^ x[10];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[11];
  assign t[141] = t[169] ^ x[19];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[20];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[18];
  assign t[148] = t[176] ^ x[26];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[178] ^ x[27];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[25];
  assign t[155] = t[183] ^ x[33];
  assign t[156] = t[184] ^ x[43];
  assign t[157] = t[185] ^ x[34];
  assign t[158] = t[186] ^ x[44];
  assign t[159] = t[187] ^ x[45];
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = t[188] ^ x[46];
  assign t[161] = t[189] ^ x[32];
  assign t[162] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[163] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[164] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[165] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[166] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[167] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[168] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[169] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[16] = ~(t[82] | t[23]);
  assign t[170] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[171] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[172] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[173] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[174] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[175] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[176] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[177] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[178] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[179] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[180] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[181] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[182] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[183] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[184] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[185] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[186] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[187] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[188] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[189] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[83] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[84] | t[29]);
  assign t[21] = ~(t[85]);
  assign t[22] = ~(t[86]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[87]);
  assign t[25] = ~(t[88]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[89]);
  assign t[28] = ~(t[90]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[91]);
  assign t[31] = ~(t[85] | t[86]);
  assign t[32] = ~(t[92]);
  assign t[33] = ~(t[87] | t[88]);
  assign t[34] = ~(t[93]);
  assign t[35] = ~(t[89] | t[90]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[85] & t[22]);
  assign t[49] = ~(t[91] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[87] & t[25]);
  assign t[51] = ~(t[92] & t[55]);
  assign t[52] = ~(t[89] & t[28]);
  assign t[53] = ~(t[93] & t[56]);
  assign t[54] = ~(t[86] & t[21]);
  assign t[55] = ~(t[88] & t[24]);
  assign t[56] = ~(t[90] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[11] ? x[53] : x[52];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = ~(t[75] & t[82]);
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = ~(t[76] & t[83]);
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = ~(t[77] & t[84]);
  assign t[75] = ~(t[78] & t[21]);
  assign t[76] = ~(t[79] & t[24]);
  assign t[77] = ~(t[80] & t[27]);
  assign t[78] = ~(t[91] & t[86]);
  assign t[79] = ~(t[92] & t[88]);
  assign t[7] = ~(t[11]);
  assign t[80] = ~(t[93] & t[90]);
  assign t[81] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[82] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[83] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[84] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[85] = (t[96] & ~t[103] & ~t[105]) | (~t[102] & t[103] & ~t[104]) | (~t[96] & ~t[103] & t[105]) | (t[102] & t[103] & t[104]);
  assign t[86] = (t[96] & ~t[103] & ~t[104]) | (~t[102] & t[103] & ~t[105]) | (~t[96] & ~t[103] & t[104]) | (t[102] & t[103] & t[105]);
  assign t[87] = (t[98] & ~t[107] & ~t[109]) | (~t[106] & t[107] & ~t[108]) | (~t[98] & ~t[107] & t[109]) | (t[106] & t[107] & t[108]);
  assign t[88] = (t[98] & ~t[107] & ~t[108]) | (~t[106] & t[107] & ~t[109]) | (~t[98] & ~t[107] & t[108]) | (t[106] & t[107] & t[109]);
  assign t[89] = (t[100] & ~t[111] & ~t[113]) | (~t[110] & t[111] & ~t[112]) | (~t[100] & ~t[111] & t[113]) | (t[110] & t[111] & t[112]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[100] & ~t[111] & ~t[112]) | (~t[110] & t[111] & ~t[113]) | (~t[100] & ~t[111] & t[112]) | (t[110] & t[111] & t[113]);
  assign t[91] = (t[96] & ~t[104]) | (~t[96] & t[104]);
  assign t[92] = (t[98] & ~t[108]) | (~t[98] & t[108]);
  assign t[93] = (t[100] & ~t[112]) | (~t[100] & t[112]);
  assign t[94] = t[114] ^ x[12];
  assign t[95] = t[115] ^ x[13];
  assign t[96] = t[116] ^ x[19];
  assign t[97] = t[117] ^ x[20];
  assign t[98] = t[118] ^ x[26];
  assign t[99] = t[119] ^ x[27];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57]) | (~t[0] & t[36] & ~t[57]) | (~t[0] & ~t[36] & t[57]) | (t[0] & t[36] & t[57]);
endmodule

module R2ind183(x, y);
 input [56:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[120] ^ x[39];
  assign t[101] = t[121] ^ x[40];
  assign t[102] = t[122] ^ x[41];
  assign t[103] = t[123] ^ x[42];
  assign t[104] = t[124] ^ x[43];
  assign t[105] = t[125] ^ x[44];
  assign t[106] = t[126] ^ x[45];
  assign t[107] = t[127] ^ x[46];
  assign t[108] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[109] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (t[135] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[136] & ~t[137] & ~t[140] & ~t[141]) | (~t[135] & t[136] & t[137] & t[138] & ~t[141]) | (~t[135] & t[136] & t[139] & t[140] & ~t[141]) | (t[135] & ~t[137] & ~t[139] & t[141]) | (~t[135] & t[137] & t[139] & t[141]);
  assign t[111] = (t[135] & t[136] & ~t[137] & t[138] & ~t[139] & ~t[141]) | (t[135] & ~t[137] & ~t[138] & t[139] & ~t[140] & t[141]) | (~t[136] & t[137] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[136] & t[137] & ~t[140] & ~t[141]) | (~t[135] & t[137] & t[138] & ~t[139] & t[140]) | (t[137] & ~t[138] & t[140] & ~t[141]);
  assign t[112] = (t[142] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[143] & ~t[144] & ~t[147] & ~t[148]) | (~t[142] & t[143] & t[144] & t[145] & ~t[148]) | (~t[142] & t[143] & t[146] & t[147] & ~t[148]) | (t[142] & ~t[144] & ~t[146] & t[148]) | (~t[142] & t[144] & t[146] & t[148]);
  assign t[113] = (t[142] & t[143] & ~t[144] & t[145] & ~t[146] & ~t[148]) | (t[142] & ~t[144] & ~t[145] & t[146] & ~t[147] & t[148]) | (~t[143] & t[144] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[143] & t[144] & ~t[147] & ~t[148]) | (~t[142] & t[144] & t[145] & ~t[146] & t[147]) | (t[144] & ~t[145] & t[147] & ~t[148]);
  assign t[114] = (t[149] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[150] & ~t[151] & ~t[154] & ~t[155]) | (~t[149] & t[150] & t[151] & t[152] & ~t[155]) | (~t[149] & t[150] & t[153] & t[154] & ~t[155]) | (t[149] & ~t[151] & ~t[153] & t[155]) | (~t[149] & t[151] & t[153] & t[155]);
  assign t[115] = (t[149] & t[150] & ~t[151] & t[152] & ~t[153] & ~t[155]) | (t[149] & ~t[151] & ~t[152] & t[153] & ~t[154] & t[155]) | (~t[150] & t[151] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[150] & t[151] & ~t[154] & ~t[155]) | (~t[149] & t[151] & t[152] & ~t[153] & t[154]) | (t[151] & ~t[152] & t[154] & ~t[155]);
  assign t[116] = (t[136] & ~t[137] & ~t[138] & ~t[139] & ~t[140]) | (~t[135] & t[136] & ~t[138] & ~t[139] & ~t[141]) | (~t[135] & t[136] & ~t[137] & ~t[140] & ~t[141]) | (t[135] & ~t[136] & t[137] & t[138] & ~t[141]) | (t[135] & ~t[136] & t[139] & t[140] & ~t[141]) | (t[136] & ~t[138] & ~t[140] & t[141]) | (~t[136] & t[138] & t[140] & t[141]);
  assign t[117] = (t[135] & t[136] & t[137] & ~t[138] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & ~t[138] & ~t[139] & t[140] & t[141]) | (~t[136] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (~t[135] & ~t[137] & t[138] & ~t[140] & ~t[141]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[141]) | (~t[136] & t[137] & t[138] & t[139] & ~t[140]) | (~t[137] & t[138] & t[139] & ~t[141]);
  assign t[118] = (t[135] & t[136] & ~t[137] & ~t[139] & t[140] & ~t[141]) | (t[135] & t[137] & ~t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & t[139] & ~t[140] & ~t[141]) | (~t[135] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[135] & ~t[136] & ~t[138] & t[139] & ~t[141]) | (~t[135] & ~t[137] & t[138] & t[139] & t[140]) | (t[138] & t[139] & ~t[140] & ~t[141]);
  assign t[119] = (t[135] & t[136] & ~t[138] & t[139] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[138] & ~t[139] & t[140] & ~t[141]) | (~t[135] & ~t[136] & ~t[137] & t[140] & ~t[141]) | (~t[136] & t[137] & ~t[138] & t[139] & t[140]) | (t[137] & ~t[139] & t[140] & ~t[141]);
  assign t[11] = ~x[2] & t[75];
  assign t[120] = (t[143] & ~t[144] & ~t[145] & ~t[146] & ~t[147]) | (~t[142] & t[143] & ~t[145] & ~t[146] & ~t[148]) | (~t[142] & t[143] & ~t[144] & ~t[147] & ~t[148]) | (t[142] & ~t[143] & t[144] & t[145] & ~t[148]) | (t[142] & ~t[143] & t[146] & t[147] & ~t[148]) | (t[143] & ~t[145] & ~t[147] & t[148]) | (~t[143] & t[145] & t[147] & t[148]);
  assign t[121] = (t[142] & t[143] & t[144] & ~t[145] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & ~t[145] & ~t[146] & t[147] & t[148]) | (~t[143] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (~t[142] & ~t[144] & t[145] & ~t[147] & ~t[148]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[148]) | (~t[143] & t[144] & t[145] & t[146] & ~t[147]) | (~t[144] & t[145] & t[146] & ~t[148]);
  assign t[122] = (t[142] & t[143] & ~t[144] & ~t[146] & t[147] & ~t[148]) | (t[142] & t[144] & ~t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & t[146] & ~t[147] & ~t[148]) | (~t[142] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[142] & ~t[143] & ~t[145] & t[146] & ~t[148]) | (~t[142] & ~t[144] & t[145] & t[146] & t[147]) | (t[145] & t[146] & ~t[147] & ~t[148]);
  assign t[123] = (t[142] & t[143] & ~t[145] & t[146] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[145] & ~t[146] & t[147] & ~t[148]) | (~t[142] & ~t[143] & ~t[144] & t[147] & ~t[148]) | (~t[143] & t[144] & ~t[145] & t[146] & t[147]) | (t[144] & ~t[146] & t[147] & ~t[148]);
  assign t[124] = (t[150] & ~t[151] & ~t[152] & ~t[153] & ~t[154]) | (~t[149] & t[150] & ~t[152] & ~t[153] & ~t[155]) | (~t[149] & t[150] & ~t[151] & ~t[154] & ~t[155]) | (t[149] & ~t[150] & t[151] & t[152] & ~t[155]) | (t[149] & ~t[150] & t[153] & t[154] & ~t[155]) | (t[150] & ~t[152] & ~t[154] & t[155]) | (~t[150] & t[152] & t[154] & t[155]);
  assign t[125] = (t[149] & t[150] & t[151] & ~t[152] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & ~t[152] & ~t[153] & t[154] & t[155]) | (~t[150] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (~t[149] & ~t[151] & t[152] & ~t[154] & ~t[155]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[155]) | (~t[150] & t[151] & t[152] & t[153] & ~t[154]) | (~t[151] & t[152] & t[153] & ~t[155]);
  assign t[126] = (t[149] & t[150] & ~t[151] & ~t[153] & t[154] & ~t[155]) | (t[149] & t[151] & ~t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & t[153] & ~t[154] & ~t[155]) | (~t[149] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[149] & ~t[150] & ~t[152] & t[153] & ~t[155]) | (~t[149] & ~t[151] & t[152] & t[153] & t[154]) | (t[152] & t[153] & ~t[154] & ~t[155]);
  assign t[127] = (t[149] & t[150] & ~t[152] & t[153] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[152] & ~t[153] & t[154] & ~t[155]) | (~t[149] & ~t[150] & ~t[151] & t[154] & ~t[155]) | (~t[150] & t[151] & ~t[152] & t[153] & t[154]) | (t[151] & ~t[153] & t[154] & ~t[155]);
  assign t[128] = t[156] ^ x[12];
  assign t[129] = t[157] ^ x[7];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[8];
  assign t[131] = t[159] ^ x[9];
  assign t[132] = t[160] ^ x[13];
  assign t[133] = t[161] ^ x[10];
  assign t[134] = t[162] ^ x[11];
  assign t[135] = t[163] ^ x[19];
  assign t[136] = t[164] ^ x[35];
  assign t[137] = t[165] ^ x[20];
  assign t[138] = t[166] ^ x[36];
  assign t[139] = t[167] ^ x[37];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[38];
  assign t[141] = t[169] ^ x[18];
  assign t[142] = t[170] ^ x[26];
  assign t[143] = t[171] ^ x[39];
  assign t[144] = t[172] ^ x[27];
  assign t[145] = t[173] ^ x[40];
  assign t[146] = t[174] ^ x[41];
  assign t[147] = t[175] ^ x[42];
  assign t[148] = t[176] ^ x[25];
  assign t[149] = t[177] ^ x[33];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[178] ^ x[43];
  assign t[151] = t[179] ^ x[34];
  assign t[152] = t[180] ^ x[44];
  assign t[153] = t[181] ^ x[45];
  assign t[154] = t[182] ^ x[46];
  assign t[155] = t[183] ^ x[32];
  assign t[156] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[157] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[158] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[159] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[163] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[164] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[165] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[166] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[167] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[168] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[169] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[16] = ~(t[76] | t[23]);
  assign t[170] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[171] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[172] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[173] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[174] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[175] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[176] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[177] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[178] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[179] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[180] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[181] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[182] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[183] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[18] = ~(t[77] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[78] | t[29]);
  assign t[21] = ~(t[79]);
  assign t[22] = ~(t[80]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[81]);
  assign t[25] = ~(t[82]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[83]);
  assign t[28] = ~(t[84]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[85]);
  assign t[31] = ~(t[79] | t[80]);
  assign t[32] = ~(t[86]);
  assign t[33] = ~(t[81] | t[82]);
  assign t[34] = ~(t[87]);
  assign t[35] = ~(t[83] | t[84]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[79] & t[22]);
  assign t[49] = ~(t[85] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[81] & t[25]);
  assign t[51] = ~(t[86] & t[55]);
  assign t[52] = ~(t[83] & t[28]);
  assign t[53] = ~(t[87] & t[56]);
  assign t[54] = ~(t[80] & t[21]);
  assign t[55] = ~(t[82] & t[24]);
  assign t[56] = ~(t[84] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[4] ? x[53] : x[52];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[54] : t[66];
  assign t[64] = x[2] ? x[55] : t[67];
  assign t[65] = x[2] ? x[56] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[15] | t[76];
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = t[17] | t[77];
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = t[19] | t[78];
  assign t[75] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[76] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[77] = (t[92] & ~t[93]) | (~t[92] & t[93]);
  assign t[78] = (t[94] & ~t[95]) | (~t[94] & t[95]);
  assign t[79] = (t[90] & ~t[97] & ~t[99]) | (~t[96] & t[97] & ~t[98]) | (~t[90] & ~t[97] & t[99]) | (t[96] & t[97] & t[98]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[90] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[99]) | (~t[90] & ~t[97] & t[98]) | (t[96] & t[97] & t[99]);
  assign t[81] = (t[92] & ~t[101] & ~t[103]) | (~t[100] & t[101] & ~t[102]) | (~t[92] & ~t[101] & t[103]) | (t[100] & t[101] & t[102]);
  assign t[82] = (t[92] & ~t[101] & ~t[102]) | (~t[100] & t[101] & ~t[103]) | (~t[92] & ~t[101] & t[102]) | (t[100] & t[101] & t[103]);
  assign t[83] = (t[94] & ~t[105] & ~t[107]) | (~t[104] & t[105] & ~t[106]) | (~t[94] & ~t[105] & t[107]) | (t[104] & t[105] & t[106]);
  assign t[84] = (t[94] & ~t[105] & ~t[106]) | (~t[104] & t[105] & ~t[107]) | (~t[94] & ~t[105] & t[106]) | (t[104] & t[105] & t[107]);
  assign t[85] = (t[90] & ~t[98]) | (~t[90] & t[98]);
  assign t[86] = (t[92] & ~t[102]) | (~t[92] & t[102]);
  assign t[87] = (t[94] & ~t[106]) | (~t[94] & t[106]);
  assign t[88] = t[108] ^ x[12];
  assign t[89] = t[109] ^ x[13];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[110] ^ x[19];
  assign t[91] = t[111] ^ x[20];
  assign t[92] = t[112] ^ x[26];
  assign t[93] = t[113] ^ x[27];
  assign t[94] = t[114] ^ x[33];
  assign t[95] = t[115] ^ x[34];
  assign t[96] = t[116] ^ x[35];
  assign t[97] = t[117] ^ x[36];
  assign t[98] = t[118] ^ x[37];
  assign t[99] = t[119] ^ x[38];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57]) | (~t[0] & t[36] & ~t[57]) | (~t[0] & ~t[36] & t[57]) | (t[0] & t[36] & t[57]);
endmodule

module R2ind184(x, y);
 input [51:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[101] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[102] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[103] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[104] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[105] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[106] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[107] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[108] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[109] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[111] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[112] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[113] = t[141] ^ x[12];
  assign t[114] = t[142] ^ x[7];
  assign t[115] = t[143] ^ x[8];
  assign t[116] = t[144] ^ x[9];
  assign t[117] = t[145] ^ x[13];
  assign t[118] = t[146] ^ x[10];
  assign t[119] = t[147] ^ x[11];
  assign t[11] = ~x[2] & t[60];
  assign t[120] = t[148] ^ x[19];
  assign t[121] = t[149] ^ x[35];
  assign t[122] = t[150] ^ x[20];
  assign t[123] = t[151] ^ x[36];
  assign t[124] = t[152] ^ x[37];
  assign t[125] = t[153] ^ x[38];
  assign t[126] = t[154] ^ x[18];
  assign t[127] = t[155] ^ x[26];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[27];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[25];
  assign t[134] = t[162] ^ x[33];
  assign t[135] = t[163] ^ x[43];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[44];
  assign t[138] = t[166] ^ x[45];
  assign t[139] = t[167] ^ x[46];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[168] ^ x[32];
  assign t[141] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[142] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[143] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[144] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[149] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[151] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[152] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[153] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[154] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[155] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[156] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[157] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[158] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[159] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[161] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[162] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[163] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[164] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[165] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[166] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[167] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[168] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[61] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[62] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[63] | t[29]);
  assign t[21] = ~(t[64]);
  assign t[22] = ~(t[65]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[66]);
  assign t[25] = ~(t[67]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[69]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[70]);
  assign t[31] = ~(t[64] | t[65]);
  assign t[32] = ~(t[71]);
  assign t[33] = ~(t[66] | t[67]);
  assign t[34] = ~(t[72]);
  assign t[35] = ~(t[68] | t[69]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[11] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[22] & t[30]);
  assign t[49] = ~(t[54] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[25] & t[32]);
  assign t[51] = ~(t[55] & t[62]);
  assign t[52] = ~(t[28] & t[34]);
  assign t[53] = ~(t[56] & t[63]);
  assign t[54] = ~(t[57] & t[21]);
  assign t[55] = ~(t[58] & t[24]);
  assign t[56] = ~(t[59] & t[27]);
  assign t[57] = ~(t[70] & t[65]);
  assign t[58] = ~(t[71] & t[67]);
  assign t[59] = ~(t[72] & t[69]);
  assign t[5] = t[8];
  assign t[60] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[61] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[62] = (t[77] & ~t[78]) | (~t[77] & t[78]);
  assign t[63] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[64] = (t[75] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[75] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[65] = (t[75] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[75] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[66] = (t[77] & ~t[86] & ~t[88]) | (~t[85] & t[86] & ~t[87]) | (~t[77] & ~t[86] & t[88]) | (t[85] & t[86] & t[87]);
  assign t[67] = (t[77] & ~t[86] & ~t[87]) | (~t[85] & t[86] & ~t[88]) | (~t[77] & ~t[86] & t[87]) | (t[85] & t[86] & t[88]);
  assign t[68] = (t[79] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[79] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[69] = (t[79] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[79] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[75] & ~t[83]) | (~t[75] & t[83]);
  assign t[71] = (t[77] & ~t[87]) | (~t[77] & t[87]);
  assign t[72] = (t[79] & ~t[91]) | (~t[79] & t[91]);
  assign t[73] = t[93] ^ x[12];
  assign t[74] = t[94] ^ x[13];
  assign t[75] = t[95] ^ x[19];
  assign t[76] = t[96] ^ x[20];
  assign t[77] = t[97] ^ x[26];
  assign t[78] = t[98] ^ x[27];
  assign t[79] = t[99] ^ x[33];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[34];
  assign t[81] = t[101] ^ x[35];
  assign t[82] = t[102] ^ x[36];
  assign t[83] = t[103] ^ x[37];
  assign t[84] = t[104] ^ x[38];
  assign t[85] = t[105] ^ x[39];
  assign t[86] = t[106] ^ x[40];
  assign t[87] = t[107] ^ x[41];
  assign t[88] = t[108] ^ x[42];
  assign t[89] = t[109] ^ x[43];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[110] ^ x[44];
  assign t[91] = t[111] ^ x[45];
  assign t[92] = t[112] ^ x[46];
  assign t[93] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[97] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[98] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[99] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind185(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[55] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[56] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[57] | t[29]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[60]);
  assign t[25] = ~(t[61]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[62]);
  assign t[28] = ~(t[63]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[64]);
  assign t[31] = ~(t[58] | t[59]);
  assign t[32] = ~(t[65]);
  assign t[33] = ~(t[60] | t[61]);
  assign t[34] = ~(t[66]);
  assign t[35] = ~(t[62] | t[63]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[48] : x[47];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[22] & t[30]);
  assign t[49] = t[15] | t[55];
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[25] & t[32]);
  assign t[51] = t[17] | t[56];
  assign t[52] = ~(t[28] & t[34]);
  assign t[53] = t[19] | t[57];
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[59] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[5] = t[8];
  assign t[60] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[61] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[62] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[63] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[64] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[65] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[66] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36]) | (~t[0] & t[36]);
endmodule

module R2ind186(x, y);
 input [51:0] x;
 output y;

 wire [165:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[101] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[102] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[103] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[104] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[105] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[106] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[107] = (t[117] & t[118] & ~t[119] & t[120] & ~t[121] & ~t[123]) | (t[117] & ~t[119] & ~t[120] & t[121] & ~t[122] & t[123]) | (~t[118] & t[119] & ~t[120] & ~t[121] & ~t[123]) | (~t[117] & t[119] & ~t[120] & ~t[121] & ~t[122]) | (~t[117] & ~t[118] & t[119] & ~t[122] & ~t[123]) | (~t[117] & t[119] & t[120] & ~t[121] & t[122]) | (t[119] & ~t[120] & t[122] & ~t[123]);
  assign t[108] = (t[124] & t[125] & ~t[126] & t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[126] & ~t[127] & t[128] & ~t[129] & t[130]) | (~t[125] & t[126] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[125] & t[126] & ~t[129] & ~t[130]) | (~t[124] & t[126] & t[127] & ~t[128] & t[129]) | (t[126] & ~t[127] & t[129] & ~t[130]);
  assign t[109] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[12];
  assign t[111] = t[139] ^ x[7];
  assign t[112] = t[140] ^ x[8];
  assign t[113] = t[141] ^ x[9];
  assign t[114] = t[142] ^ x[13];
  assign t[115] = t[143] ^ x[10];
  assign t[116] = t[144] ^ x[11];
  assign t[117] = t[145] ^ x[19];
  assign t[118] = t[146] ^ x[20];
  assign t[119] = t[147] ^ x[49];
  assign t[11] = ~x[2] & t[57];
  assign t[120] = t[148] ^ x[21];
  assign t[121] = t[149] ^ x[22];
  assign t[122] = t[150] ^ x[23];
  assign t[123] = t[151] ^ x[18];
  assign t[124] = t[152] ^ x[29];
  assign t[125] = t[153] ^ x[30];
  assign t[126] = t[154] ^ x[50];
  assign t[127] = t[155] ^ x[31];
  assign t[128] = t[156] ^ x[32];
  assign t[129] = t[157] ^ x[33];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[28];
  assign t[131] = t[159] ^ x[39];
  assign t[132] = t[160] ^ x[40];
  assign t[133] = t[161] ^ x[51];
  assign t[134] = t[162] ^ x[41];
  assign t[135] = t[163] ^ x[42];
  assign t[136] = t[164] ^ x[43];
  assign t[137] = t[165] ^ x[38];
  assign t[138] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[139] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[141] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[142] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[146] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[147] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[148] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[149] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[151] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[152] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[153] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[154] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[155] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[156] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[157] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[158] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[159] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[15] = ~(t[58] & t[21]);
  assign t[160] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[161] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[162] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[163] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[164] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[165] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[59] & t[22]);
  assign t[17] = ~(t[60] & t[23]);
  assign t[18] = ~(t[61] & t[24]);
  assign t[19] = ~(t[62] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[63] & t[26]);
  assign t[21] = ~(t[64]);
  assign t[22] = ~(t[64] & t[27]);
  assign t[23] = ~(t[65]);
  assign t[24] = ~(t[65] & t[28]);
  assign t[25] = ~(t[66]);
  assign t[26] = ~(t[66] & t[29]);
  assign t[27] = ~(t[58]);
  assign t[28] = ~(t[60]);
  assign t[29] = ~(t[62]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[11] ? x[45] : x[44];
  assign t[33] = ~(t[34] ^ t[35]);
  assign t[34] = t[36];
  assign t[35] = ~(t[37] ^ t[38]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = ~(t[49] & t[67]);
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = ~(t[51] & t[68]);
  assign t[46] = ~(t[25] & t[52]);
  assign t[47] = ~(t[53] & t[69]);
  assign t[48] = ~(t[59]);
  assign t[49] = ~(t[54] & t[27]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[61]);
  assign t[51] = ~(t[55] & t[28]);
  assign t[52] = ~(t[63]);
  assign t[53] = ~(t[56] & t[29]);
  assign t[54] = ~(t[59] & t[64]);
  assign t[55] = ~(t[61] & t[65]);
  assign t[56] = ~(t[63] & t[66]);
  assign t[57] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[58] = (t[72] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[72] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[59] = (t[72] & ~t[75]) | (~t[72] & t[75]);
  assign t[5] = t[8];
  assign t[60] = (t[77] & ~t[79] & ~t[81]) | (~t[78] & t[79] & ~t[80]) | (~t[77] & ~t[79] & t[81]) | (t[78] & t[79] & t[80]);
  assign t[61] = (t[77] & ~t[80]) | (~t[77] & t[80]);
  assign t[62] = (t[82] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[82] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[63] = (t[82] & ~t[85]) | (~t[82] & t[85]);
  assign t[64] = (t[72] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[72] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[65] = (t[77] & ~t[79] & ~t[80]) | (~t[78] & t[79] & ~t[81]) | (~t[77] & ~t[79] & t[80]) | (t[78] & t[79] & t[81]);
  assign t[66] = (t[82] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[82] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[67] = (t[72] & ~t[87]) | (~t[72] & t[87]);
  assign t[68] = (t[77] & ~t[88]) | (~t[77] & t[88]);
  assign t[69] = (t[82] & ~t[89]) | (~t[82] & t[89]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[12];
  assign t[71] = t[91] ^ x[13];
  assign t[72] = t[92] ^ x[19];
  assign t[73] = t[93] ^ x[20];
  assign t[74] = t[94] ^ x[21];
  assign t[75] = t[95] ^ x[22];
  assign t[76] = t[96] ^ x[23];
  assign t[77] = t[97] ^ x[29];
  assign t[78] = t[98] ^ x[30];
  assign t[79] = t[99] ^ x[31];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[32];
  assign t[81] = t[101] ^ x[33];
  assign t[82] = t[102] ^ x[39];
  assign t[83] = t[103] ^ x[40];
  assign t[84] = t[104] ^ x[41];
  assign t[85] = t[105] ^ x[42];
  assign t[86] = t[106] ^ x[43];
  assign t[87] = t[107] ^ x[49];
  assign t[88] = t[108] ^ x[50];
  assign t[89] = t[109] ^ x[51];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[110] & ~t[112] & ~t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[113] & ~t[114] & ~t[116]) | (t[110] & ~t[111] & ~t[112] & ~t[115] & ~t[116]) | (~t[110] & t[111] & t[112] & t[113] & ~t[116]) | (~t[110] & t[111] & t[114] & t[115] & ~t[116]) | (t[110] & ~t[112] & ~t[114] & t[116]) | (~t[110] & t[112] & t[114] & t[116]);
  assign t[91] = (t[110] & t[111] & ~t[112] & ~t[114] & t[115] & ~t[116]) | (t[110] & t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[116]) | (~t[110] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[110] & ~t[111] & ~t[113] & t[114] & ~t[116]) | (~t[110] & ~t[112] & t[113] & t[114] & t[115]) | (t[113] & t[114] & ~t[115] & ~t[116]);
  assign t[92] = (t[117] & ~t[119] & ~t[120] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & ~t[120] & ~t[121] & ~t[123]) | (t[117] & ~t[118] & ~t[119] & ~t[122] & ~t[123]) | (~t[117] & t[118] & t[119] & t[120] & ~t[123]) | (~t[117] & t[118] & t[121] & t[122] & ~t[123]) | (t[117] & ~t[119] & ~t[121] & t[123]) | (~t[117] & t[119] & t[121] & t[123]);
  assign t[93] = (t[118] & ~t[119] & ~t[120] & ~t[121] & ~t[122]) | (~t[117] & t[118] & ~t[120] & ~t[121] & ~t[123]) | (~t[117] & t[118] & ~t[119] & ~t[122] & ~t[123]) | (t[117] & ~t[118] & t[119] & t[120] & ~t[123]) | (t[117] & ~t[118] & t[121] & t[122] & ~t[123]) | (t[118] & ~t[120] & ~t[122] & t[123]) | (~t[118] & t[120] & t[122] & t[123]);
  assign t[94] = (t[117] & t[118] & t[119] & ~t[120] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[120] & ~t[121] & t[122] & t[123]) | (~t[118] & ~t[119] & t[120] & ~t[121] & ~t[122]) | (~t[117] & ~t[119] & t[120] & ~t[122] & ~t[123]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[123]) | (~t[118] & t[119] & t[120] & t[121] & ~t[122]) | (~t[119] & t[120] & t[121] & ~t[123]);
  assign t[95] = (t[117] & t[118] & ~t[119] & ~t[121] & t[122] & ~t[123]) | (t[117] & t[119] & ~t[120] & ~t[121] & ~t[122] & t[123]) | (~t[118] & ~t[119] & t[121] & ~t[122] & ~t[123]) | (~t[117] & ~t[119] & ~t[120] & t[121] & ~t[122]) | (~t[117] & ~t[118] & ~t[120] & t[121] & ~t[123]) | (~t[117] & ~t[119] & t[120] & t[121] & t[122]) | (t[120] & t[121] & ~t[122] & ~t[123]);
  assign t[96] = (t[117] & t[118] & ~t[120] & t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & t[120] & ~t[121] & ~t[122] & t[123]) | (~t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[117] & ~t[118] & ~t[119] & t[122] & ~t[123]) | (~t[118] & t[119] & ~t[120] & t[121] & t[122]) | (t[119] & ~t[121] & t[122] & ~t[123]);
  assign t[97] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[98] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[99] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[30]) | (~t[0] & t[30]);
endmodule

module R2ind187(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[101] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[102] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[103] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[104] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[105] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[106] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[12];
  assign t[108] = t[136] ^ x[7];
  assign t[109] = t[137] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[138] ^ x[9];
  assign t[111] = t[139] ^ x[13];
  assign t[112] = t[140] ^ x[10];
  assign t[113] = t[141] ^ x[11];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[20];
  assign t[116] = t[144] ^ x[49];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[23];
  assign t[11] = ~x[2] & t[54];
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[30];
  assign t[123] = t[151] ^ x[50];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[33];
  assign t[127] = t[155] ^ x[28];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[40];
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = t[158] ^ x[51];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[43];
  assign t[134] = t[162] ^ x[38];
  assign t[135] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[136] = (x[6] & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0);
  assign t[137] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[138] = (x[6] & ~1'b0) | (~x[6] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[17] & t[18]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[151] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[152] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[153] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[154] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[155] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[156] = (x[34] & ~x[35] & ~x[36]) | (~x[34] & x[35] & ~x[36]) | (~x[34] & ~x[35] & x[36]) | (x[34] & x[35] & x[36]);
  assign t[157] = (x[34] & ~x[35] & ~x[37]) | (~x[34] & x[35] & ~x[37]) | (~x[34] & ~x[35] & x[37]) | (x[34] & x[35] & x[37]);
  assign t[158] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[159] = (x[34] & ~x[37]) | (~x[34] & x[37]);
  assign t[15] = ~(t[55] & t[21]);
  assign t[160] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[161] = (x[35] & ~x[37]) | (~x[35] & x[37]);
  assign t[162] = (x[36] & ~x[37]) | (~x[36] & x[37]);
  assign t[16] = ~(t[56] & t[22]);
  assign t[17] = ~(t[57] & t[23]);
  assign t[18] = ~(t[58] & t[24]);
  assign t[19] = ~(t[59] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[60] & t[26]);
  assign t[21] = ~(t[61]);
  assign t[22] = ~(t[61] & t[27]);
  assign t[23] = ~(t[62]);
  assign t[24] = ~(t[62] & t[28]);
  assign t[25] = ~(t[63]);
  assign t[26] = ~(t[63] & t[29]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[59]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[4] ? x[45] : x[44];
  assign t[33] = ~(t[34] ^ t[35]);
  assign t[34] = t[36];
  assign t[35] = ~(t[37] ^ t[38]);
  assign t[36] = x[2] ? x[46] : t[39];
  assign t[37] = x[2] ? x[47] : t[40];
  assign t[38] = x[2] ? x[48] : t[41];
  assign t[39] = ~(t[42] & t[43]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[44] & t[45]);
  assign t[41] = ~(t[46] & t[47]);
  assign t[42] = ~(t[21] & t[48]);
  assign t[43] = t[49] | t[64];
  assign t[44] = ~(t[23] & t[50]);
  assign t[45] = t[51] | t[65];
  assign t[46] = ~(t[25] & t[52]);
  assign t[47] = t[53] | t[66];
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[27] | t[21]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[58]);
  assign t[51] = ~(t[28] | t[23]);
  assign t[52] = ~(t[60]);
  assign t[53] = ~(t[29] | t[25]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[69] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = (t[69] & ~t[72]) | (~t[69] & t[72]);
  assign t[57] = (t[74] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[74] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[58] = (t[74] & ~t[77]) | (~t[74] & t[77]);
  assign t[59] = (t[79] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[79] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[5] = t[8];
  assign t[60] = (t[79] & ~t[82]) | (~t[79] & t[82]);
  assign t[61] = (t[69] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[69] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[62] = (t[74] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[74] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[63] = (t[79] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[79] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[64] = (t[69] & ~t[84]) | (~t[69] & t[84]);
  assign t[65] = (t[74] & ~t[85]) | (~t[74] & t[85]);
  assign t[66] = (t[79] & ~t[86]) | (~t[79] & t[86]);
  assign t[67] = t[87] ^ x[12];
  assign t[68] = t[88] ^ x[13];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[21];
  assign t[72] = t[92] ^ x[22];
  assign t[73] = t[93] ^ x[23];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[31];
  assign t[77] = t[97] ^ x[32];
  assign t[78] = t[98] ^ x[33];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = ~(t[11]);
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[49];
  assign t[85] = t[105] ^ x[50];
  assign t[86] = t[106] ^ x[51];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[91] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[92] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[93] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[94] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[95] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[96] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[97] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[98] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[99] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[30]) | (~t[0] & t[30]);
endmodule

module R2ind188(x, y);
 input [51:0] x;
 output y;

 wire [162:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[129] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & t[129] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[129] & ~t[130] & ~t[133] & ~t[134]) | (t[128] & ~t[129] & t[130] & t[131] & ~t[134]) | (t[128] & ~t[129] & t[132] & t[133] & ~t[134]) | (t[129] & ~t[131] & ~t[133] & t[134]) | (~t[129] & t[131] & t[133] & t[134]);
  assign t[104] = (t[128] & t[129] & t[130] & ~t[131] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[131] & ~t[132] & t[133] & t[134]) | (~t[129] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[130] & t[131] & ~t[133] & ~t[134]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[134]) | (~t[129] & t[130] & t[131] & t[132] & ~t[133]) | (~t[130] & t[131] & t[132] & ~t[134]);
  assign t[105] = (t[128] & t[129] & ~t[130] & ~t[132] & t[133] & ~t[134]) | (t[128] & t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[134]) | (~t[128] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[128] & ~t[129] & ~t[131] & t[132] & ~t[134]) | (~t[128] & ~t[130] & t[131] & t[132] & t[133]) | (t[131] & t[132] & ~t[133] & ~t[134]);
  assign t[106] = (t[128] & t[129] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[128] & ~t[129] & ~t[130] & t[133] & ~t[134]) | (~t[129] & t[130] & ~t[131] & t[132] & t[133]) | (t[130] & ~t[132] & t[133] & ~t[134]);
  assign t[107] = t[135] ^ x[9];
  assign t[108] = t[136] ^ x[4];
  assign t[109] = t[137] ^ x[5];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[138] ^ x[6];
  assign t[111] = t[139] ^ x[10];
  assign t[112] = t[140] ^ x[7];
  assign t[113] = t[141] ^ x[8];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[35];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[36];
  assign t[118] = t[146] ^ x[37];
  assign t[119] = t[147] ^ x[38];
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = t[148] ^ x[18];
  assign t[121] = t[149] ^ x[26];
  assign t[122] = t[150] ^ x[39];
  assign t[123] = t[151] ^ x[27];
  assign t[124] = t[152] ^ x[40];
  assign t[125] = t[153] ^ x[41];
  assign t[126] = t[154] ^ x[42];
  assign t[127] = t[155] ^ x[25];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = t[157] ^ x[43];
  assign t[12] = ~(t[17] & t[18]);
  assign t[130] = t[158] ^ x[34];
  assign t[131] = t[159] ^ x[44];
  assign t[132] = t[160] ^ x[45];
  assign t[133] = t[161] ^ x[46];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[136] = (x[3] & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0);
  assign t[137] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[138] = (x[3] & ~1'b0) | (~x[3] & 1'b0);
  assign t[139] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[13] = ~(t[19] & t[20]);
  assign t[140] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[141] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[142] = (x[14] & ~x[15] & ~x[16]) | (~x[14] & x[15] & ~x[16]) | (~x[14] & ~x[15] & x[16]) | (x[14] & x[15] & x[16]);
  assign t[143] = (x[14] & ~x[15] & ~x[17]) | (~x[14] & x[15] & ~x[17]) | (~x[14] & ~x[15] & x[17]) | (x[14] & x[15] & x[17]);
  assign t[144] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[145] = (x[14] & ~x[17]) | (~x[14] & x[17]);
  assign t[146] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[147] = (x[15] & ~x[17]) | (~x[15] & x[17]);
  assign t[148] = (x[16] & ~x[17]) | (~x[16] & x[17]);
  assign t[149] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[14] = ~(t[21] & t[55]);
  assign t[150] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[151] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[152] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[153] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[154] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[155] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[156] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[157] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[158] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[159] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[160] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[161] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[162] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[16] = ~(t[24] & t[56]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[57]);
  assign t[19] = ~(t[58]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[59]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[60]);
  assign t[23] = ~(t[61]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[62]);
  assign t[26] = ~(t[63]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[59] & t[58]);
  assign t[29] = ~(t[64]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[61] & t[60]);
  assign t[31] = ~(t[65]);
  assign t[32] = ~(t[63] & t[62]);
  assign t[33] = ~(t[66]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[38] ? x[48] : x[47];
  assign t[37] = ~(t[39] ^ t[40]);
  assign t[38] = ~(t[41]);
  assign t[39] = t[42];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[43] ^ t[44]);
  assign t[41] = ~(t[4]);
  assign t[42] = x[2] ? x[49] : t[45];
  assign t[43] = x[2] ? x[50] : t[46];
  assign t[44] = x[2] ? x[51] : t[47];
  assign t[45] = ~(t[13] & t[48]);
  assign t[46] = ~(t[15] & t[49]);
  assign t[47] = ~(t[17] & t[50]);
  assign t[48] = t[51] | t[55];
  assign t[49] = t[52] | t[56];
  assign t[4] = ~x[2] & t[54];
  assign t[50] = t[53] | t[57];
  assign t[51] = ~(t[29] | t[19]);
  assign t[52] = ~(t[31] | t[22]);
  assign t[53] = ~(t[33] | t[25]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[58] = (t[69] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[69] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[59] = (t[69] & ~t[77]) | (~t[69] & t[77]);
  assign t[5] = t[7];
  assign t[60] = (t[71] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[71] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[61] = (t[71] & ~t[81]) | (~t[71] & t[81]);
  assign t[62] = (t[73] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[73] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[63] = (t[73] & ~t[85]) | (~t[73] & t[85]);
  assign t[64] = (t[69] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[69] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[65] = (t[71] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[71] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[66] = (t[73] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[73] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[67] = t[87] ^ x[9];
  assign t[68] = t[88] ^ x[10];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[20];
  assign t[71] = t[91] ^ x[26];
  assign t[72] = t[92] ^ x[27];
  assign t[73] = t[93] ^ x[33];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[35];
  assign t[76] = t[96] ^ x[36];
  assign t[77] = t[97] ^ x[37];
  assign t[78] = t[98] ^ x[38];
  assign t[79] = t[99] ^ x[39];
  assign t[7] = x[2] ? x[11] : t[10];
  assign t[80] = t[100] ^ x[40];
  assign t[81] = t[101] ^ x[41];
  assign t[82] = t[102] ^ x[42];
  assign t[83] = t[103] ^ x[43];
  assign t[84] = t[104] ^ x[44];
  assign t[85] = t[105] ^ x[45];
  assign t[86] = t[106] ^ x[46];
  assign t[87] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[88] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[89] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[8] = x[2] ? x[12] : t[11];
  assign t[90] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[91] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[92] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[130] & ~t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[129] & ~t[130] & ~t[133] & ~t[134]) | (~t[128] & t[129] & t[130] & t[131] & ~t[134]) | (~t[128] & t[129] & t[132] & t[133] & ~t[134]) | (t[128] & ~t[130] & ~t[132] & t[134]) | (~t[128] & t[130] & t[132] & t[134]);
  assign t[94] = (t[128] & t[129] & ~t[130] & t[131] & ~t[132] & ~t[134]) | (t[128] & ~t[130] & ~t[131] & t[132] & ~t[133] & t[134]) | (~t[129] & t[130] & ~t[131] & ~t[132] & ~t[134]) | (~t[128] & t[130] & ~t[131] & ~t[132] & ~t[133]) | (~t[128] & ~t[129] & t[130] & ~t[133] & ~t[134]) | (~t[128] & t[130] & t[131] & ~t[132] & t[133]) | (t[130] & ~t[131] & t[133] & ~t[134]);
  assign t[95] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[96] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[97] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[98] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = x[2] ? x[13] : t[12];
  assign y = (t[0] & ~t[34]) | (~t[0] & t[34]);
endmodule

module R2_ind(x, y);
 input [448:0] x;
 output [188:0] y;

  R2ind0 R2ind0_inst(.x({x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[6], x[5], x[4], x[3], x[2], x[7], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[6], x[5], x[4], x[3], x[1], x[7], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[6], x[5], x[4], x[2], x[1], x[7], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[6], x[5], x[3], x[2], x[1], x[7], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[5], x[6], x[4], x[3], x[2], x[1], x[7], x[0]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[6], x[5], x[4], x[3], x[2], x[1], x[7], x[0]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.y(y[19]));
  R2ind20 R2ind20_inst(.y(y[20]));
  R2ind21 R2ind21_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[8]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[8]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[8]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[8]}), .y(y[24]));
  R2ind25 R2ind25_inst(.y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8]}), .y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.y(y[34]));
  R2ind35 R2ind35_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[8]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[8]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[8]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[8]}), .y(y[38]));
  R2ind39 R2ind39_inst(.y(y[39]));
  R2ind40 R2ind40_inst(.y(y[40]));
  R2ind41 R2ind41_inst(.y(y[41]));
  R2ind42 R2ind42_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[8]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[8]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[8]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[8]}), .y(y[45]));
  R2ind46 R2ind46_inst(.y(y[46]));
  R2ind47 R2ind47_inst(.y(y[47]));
  R2ind48 R2ind48_inst(.y(y[48]));
  R2ind49 R2ind49_inst(.x({x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[52]));
  R2ind53 R2ind53_inst(.y(y[53]));
  R2ind54 R2ind54_inst(.y(y[54]));
  R2ind55 R2ind55_inst(.y(y[55]));
  R2ind56 R2ind56_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8]}), .y(y[59]));
  R2ind60 R2ind60_inst(.y(y[60]));
  R2ind61 R2ind61_inst(.y(y[61]));
  R2ind62 R2ind62_inst(.y(y[62]));
  R2ind63 R2ind63_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8]}), .y(y[66]));
  R2ind67 R2ind67_inst(.y(y[67]));
  R2ind68 R2ind68_inst(.y(y[68]));
  R2ind69 R2ind69_inst(.y(y[69]));
  R2ind70 R2ind70_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[8]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[8]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[8]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[8]}), .y(y[73]));
  R2ind74 R2ind74_inst(.y(y[74]));
  R2ind75 R2ind75_inst(.y(y[75]));
  R2ind76 R2ind76_inst(.y(y[76]));
  R2ind77 R2ind77_inst(.x({x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[8], x[82], x[81]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[103], x[102], x[101], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[8], x[82], x[81]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[100], x[99], x[98], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[8], x[82], x[81]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[103], x[102], x[101], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[8], x[82], x[81]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[90], x[100], x[99], x[98], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[94], x[93], x[92], x[91], x[89], x[88], x[87], x[86], x[85], x[84], x[97], x[8], x[96], x[95]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[90], x[103], x[102], x[101], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[94], x[93], x[92], x[91], x[89], x[88], x[87], x[86], x[85], x[84], x[97], x[8], x[96], x[95]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[103], x[102], x[101], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[100], x[8], x[99], x[98]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[8], x[105], x[104]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[126], x[125], x[124], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[8], x[105], x[104]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[123], x[122], x[121], x[117], x[116], x[115], x[114], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[8], x[105], x[104]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[126], x[125], x[124], x[117], x[116], x[115], x[114], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[8], x[105], x[104]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[113], x[123], x[122], x[121], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[117], x[116], x[115], x[114], x[112], x[111], x[110], x[109], x[108], x[107], x[120], x[8], x[119], x[118]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[113], x[126], x[125], x[124], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[117], x[116], x[115], x[114], x[112], x[111], x[110], x[109], x[108], x[107], x[120], x[8], x[119], x[118]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[126], x[125], x[124], x[117], x[116], x[115], x[114], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[123], x[8], x[122], x[121]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[8], x[128], x[127]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[149], x[148], x[147], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[8], x[128], x[127]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[146], x[145], x[144], x[140], x[139], x[138], x[137], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[8], x[128], x[127]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[149], x[148], x[147], x[140], x[139], x[138], x[137], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[8], x[128], x[127]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[136], x[146], x[145], x[144], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[140], x[139], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[143], x[8], x[142], x[141]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[136], x[149], x[148], x[147], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[140], x[139], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[143], x[8], x[142], x[141]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[149], x[148], x[147], x[140], x[139], x[138], x[137], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[146], x[8], x[145], x[144]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[8], x[151], x[150]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[172], x[171], x[170], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[8], x[151], x[150]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[169], x[168], x[167], x[163], x[162], x[161], x[160], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[8], x[151], x[150]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[172], x[171], x[170], x[163], x[162], x[161], x[160], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[8], x[151], x[150]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[159], x[169], x[168], x[167], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[163], x[162], x[161], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[166], x[8], x[165], x[164]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[159], x[172], x[171], x[170], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[163], x[162], x[161], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[166], x[8], x[165], x[164]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[172], x[171], x[170], x[163], x[162], x[161], x[160], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[169], x[8], x[168], x[167]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[8], x[174], x[173]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[195], x[194], x[193], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[8], x[174], x[173]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[192], x[191], x[190], x[186], x[185], x[184], x[183], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[8], x[174], x[173]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[195], x[194], x[193], x[186], x[185], x[184], x[183], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[8], x[174], x[173]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[182], x[192], x[191], x[190], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[189], x[8], x[188], x[187]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[182], x[195], x[194], x[193], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[189], x[8], x[188], x[187]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[195], x[194], x[193], x[186], x[185], x[184], x[183], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[192], x[8], x[191], x[190]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[8], x[197], x[196]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[218], x[217], x[216], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[8], x[197], x[196]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[215], x[214], x[213], x[209], x[208], x[207], x[206], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[8], x[197], x[196]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[218], x[217], x[216], x[209], x[208], x[207], x[206], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[8], x[197], x[196]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[205], x[215], x[214], x[213], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[209], x[208], x[207], x[206], x[204], x[203], x[202], x[201], x[200], x[199], x[212], x[8], x[211], x[210]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[205], x[218], x[217], x[216], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[209], x[208], x[207], x[206], x[204], x[203], x[202], x[201], x[200], x[199], x[212], x[8], x[211], x[210]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[218], x[217], x[216], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[215], x[8], x[214], x[213]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[221], x[8], x[220], x[219]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[241], x[240], x[239], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[221], x[8], x[220], x[219]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[238], x[237], x[236], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[221], x[8], x[220], x[219]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[241], x[240], x[239], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[221], x[8], x[220], x[219]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[228], x[238], x[237], x[236], x[232], x[231], x[230], x[229], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[235], x[8], x[234], x[233]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[228], x[241], x[240], x[239], x[232], x[231], x[230], x[229], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[235], x[8], x[234], x[233]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[241], x[240], x[239], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[238], x[8], x[237], x[236]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[261], x[260], x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[8], x[243], x[242]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[264], x[263], x[262], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[8], x[243], x[242]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[261], x[260], x[259], x[255], x[254], x[253], x[252], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[8], x[243], x[242]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[264], x[263], x[262], x[255], x[254], x[253], x[252], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[8], x[243], x[242]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[251], x[261], x[260], x[259], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[255], x[254], x[253], x[252], x[250], x[249], x[248], x[247], x[246], x[245], x[258], x[8], x[257], x[256]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[251], x[264], x[263], x[262], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[255], x[254], x[253], x[252], x[250], x[249], x[248], x[247], x[246], x[245], x[258], x[8], x[257], x[256]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[264], x[263], x[262], x[255], x[254], x[253], x[252], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[261], x[8], x[260], x[259]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[284], x[100], x[283], x[282], x[281], x[97], x[280], x[279], x[278], x[277], x[276], x[275], x[94], x[93], x[92], x[91], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[267], x[83], x[8], x[266], x[265]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[287], x[103], x[286], x[285], x[281], x[97], x[280], x[279], x[278], x[277], x[276], x[275], x[94], x[93], x[92], x[91], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[267], x[83], x[8], x[266], x[265]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[284], x[100], x[283], x[282], x[278], x[277], x[276], x[275], x[94], x[93], x[92], x[91], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[267], x[83], x[8], x[266], x[265]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[287], x[103], x[286], x[285], x[278], x[277], x[276], x[275], x[94], x[93], x[92], x[91], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[267], x[83], x[8], x[266], x[265]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[274], x[90], x[284], x[100], x[283], x[282], x[278], x[277], x[276], x[275], x[273], x[272], x[271], x[270], x[269], x[268], x[94], x[93], x[92], x[91], x[89], x[88], x[87], x[86], x[85], x[84], x[281], x[97], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[280], x[279]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[274], x[90], x[287], x[103], x[286], x[285], x[278], x[277], x[276], x[275], x[273], x[272], x[271], x[270], x[269], x[268], x[94], x[93], x[92], x[91], x[89], x[88], x[87], x[86], x[85], x[84], x[281], x[97], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[280], x[279]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[287], x[103], x[286], x[285], x[278], x[277], x[276], x[275], x[94], x[93], x[92], x[91], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[284], x[100], x[8], x[283], x[282]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[307], x[123], x[306], x[305], x[304], x[120], x[303], x[302], x[301], x[300], x[299], x[298], x[117], x[116], x[115], x[114], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[290], x[106], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[289], x[288]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[310], x[126], x[309], x[308], x[304], x[120], x[303], x[302], x[301], x[300], x[299], x[298], x[117], x[116], x[115], x[114], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[290], x[106], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[289], x[288]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[307], x[123], x[306], x[305], x[301], x[300], x[299], x[298], x[117], x[116], x[115], x[114], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[290], x[106], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[289], x[288]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[310], x[126], x[309], x[308], x[301], x[300], x[299], x[298], x[117], x[116], x[115], x[114], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[290], x[106], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[289], x[288]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[297], x[113], x[307], x[123], x[306], x[305], x[301], x[300], x[299], x[298], x[296], x[295], x[294], x[293], x[292], x[291], x[117], x[116], x[115], x[114], x[112], x[111], x[110], x[109], x[108], x[107], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[304], x[120], x[8], x[303], x[302]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[297], x[113], x[310], x[126], x[309], x[308], x[301], x[300], x[299], x[298], x[296], x[295], x[294], x[293], x[292], x[291], x[117], x[116], x[115], x[114], x[112], x[111], x[110], x[109], x[108], x[107], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[304], x[120], x[8], x[303], x[302]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[310], x[126], x[309], x[308], x[301], x[300], x[299], x[298], x[117], x[116], x[115], x[114], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[307], x[123], x[8], x[306], x[305]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[330], x[146], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[329], x[328], x[327], x[143], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[326], x[325], x[324], x[323], x[322], x[321], x[140], x[139], x[138], x[137], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[313], x[129], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[8], x[312], x[311]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[333], x[149], x[332], x[331], x[327], x[143], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[326], x[325], x[324], x[323], x[322], x[321], x[140], x[139], x[138], x[137], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[313], x[129], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[8], x[312], x[311]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[330], x[146], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[329], x[328], x[324], x[323], x[322], x[321], x[140], x[139], x[138], x[137], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[313], x[129], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[8], x[312], x[311]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[333], x[149], x[332], x[331], x[324], x[323], x[322], x[321], x[140], x[139], x[138], x[137], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[313], x[129], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[8], x[312], x[311]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[320], x[136], x[330], x[146], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[329], x[328], x[324], x[323], x[322], x[321], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[140], x[139], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[327], x[143], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8], x[326], x[325]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[320], x[136], x[333], x[149], x[332], x[331], x[324], x[323], x[322], x[321], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[140], x[139], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[327], x[143], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[8], x[326], x[325]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[333], x[149], x[332], x[331], x[324], x[323], x[322], x[321], x[140], x[139], x[138], x[137], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[330], x[146], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[8], x[329], x[328]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[353], x[169], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[352], x[351], x[350], x[166], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[349], x[348], x[347], x[346], x[345], x[344], x[163], x[162], x[161], x[160], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[336], x[152], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8], x[335], x[334]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[356], x[172], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[355], x[354], x[350], x[166], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[349], x[348], x[347], x[346], x[345], x[344], x[163], x[162], x[161], x[160], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[336], x[152], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8], x[335], x[334]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[353], x[169], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[352], x[351], x[347], x[346], x[345], x[344], x[163], x[162], x[161], x[160], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[336], x[152], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8], x[335], x[334]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[356], x[172], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[355], x[354], x[347], x[346], x[345], x[344], x[163], x[162], x[161], x[160], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[336], x[152], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[8], x[335], x[334]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[343], x[159], x[353], x[169], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[352], x[351], x[347], x[346], x[345], x[344], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[163], x[162], x[161], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[350], x[166], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[8], x[349], x[348]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[343], x[159], x[356], x[172], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[355], x[354], x[347], x[346], x[345], x[344], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[163], x[162], x[161], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[350], x[166], x[56], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[8], x[349], x[348]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[356], x[172], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[355], x[354], x[347], x[346], x[345], x[344], x[163], x[162], x[161], x[160], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[353], x[169], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[8], x[352], x[351]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[100], x[192], x[376], x[375], x[374], x[97], x[189], x[373], x[372], x[371], x[94], x[93], x[92], x[91], x[186], x[185], x[184], x[183], x[370], x[369], x[368], x[367], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[175], x[359], x[8], x[358], x[357]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[103], x[195], x[379], x[378], x[377], x[97], x[189], x[373], x[372], x[371], x[94], x[93], x[92], x[91], x[186], x[185], x[184], x[183], x[370], x[369], x[368], x[367], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[175], x[359], x[8], x[358], x[357]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[100], x[192], x[376], x[375], x[374], x[94], x[93], x[92], x[91], x[186], x[185], x[184], x[183], x[370], x[369], x[368], x[367], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[175], x[359], x[8], x[358], x[357]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[103], x[195], x[379], x[378], x[377], x[94], x[93], x[92], x[91], x[186], x[185], x[184], x[183], x[370], x[369], x[368], x[367], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[83], x[175], x[359], x[8], x[358], x[357]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[90], x[182], x[366], x[100], x[192], x[376], x[375], x[374], x[94], x[93], x[92], x[91], x[89], x[88], x[87], x[86], x[85], x[84], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[370], x[369], x[368], x[367], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[97], x[189], x[373], x[8], x[372], x[371]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[90], x[182], x[366], x[103], x[195], x[379], x[378], x[377], x[94], x[93], x[92], x[91], x[89], x[88], x[87], x[86], x[85], x[84], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[370], x[369], x[368], x[367], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[97], x[189], x[373], x[8], x[372], x[371]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[103], x[195], x[379], x[378], x[377], x[94], x[93], x[92], x[91], x[186], x[185], x[184], x[183], x[370], x[369], x[368], x[367], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[366], x[365], x[364], x[363], x[362], x[361], x[360], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[100], x[192], x[376], x[8], x[375], x[374]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[123], x[215], x[399], x[398], x[397], x[120], x[212], x[396], x[395], x[394], x[117], x[116], x[115], x[114], x[209], x[208], x[207], x[206], x[393], x[392], x[391], x[390], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[106], x[198], x[382], x[8], x[381], x[380]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[126], x[218], x[402], x[401], x[400], x[120], x[212], x[396], x[395], x[394], x[117], x[116], x[115], x[114], x[209], x[208], x[207], x[206], x[393], x[392], x[391], x[390], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[106], x[198], x[382], x[8], x[381], x[380]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[123], x[215], x[399], x[398], x[397], x[117], x[116], x[115], x[114], x[209], x[208], x[207], x[206], x[393], x[392], x[391], x[390], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[106], x[198], x[382], x[8], x[381], x[380]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[126], x[218], x[402], x[401], x[400], x[117], x[116], x[115], x[114], x[209], x[208], x[207], x[206], x[393], x[392], x[391], x[390], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[106], x[198], x[382], x[8], x[381], x[380]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[113], x[205], x[389], x[123], x[215], x[399], x[398], x[397], x[117], x[116], x[115], x[114], x[112], x[111], x[110], x[109], x[108], x[107], x[209], x[208], x[207], x[206], x[204], x[203], x[202], x[201], x[200], x[199], x[393], x[392], x[391], x[390], x[388], x[387], x[386], x[385], x[384], x[383], x[120], x[212], x[396], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[395], x[394]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[113], x[205], x[389], x[126], x[218], x[402], x[401], x[400], x[117], x[116], x[115], x[114], x[112], x[111], x[110], x[109], x[108], x[107], x[209], x[208], x[207], x[206], x[204], x[203], x[202], x[201], x[200], x[199], x[393], x[392], x[391], x[390], x[388], x[387], x[386], x[385], x[384], x[383], x[120], x[212], x[396], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[395], x[394]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[126], x[218], x[402], x[401], x[400], x[117], x[116], x[115], x[114], x[209], x[208], x[207], x[206], x[393], x[392], x[391], x[390], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[123], x[215], x[399], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[398], x[397]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[146], x[238], x[422], x[421], x[420], x[143], x[235], x[419], x[418], x[417], x[140], x[139], x[138], x[137], x[232], x[231], x[230], x[229], x[416], x[415], x[414], x[413], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[129], x[221], x[405], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[404], x[403]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[149], x[241], x[425], x[424], x[423], x[143], x[235], x[419], x[418], x[417], x[140], x[139], x[138], x[137], x[232], x[231], x[230], x[229], x[416], x[415], x[414], x[413], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[129], x[221], x[405], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[404], x[403]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[146], x[238], x[422], x[421], x[420], x[140], x[139], x[138], x[137], x[232], x[231], x[230], x[229], x[416], x[415], x[414], x[413], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[129], x[221], x[405], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[404], x[403]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[149], x[241], x[425], x[424], x[423], x[140], x[139], x[138], x[137], x[232], x[231], x[230], x[229], x[416], x[415], x[414], x[413], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[129], x[221], x[405], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[404], x[403]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[136], x[228], x[412], x[146], x[238], x[422], x[421], x[420], x[140], x[139], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[232], x[231], x[230], x[229], x[227], x[226], x[225], x[224], x[223], x[222], x[416], x[415], x[414], x[413], x[411], x[410], x[409], x[408], x[407], x[406], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[143], x[235], x[419], x[8], x[418], x[417]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[136], x[228], x[412], x[149], x[241], x[425], x[424], x[423], x[140], x[139], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[232], x[231], x[230], x[229], x[227], x[226], x[225], x[224], x[223], x[222], x[416], x[415], x[414], x[413], x[411], x[410], x[409], x[408], x[407], x[406], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[143], x[235], x[419], x[8], x[418], x[417]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[149], x[241], x[425], x[424], x[423], x[140], x[139], x[138], x[137], x[232], x[231], x[230], x[229], x[416], x[415], x[414], x[413], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[146], x[238], x[422], x[8], x[421], x[420]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[169], x[261], x[445], x[444], x[443], x[166], x[258], x[442], x[441], x[440], x[163], x[162], x[161], x[160], x[255], x[254], x[253], x[252], x[439], x[438], x[437], x[436], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[152], x[244], x[428], x[8], x[427], x[426]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[172], x[264], x[448], x[447], x[446], x[166], x[258], x[442], x[441], x[440], x[163], x[162], x[161], x[160], x[255], x[254], x[253], x[252], x[439], x[438], x[437], x[436], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[152], x[244], x[428], x[8], x[427], x[426]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[169], x[261], x[445], x[444], x[443], x[163], x[162], x[161], x[160], x[255], x[254], x[253], x[252], x[439], x[438], x[437], x[436], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[152], x[244], x[428], x[8], x[427], x[426]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[172], x[264], x[448], x[447], x[446], x[163], x[162], x[161], x[160], x[255], x[254], x[253], x[252], x[439], x[438], x[437], x[436], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[152], x[244], x[428], x[8], x[427], x[426]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[159], x[251], x[435], x[169], x[261], x[445], x[444], x[443], x[163], x[162], x[161], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[255], x[254], x[253], x[252], x[250], x[249], x[248], x[247], x[246], x[245], x[439], x[438], x[437], x[436], x[434], x[433], x[432], x[431], x[430], x[429], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[166], x[258], x[442], x[8], x[441], x[440]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[159], x[251], x[435], x[172], x[264], x[448], x[447], x[446], x[163], x[162], x[161], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[255], x[254], x[253], x[252], x[250], x[249], x[248], x[247], x[246], x[245], x[439], x[438], x[437], x[436], x[434], x[433], x[432], x[431], x[430], x[429], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[166], x[258], x[442], x[8], x[441], x[440]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[172], x[264], x[448], x[447], x[446], x[163], x[162], x[161], x[160], x[255], x[254], x[253], x[252], x[439], x[438], x[437], x[436], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[169], x[261], x[445], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[8], x[444], x[443]}), .y(y[188]));
endmodule

