/* modified netlist. Source: module AES in file /mnt/c/Users/Amir/Desktop/Papers_in_progress/AGEMA/Designs/AES_serial/AGEMA/sbox_opt3/AES.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module AES_HPC2_BDDsylvan_Pipeline_d1 (plaintext_s0, key_s0, clk, start, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [430:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_677 ;
    wire signal_679 ;
    wire signal_681 ;
    wire signal_683 ;
    wire signal_685 ;
    wire signal_687 ;
    wire signal_689 ;
    wire signal_691 ;
    wire signal_693 ;
    wire signal_695 ;
    wire signal_697 ;
    wire signal_699 ;
    wire signal_701 ;
    wire signal_703 ;
    wire signal_705 ;
    wire signal_707 ;
    wire signal_709 ;
    wire signal_711 ;
    wire signal_713 ;
    wire signal_715 ;
    wire signal_717 ;
    wire signal_719 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2447 ;
    wire signal_2450 ;
    wire signal_2453 ;
    wire signal_2456 ;
    wire signal_2459 ;
    wire signal_2462 ;
    wire signal_2465 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2474 ;
    wire signal_2476 ;
    wire signal_2478 ;
    wire signal_2481 ;
    wire signal_2483 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2579 ;
    wire signal_2582 ;
    wire signal_2585 ;
    wire signal_2588 ;
    wire signal_2591 ;
    wire signal_2594 ;
    wire signal_2597 ;
    wire signal_2600 ;
    wire signal_2603 ;
    wire signal_2606 ;
    wire signal_2609 ;
    wire signal_2612 ;
    wire signal_2615 ;
    wire signal_2618 ;
    wire signal_2621 ;
    wire signal_2624 ;
    wire signal_2627 ;
    wire signal_2630 ;
    wire signal_2633 ;
    wire signal_2636 ;
    wire signal_2639 ;
    wire signal_2642 ;
    wire signal_2645 ;
    wire signal_2648 ;
    wire signal_2651 ;
    wire signal_2654 ;
    wire signal_2657 ;
    wire signal_2660 ;
    wire signal_2663 ;
    wire signal_2666 ;
    wire signal_2669 ;
    wire signal_2672 ;
    wire signal_2675 ;
    wire signal_2678 ;
    wire signal_2681 ;
    wire signal_2684 ;
    wire signal_2687 ;
    wire signal_2690 ;
    wire signal_2693 ;
    wire signal_2696 ;
    wire signal_2699 ;
    wire signal_2702 ;
    wire signal_2705 ;
    wire signal_2708 ;
    wire signal_2711 ;
    wire signal_2714 ;
    wire signal_2717 ;
    wire signal_2720 ;
    wire signal_2723 ;
    wire signal_2726 ;
    wire signal_2729 ;
    wire signal_2732 ;
    wire signal_2735 ;
    wire signal_2738 ;
    wire signal_2741 ;
    wire signal_2744 ;
    wire signal_2747 ;
    wire signal_2750 ;
    wire signal_2753 ;
    wire signal_2756 ;
    wire signal_2759 ;
    wire signal_2762 ;
    wire signal_2765 ;
    wire signal_2768 ;
    wire signal_2771 ;
    wire signal_2774 ;
    wire signal_2777 ;
    wire signal_2780 ;
    wire signal_2783 ;
    wire signal_2786 ;
    wire signal_2789 ;
    wire signal_2792 ;
    wire signal_2795 ;
    wire signal_2798 ;
    wire signal_2801 ;
    wire signal_2804 ;
    wire signal_2807 ;
    wire signal_2810 ;
    wire signal_2813 ;
    wire signal_2816 ;
    wire signal_2819 ;
    wire signal_2822 ;
    wire signal_2825 ;
    wire signal_2828 ;
    wire signal_2831 ;
    wire signal_2834 ;
    wire signal_2837 ;
    wire signal_2840 ;
    wire signal_2843 ;
    wire signal_2846 ;
    wire signal_2849 ;
    wire signal_2852 ;
    wire signal_2855 ;
    wire signal_2858 ;
    wire signal_2861 ;
    wire signal_2864 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3202 ;
    wire signal_3204 ;
    wire signal_3206 ;
    wire signal_3208 ;
    wire signal_3210 ;
    wire signal_3212 ;
    wire signal_3214 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3628 ;
    wire signal_3630 ;
    wire signal_3632 ;
    wire signal_3634 ;
    wire signal_3636 ;
    wire signal_3638 ;
    wire signal_3640 ;
    wire signal_3642 ;
    wire signal_3644 ;
    wire signal_3646 ;
    wire signal_3648 ;
    wire signal_3650 ;
    wire signal_3652 ;
    wire signal_3654 ;
    wire signal_3656 ;
    wire signal_3658 ;
    wire signal_3660 ;
    wire signal_3662 ;
    wire signal_3664 ;
    wire signal_3666 ;
    wire signal_3668 ;
    wire signal_3670 ;
    wire signal_3672 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3941 ;
    wire signal_3943 ;
    wire signal_3945 ;
    wire signal_3947 ;
    wire signal_3949 ;
    wire signal_3951 ;
    wire signal_3953 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4221 ;
    wire signal_4223 ;
    wire signal_4225 ;
    wire signal_4227 ;
    wire signal_4229 ;
    wire signal_4231 ;
    wire signal_4233 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7759 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7762 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7765 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7768 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7771 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7774 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7777 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7780 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7783 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7786 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7789 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7792 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7795 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7798 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7801 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7804 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7807 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7810 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7813 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7816 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7819 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7822 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7825 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7828 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7831 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7834 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7837 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7840 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;
    wire signal_7973 ;
    wire signal_7974 ;
    wire signal_7975 ;
    wire signal_7976 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_8256 ;
    wire signal_8257 ;
    wire signal_8258 ;
    wire signal_8259 ;
    wire signal_8260 ;
    wire signal_8261 ;
    wire signal_8262 ;
    wire signal_8263 ;
    wire signal_8264 ;
    wire signal_8265 ;
    wire signal_8266 ;
    wire signal_8267 ;
    wire signal_8268 ;
    wire signal_8269 ;
    wire signal_8270 ;
    wire signal_8271 ;
    wire signal_8272 ;
    wire signal_8273 ;
    wire signal_8274 ;
    wire signal_8275 ;
    wire signal_8276 ;
    wire signal_8277 ;
    wire signal_8278 ;
    wire signal_8279 ;
    wire signal_8280 ;
    wire signal_8281 ;
    wire signal_8282 ;
    wire signal_8283 ;
    wire signal_8284 ;
    wire signal_8285 ;
    wire signal_8286 ;
    wire signal_8287 ;
    wire signal_8288 ;
    wire signal_8289 ;
    wire signal_8290 ;
    wire signal_8291 ;
    wire signal_8292 ;
    wire signal_8293 ;
    wire signal_8294 ;
    wire signal_8295 ;
    wire signal_8296 ;
    wire signal_8297 ;
    wire signal_8298 ;
    wire signal_8299 ;
    wire signal_8300 ;
    wire signal_8301 ;
    wire signal_8302 ;
    wire signal_8303 ;
    wire signal_8304 ;
    wire signal_8305 ;
    wire signal_8306 ;
    wire signal_8307 ;
    wire signal_8308 ;
    wire signal_8309 ;
    wire signal_8310 ;
    wire signal_8311 ;
    wire signal_8312 ;
    wire signal_8313 ;
    wire signal_8314 ;
    wire signal_8315 ;
    wire signal_8316 ;
    wire signal_8317 ;
    wire signal_8318 ;
    wire signal_8319 ;
    wire signal_8320 ;
    wire signal_8321 ;
    wire signal_8322 ;
    wire signal_8323 ;
    wire signal_8324 ;
    wire signal_8325 ;
    wire signal_8326 ;
    wire signal_8327 ;
    wire signal_8328 ;
    wire signal_8329 ;
    wire signal_8330 ;
    wire signal_8331 ;
    wire signal_8332 ;
    wire signal_8333 ;
    wire signal_8334 ;
    wire signal_8335 ;
    wire signal_8336 ;
    wire signal_8337 ;
    wire signal_8338 ;
    wire signal_8339 ;
    wire signal_8340 ;
    wire signal_8341 ;
    wire signal_8342 ;
    wire signal_8343 ;
    wire signal_8344 ;
    wire signal_8345 ;
    wire signal_8346 ;
    wire signal_8347 ;
    wire signal_8348 ;
    wire signal_8349 ;
    wire signal_8350 ;
    wire signal_8351 ;
    wire signal_8352 ;
    wire signal_8353 ;
    wire signal_8354 ;
    wire signal_8355 ;
    wire signal_8356 ;
    wire signal_8357 ;
    wire signal_8358 ;
    wire signal_8359 ;
    wire signal_8360 ;
    wire signal_8361 ;
    wire signal_8362 ;
    wire signal_8363 ;
    wire signal_8364 ;
    wire signal_8365 ;
    wire signal_8366 ;
    wire signal_8367 ;
    wire signal_8368 ;
    wire signal_8369 ;
    wire signal_8370 ;
    wire signal_8371 ;
    wire signal_8372 ;
    wire signal_8373 ;
    wire signal_8374 ;
    wire signal_8375 ;
    wire signal_8376 ;
    wire signal_8377 ;
    wire signal_8378 ;
    wire signal_8379 ;
    wire signal_8380 ;
    wire signal_8381 ;
    wire signal_8382 ;
    wire signal_8383 ;
    wire signal_8384 ;
    wire signal_8385 ;
    wire signal_8386 ;
    wire signal_8387 ;
    wire signal_8388 ;
    wire signal_8389 ;
    wire signal_8390 ;
    wire signal_8391 ;
    wire signal_8392 ;
    wire signal_8393 ;
    wire signal_8394 ;
    wire signal_8395 ;
    wire signal_8396 ;
    wire signal_8397 ;
    wire signal_8398 ;
    wire signal_8399 ;
    wire signal_8400 ;
    wire signal_8401 ;
    wire signal_8402 ;
    wire signal_8403 ;
    wire signal_8404 ;
    wire signal_8405 ;
    wire signal_8406 ;
    wire signal_8407 ;
    wire signal_8408 ;
    wire signal_8409 ;
    wire signal_8410 ;
    wire signal_8411 ;
    wire signal_8412 ;
    wire signal_8413 ;
    wire signal_8414 ;
    wire signal_8415 ;
    wire signal_8416 ;
    wire signal_8417 ;
    wire signal_8418 ;
    wire signal_8419 ;
    wire signal_8420 ;
    wire signal_8421 ;
    wire signal_8422 ;
    wire signal_8423 ;
    wire signal_8424 ;
    wire signal_8425 ;
    wire signal_8426 ;
    wire signal_8427 ;
    wire signal_8428 ;
    wire signal_8429 ;
    wire signal_8430 ;
    wire signal_8431 ;
    wire signal_8432 ;
    wire signal_8433 ;
    wire signal_8434 ;
    wire signal_8435 ;
    wire signal_8436 ;
    wire signal_8437 ;
    wire signal_8438 ;
    wire signal_8439 ;
    wire signal_8440 ;
    wire signal_8441 ;
    wire signal_8442 ;
    wire signal_8443 ;
    wire signal_8444 ;
    wire signal_8445 ;
    wire signal_8446 ;
    wire signal_8447 ;
    wire signal_8448 ;
    wire signal_8449 ;
    wire signal_8450 ;
    wire signal_8451 ;
    wire signal_8452 ;
    wire signal_8453 ;
    wire signal_8454 ;
    wire signal_8455 ;
    wire signal_8456 ;
    wire signal_8457 ;
    wire signal_8458 ;
    wire signal_8459 ;
    wire signal_8460 ;
    wire signal_8461 ;
    wire signal_8462 ;
    wire signal_8463 ;
    wire signal_8464 ;
    wire signal_8465 ;
    wire signal_8466 ;
    wire signal_8467 ;
    wire signal_8468 ;
    wire signal_8469 ;
    wire signal_8470 ;
    wire signal_8471 ;
    wire signal_8472 ;
    wire signal_8473 ;
    wire signal_8474 ;
    wire signal_8475 ;
    wire signal_8476 ;
    wire signal_8477 ;
    wire signal_8478 ;
    wire signal_8479 ;
    wire signal_8480 ;
    wire signal_8481 ;
    wire signal_8482 ;
    wire signal_8483 ;
    wire signal_8484 ;
    wire signal_8485 ;
    wire signal_8486 ;
    wire signal_8487 ;
    wire signal_8488 ;
    wire signal_8489 ;
    wire signal_8490 ;
    wire signal_8491 ;
    wire signal_8492 ;
    wire signal_8493 ;
    wire signal_8494 ;
    wire signal_8495 ;
    wire signal_8496 ;
    wire signal_8497 ;
    wire signal_8498 ;
    wire signal_8499 ;
    wire signal_8500 ;
    wire signal_8501 ;
    wire signal_8502 ;
    wire signal_8503 ;
    wire signal_8504 ;
    wire signal_8505 ;
    wire signal_8506 ;
    wire signal_8507 ;
    wire signal_8508 ;
    wire signal_8509 ;
    wire signal_8510 ;
    wire signal_8511 ;
    wire signal_8512 ;
    wire signal_8513 ;
    wire signal_8514 ;
    wire signal_8515 ;
    wire signal_8516 ;
    wire signal_8517 ;
    wire signal_8518 ;
    wire signal_8519 ;
    wire signal_8520 ;
    wire signal_8521 ;
    wire signal_8522 ;
    wire signal_8523 ;
    wire signal_8524 ;
    wire signal_8525 ;
    wire signal_8526 ;
    wire signal_8527 ;
    wire signal_8528 ;
    wire signal_8529 ;
    wire signal_8530 ;
    wire signal_8531 ;
    wire signal_8532 ;
    wire signal_8533 ;
    wire signal_8534 ;
    wire signal_8535 ;
    wire signal_8536 ;
    wire signal_8537 ;
    wire signal_8538 ;
    wire signal_8539 ;
    wire signal_8540 ;
    wire signal_8541 ;
    wire signal_8542 ;
    wire signal_8543 ;
    wire signal_8544 ;
    wire signal_8545 ;
    wire signal_8546 ;
    wire signal_8547 ;
    wire signal_8548 ;
    wire signal_8549 ;
    wire signal_8550 ;
    wire signal_8551 ;
    wire signal_8552 ;
    wire signal_8553 ;
    wire signal_8554 ;
    wire signal_8555 ;
    wire signal_8556 ;
    wire signal_8557 ;
    wire signal_8558 ;
    wire signal_8559 ;
    wire signal_8560 ;
    wire signal_8561 ;
    wire signal_8562 ;
    wire signal_8563 ;
    wire signal_8564 ;
    wire signal_8565 ;
    wire signal_8566 ;
    wire signal_8567 ;
    wire signal_8568 ;
    wire signal_8569 ;
    wire signal_8570 ;
    wire signal_8571 ;
    wire signal_8572 ;
    wire signal_8573 ;
    wire signal_8574 ;
    wire signal_8575 ;
    wire signal_8576 ;
    wire signal_8577 ;
    wire signal_8578 ;
    wire signal_8579 ;
    wire signal_8580 ;
    wire signal_8581 ;
    wire signal_8582 ;
    wire signal_8583 ;
    wire signal_8584 ;
    wire signal_8585 ;
    wire signal_8586 ;
    wire signal_8587 ;
    wire signal_8588 ;
    wire signal_8589 ;
    wire signal_8590 ;
    wire signal_8591 ;
    wire signal_8592 ;
    wire signal_8593 ;
    wire signal_8594 ;
    wire signal_8595 ;
    wire signal_8596 ;
    wire signal_8597 ;
    wire signal_8598 ;
    wire signal_8599 ;
    wire signal_8600 ;
    wire signal_8601 ;
    wire signal_8602 ;
    wire signal_8603 ;
    wire signal_8604 ;
    wire signal_8605 ;
    wire signal_8606 ;
    wire signal_8607 ;
    wire signal_8608 ;
    wire signal_8609 ;
    wire signal_8610 ;
    wire signal_8611 ;
    wire signal_8612 ;
    wire signal_8613 ;
    wire signal_8614 ;
    wire signal_8615 ;
    wire signal_8616 ;
    wire signal_8617 ;
    wire signal_8618 ;
    wire signal_8619 ;
    wire signal_8620 ;
    wire signal_8621 ;
    wire signal_8622 ;
    wire signal_8623 ;
    wire signal_8624 ;
    wire signal_8625 ;
    wire signal_8626 ;
    wire signal_8627 ;
    wire signal_8628 ;
    wire signal_8629 ;
    wire signal_8630 ;
    wire signal_8631 ;
    wire signal_8632 ;
    wire signal_8633 ;
    wire signal_8634 ;
    wire signal_8635 ;
    wire signal_8636 ;
    wire signal_8637 ;
    wire signal_8638 ;
    wire signal_8639 ;
    wire signal_8640 ;
    wire signal_8641 ;
    wire signal_8642 ;
    wire signal_8643 ;
    wire signal_8644 ;
    wire signal_8645 ;
    wire signal_8646 ;
    wire signal_8647 ;
    wire signal_8648 ;
    wire signal_8649 ;
    wire signal_8650 ;
    wire signal_8651 ;
    wire signal_8652 ;
    wire signal_8653 ;
    wire signal_8654 ;
    wire signal_8655 ;
    wire signal_8656 ;
    wire signal_8657 ;
    wire signal_8658 ;
    wire signal_8659 ;
    wire signal_8660 ;
    wire signal_8661 ;
    wire signal_8662 ;
    wire signal_8663 ;
    wire signal_8664 ;
    wire signal_8665 ;
    wire signal_8666 ;
    wire signal_8667 ;
    wire signal_8668 ;
    wire signal_8669 ;
    wire signal_8670 ;
    wire signal_8671 ;
    wire signal_8672 ;
    wire signal_8673 ;
    wire signal_8674 ;
    wire signal_8675 ;
    wire signal_8676 ;
    wire signal_8677 ;
    wire signal_8678 ;
    wire signal_8679 ;
    wire signal_8680 ;
    wire signal_8681 ;
    wire signal_8682 ;
    wire signal_8683 ;
    wire signal_8684 ;
    wire signal_8685 ;
    wire signal_8686 ;
    wire signal_8687 ;
    wire signal_8688 ;
    wire signal_8689 ;
    wire signal_8690 ;
    wire signal_8691 ;
    wire signal_8692 ;
    wire signal_8693 ;
    wire signal_8694 ;
    wire signal_8695 ;
    wire signal_8696 ;
    wire signal_8697 ;
    wire signal_8698 ;
    wire signal_8699 ;
    wire signal_8700 ;
    wire signal_8701 ;
    wire signal_8702 ;
    wire signal_8703 ;
    wire signal_8704 ;
    wire signal_8705 ;
    wire signal_8706 ;
    wire signal_8707 ;
    wire signal_8708 ;
    wire signal_8709 ;
    wire signal_8710 ;
    wire signal_8711 ;
    wire signal_8712 ;
    wire signal_8713 ;
    wire signal_8714 ;
    wire signal_8715 ;
    wire signal_8716 ;
    wire signal_8717 ;
    wire signal_8718 ;
    wire signal_8719 ;
    wire signal_8720 ;
    wire signal_8721 ;
    wire signal_8722 ;
    wire signal_8723 ;
    wire signal_8724 ;
    wire signal_8725 ;
    wire signal_8726 ;
    wire signal_8727 ;
    wire signal_8728 ;
    wire signal_8729 ;
    wire signal_8730 ;
    wire signal_8731 ;
    wire signal_8732 ;
    wire signal_8733 ;
    wire signal_8734 ;
    wire signal_8735 ;
    wire signal_8736 ;
    wire signal_8737 ;
    wire signal_8738 ;
    wire signal_8739 ;
    wire signal_8740 ;
    wire signal_8741 ;
    wire signal_8742 ;
    wire signal_8743 ;
    wire signal_8744 ;
    wire signal_8745 ;
    wire signal_8746 ;
    wire signal_8747 ;
    wire signal_8748 ;
    wire signal_8749 ;
    wire signal_8750 ;
    wire signal_8751 ;
    wire signal_8752 ;
    wire signal_8753 ;
    wire signal_8754 ;
    wire signal_8755 ;
    wire signal_8756 ;
    wire signal_8757 ;
    wire signal_8758 ;
    wire signal_8759 ;
    wire signal_8760 ;
    wire signal_8761 ;
    wire signal_8762 ;
    wire signal_8763 ;
    wire signal_8764 ;
    wire signal_8765 ;
    wire signal_8766 ;
    wire signal_8767 ;
    wire signal_8768 ;
    wire signal_8769 ;
    wire signal_8770 ;
    wire signal_8771 ;
    wire signal_8772 ;
    wire signal_8773 ;
    wire signal_8774 ;
    wire signal_8775 ;
    wire signal_8776 ;
    wire signal_8777 ;
    wire signal_8778 ;
    wire signal_8779 ;
    wire signal_8780 ;
    wire signal_8781 ;
    wire signal_8782 ;
    wire signal_8783 ;
    wire signal_8784 ;
    wire signal_8785 ;
    wire signal_8786 ;
    wire signal_8787 ;
    wire signal_8788 ;
    wire signal_8789 ;
    wire signal_8790 ;
    wire signal_8791 ;
    wire signal_8792 ;
    wire signal_8793 ;
    wire signal_8794 ;
    wire signal_8795 ;
    wire signal_8796 ;
    wire signal_8797 ;
    wire signal_8798 ;
    wire signal_8799 ;
    wire signal_8800 ;
    wire signal_8801 ;
    wire signal_8802 ;
    wire signal_8803 ;
    wire signal_8804 ;
    wire signal_8805 ;
    wire signal_8806 ;
    wire signal_8807 ;
    wire signal_8808 ;
    wire signal_8809 ;
    wire signal_8810 ;
    wire signal_8811 ;
    wire signal_8812 ;
    wire signal_8813 ;
    wire signal_8814 ;
    wire signal_8815 ;
    wire signal_8816 ;
    wire signal_8817 ;
    wire signal_8818 ;
    wire signal_8819 ;
    wire signal_8820 ;
    wire signal_8821 ;
    wire signal_8822 ;
    wire signal_8823 ;
    wire signal_8824 ;
    wire signal_8825 ;
    wire signal_8826 ;
    wire signal_8827 ;
    wire signal_8828 ;
    wire signal_8829 ;
    wire signal_8830 ;
    wire signal_8831 ;
    wire signal_8832 ;
    wire signal_8833 ;
    wire signal_8834 ;
    wire signal_8835 ;
    wire signal_8836 ;
    wire signal_8837 ;
    wire signal_8838 ;
    wire signal_8839 ;
    wire signal_8840 ;
    wire signal_8841 ;
    wire signal_8842 ;
    wire signal_8843 ;
    wire signal_8844 ;
    wire signal_8845 ;
    wire signal_8846 ;
    wire signal_8847 ;
    wire signal_8848 ;
    wire signal_8849 ;
    wire signal_8850 ;
    wire signal_8851 ;
    wire signal_8852 ;
    wire signal_8853 ;
    wire signal_8854 ;
    wire signal_8855 ;
    wire signal_8856 ;
    wire signal_8857 ;
    wire signal_8858 ;
    wire signal_8859 ;
    wire signal_8860 ;
    wire signal_8861 ;
    wire signal_8862 ;
    wire signal_8863 ;
    wire signal_8864 ;
    wire signal_8865 ;
    wire signal_8866 ;
    wire signal_8867 ;
    wire signal_8868 ;
    wire signal_8869 ;
    wire signal_8870 ;
    wire signal_8871 ;
    wire signal_8872 ;
    wire signal_8873 ;
    wire signal_8874 ;
    wire signal_8875 ;
    wire signal_8876 ;
    wire signal_8877 ;
    wire signal_8878 ;
    wire signal_8879 ;
    wire signal_8880 ;
    wire signal_8881 ;
    wire signal_8882 ;
    wire signal_8883 ;
    wire signal_8884 ;
    wire signal_8885 ;
    wire signal_8886 ;
    wire signal_8887 ;
    wire signal_8888 ;
    wire signal_8889 ;
    wire signal_8890 ;
    wire signal_8891 ;
    wire signal_8892 ;
    wire signal_8893 ;
    wire signal_8894 ;
    wire signal_8895 ;
    wire signal_8896 ;
    wire signal_8897 ;
    wire signal_8898 ;
    wire signal_8899 ;
    wire signal_8900 ;
    wire signal_8901 ;
    wire signal_8902 ;
    wire signal_8903 ;
    wire signal_8904 ;
    wire signal_8905 ;
    wire signal_8906 ;
    wire signal_8907 ;
    wire signal_8908 ;
    wire signal_8909 ;
    wire signal_8910 ;
    wire signal_8911 ;
    wire signal_8912 ;
    wire signal_8913 ;
    wire signal_8914 ;
    wire signal_8915 ;
    wire signal_8916 ;
    wire signal_8917 ;
    wire signal_8918 ;
    wire signal_8919 ;
    wire signal_8920 ;
    wire signal_8921 ;
    wire signal_8922 ;
    wire signal_8923 ;
    wire signal_8924 ;
    wire signal_8925 ;
    wire signal_8926 ;
    wire signal_8927 ;
    wire signal_8928 ;
    wire signal_8929 ;
    wire signal_8930 ;
    wire signal_8931 ;
    wire signal_8932 ;
    wire signal_8933 ;
    wire signal_8934 ;
    wire signal_8935 ;
    wire signal_8936 ;
    wire signal_8937 ;
    wire signal_8938 ;
    wire signal_8939 ;
    wire signal_8940 ;
    wire signal_8941 ;
    wire signal_8942 ;
    wire signal_8943 ;
    wire signal_8944 ;
    wire signal_8945 ;
    wire signal_8946 ;
    wire signal_8947 ;
    wire signal_8948 ;
    wire signal_8949 ;
    wire signal_8950 ;
    wire signal_8951 ;
    wire signal_8952 ;
    wire signal_8953 ;
    wire signal_8954 ;
    wire signal_8955 ;
    wire signal_8956 ;
    wire signal_8957 ;
    wire signal_8958 ;
    wire signal_8959 ;
    wire signal_8960 ;
    wire signal_8961 ;
    wire signal_8962 ;
    wire signal_8963 ;
    wire signal_8964 ;
    wire signal_8965 ;
    wire signal_8966 ;
    wire signal_8967 ;
    wire signal_8968 ;
    wire signal_8969 ;
    wire signal_8970 ;
    wire signal_8971 ;
    wire signal_8972 ;
    wire signal_8973 ;
    wire signal_8974 ;
    wire signal_8975 ;
    wire signal_8976 ;
    wire signal_8977 ;
    wire signal_8978 ;
    wire signal_8979 ;
    wire signal_8980 ;
    wire signal_8981 ;
    wire signal_8982 ;
    wire signal_8983 ;
    wire signal_8984 ;
    wire signal_8985 ;
    wire signal_8986 ;
    wire signal_8987 ;
    wire signal_8988 ;
    wire signal_8989 ;
    wire signal_8990 ;
    wire signal_8991 ;
    wire signal_8992 ;
    wire signal_8993 ;
    wire signal_8994 ;
    wire signal_8995 ;
    wire signal_8996 ;
    wire signal_8997 ;
    wire signal_8998 ;
    wire signal_8999 ;
    wire signal_9000 ;
    wire signal_9001 ;
    wire signal_9002 ;
    wire signal_9003 ;
    wire signal_9004 ;
    wire signal_9005 ;
    wire signal_9006 ;
    wire signal_9007 ;
    wire signal_9008 ;
    wire signal_9009 ;
    wire signal_9010 ;
    wire signal_9011 ;
    wire signal_9012 ;
    wire signal_9013 ;
    wire signal_9014 ;
    wire signal_9015 ;
    wire signal_9016 ;
    wire signal_9017 ;
    wire signal_9018 ;
    wire signal_9019 ;
    wire signal_9020 ;
    wire signal_9021 ;
    wire signal_9022 ;
    wire signal_9023 ;
    wire signal_9024 ;
    wire signal_9025 ;
    wire signal_9026 ;
    wire signal_9027 ;
    wire signal_9028 ;
    wire signal_9029 ;
    wire signal_9030 ;
    wire signal_9031 ;
    wire signal_9032 ;
    wire signal_9033 ;
    wire signal_9034 ;
    wire signal_9035 ;
    wire signal_9036 ;
    wire signal_9037 ;
    wire signal_9038 ;
    wire signal_9039 ;
    wire signal_9040 ;
    wire signal_9041 ;
    wire signal_9042 ;
    wire signal_9043 ;
    wire signal_9044 ;
    wire signal_9045 ;
    wire signal_9046 ;
    wire signal_9047 ;
    wire signal_9048 ;
    wire signal_9049 ;
    wire signal_9050 ;
    wire signal_9051 ;
    wire signal_9052 ;
    wire signal_9053 ;
    wire signal_9054 ;
    wire signal_9055 ;
    wire signal_9056 ;
    wire signal_9057 ;
    wire signal_9058 ;
    wire signal_9059 ;
    wire signal_9060 ;
    wire signal_9061 ;
    wire signal_9062 ;
    wire signal_9063 ;
    wire signal_9064 ;
    wire signal_9065 ;
    wire signal_9066 ;
    wire signal_9067 ;
    wire signal_9068 ;
    wire signal_9069 ;
    wire signal_9070 ;
    wire signal_9071 ;
    wire signal_9072 ;
    wire signal_9073 ;
    wire signal_9074 ;
    wire signal_9075 ;
    wire signal_9076 ;
    wire signal_9077 ;
    wire signal_9078 ;
    wire signal_9079 ;
    wire signal_9080 ;
    wire signal_9081 ;
    wire signal_9082 ;
    wire signal_9083 ;
    wire signal_9084 ;
    wire signal_9085 ;
    wire signal_9086 ;
    wire signal_9087 ;
    wire signal_9088 ;
    wire signal_9089 ;
    wire signal_9090 ;
    wire signal_9091 ;
    wire signal_9092 ;
    wire signal_9093 ;
    wire signal_9094 ;
    wire signal_9095 ;
    wire signal_9096 ;
    wire signal_9097 ;
    wire signal_9098 ;
    wire signal_9099 ;
    wire signal_9100 ;
    wire signal_9101 ;
    wire signal_9102 ;
    wire signal_9103 ;
    wire signal_9104 ;
    wire signal_9105 ;
    wire signal_9106 ;
    wire signal_9107 ;
    wire signal_9108 ;
    wire signal_9109 ;
    wire signal_9110 ;
    wire signal_9111 ;
    wire signal_9112 ;
    wire signal_9113 ;
    wire signal_9114 ;
    wire signal_9115 ;
    wire signal_9116 ;
    wire signal_9117 ;
    wire signal_9118 ;
    wire signal_9119 ;
    wire signal_9120 ;
    wire signal_9121 ;
    wire signal_9122 ;
    wire signal_9123 ;
    wire signal_9124 ;
    wire signal_9125 ;
    wire signal_9126 ;
    wire signal_9127 ;
    wire signal_9128 ;
    wire signal_9129 ;
    wire signal_9130 ;
    wire signal_9131 ;
    wire signal_9132 ;
    wire signal_9133 ;
    wire signal_9134 ;
    wire signal_9135 ;
    wire signal_9136 ;
    wire signal_9137 ;
    wire signal_9138 ;
    wire signal_9139 ;
    wire signal_9140 ;
    wire signal_9141 ;
    wire signal_9142 ;
    wire signal_9143 ;
    wire signal_9144 ;
    wire signal_9145 ;
    wire signal_9146 ;
    wire signal_9147 ;
    wire signal_9148 ;
    wire signal_9149 ;
    wire signal_9150 ;
    wire signal_9151 ;
    wire signal_9152 ;
    wire signal_9153 ;
    wire signal_9154 ;
    wire signal_9155 ;
    wire signal_9156 ;
    wire signal_9157 ;
    wire signal_9158 ;
    wire signal_9159 ;
    wire signal_9160 ;
    wire signal_9161 ;
    wire signal_9162 ;
    wire signal_9163 ;
    wire signal_9164 ;
    wire signal_9165 ;
    wire signal_9166 ;
    wire signal_9167 ;
    wire signal_9168 ;
    wire signal_9169 ;
    wire signal_9170 ;
    wire signal_9171 ;
    wire signal_9172 ;
    wire signal_9173 ;
    wire signal_9174 ;
    wire signal_9175 ;
    wire signal_9176 ;
    wire signal_9177 ;
    wire signal_9178 ;
    wire signal_9179 ;
    wire signal_9180 ;
    wire signal_9181 ;
    wire signal_9182 ;
    wire signal_9183 ;
    wire signal_9184 ;
    wire signal_9185 ;
    wire signal_9186 ;
    wire signal_9187 ;
    wire signal_9188 ;
    wire signal_9189 ;
    wire signal_9190 ;
    wire signal_9191 ;
    wire signal_9192 ;
    wire signal_9193 ;
    wire signal_9194 ;
    wire signal_9195 ;
    wire signal_9196 ;
    wire signal_9197 ;
    wire signal_9198 ;
    wire signal_9199 ;
    wire signal_9200 ;
    wire signal_9201 ;
    wire signal_9202 ;
    wire signal_9203 ;
    wire signal_9204 ;
    wire signal_9205 ;
    wire signal_9206 ;
    wire signal_9207 ;
    wire signal_9208 ;
    wire signal_9209 ;
    wire signal_9210 ;
    wire signal_9211 ;
    wire signal_9212 ;
    wire signal_9213 ;
    wire signal_9214 ;
    wire signal_9215 ;
    wire signal_9216 ;
    wire signal_9217 ;
    wire signal_9218 ;
    wire signal_9219 ;
    wire signal_9220 ;
    wire signal_9221 ;
    wire signal_9222 ;
    wire signal_9223 ;
    wire signal_9224 ;
    wire signal_9225 ;
    wire signal_9226 ;
    wire signal_9227 ;
    wire signal_9228 ;
    wire signal_9229 ;
    wire signal_9230 ;
    wire signal_9231 ;
    wire signal_9232 ;
    wire signal_9233 ;
    wire signal_9234 ;
    wire signal_9235 ;
    wire signal_9236 ;
    wire signal_9237 ;
    wire signal_9238 ;
    wire signal_9239 ;
    wire signal_9240 ;
    wire signal_9241 ;
    wire signal_9242 ;
    wire signal_9243 ;
    wire signal_9244 ;
    wire signal_9245 ;
    wire signal_9246 ;
    wire signal_9247 ;
    wire signal_9248 ;
    wire signal_9249 ;
    wire signal_9250 ;
    wire signal_9251 ;
    wire signal_9252 ;
    wire signal_9253 ;
    wire signal_9254 ;
    wire signal_9255 ;
    wire signal_9256 ;
    wire signal_9257 ;
    wire signal_9258 ;
    wire signal_9259 ;
    wire signal_9260 ;
    wire signal_9261 ;
    wire signal_9262 ;
    wire signal_9263 ;
    wire signal_9264 ;
    wire signal_9265 ;
    wire signal_9266 ;
    wire signal_9267 ;
    wire signal_9268 ;
    wire signal_9269 ;
    wire signal_9270 ;
    wire signal_9271 ;
    wire signal_9272 ;
    wire signal_9273 ;
    wire signal_9274 ;
    wire signal_9275 ;
    wire signal_9276 ;
    wire signal_9277 ;
    wire signal_9278 ;
    wire signal_9279 ;
    wire signal_9280 ;
    wire signal_9281 ;
    wire signal_9282 ;
    wire signal_9283 ;
    wire signal_9284 ;
    wire signal_9285 ;
    wire signal_9286 ;
    wire signal_9287 ;
    wire signal_9288 ;
    wire signal_9289 ;
    wire signal_9290 ;
    wire signal_9291 ;
    wire signal_9292 ;
    wire signal_9293 ;
    wire signal_9294 ;
    wire signal_9295 ;
    wire signal_9296 ;
    wire signal_9297 ;
    wire signal_9298 ;
    wire signal_9299 ;
    wire signal_9300 ;
    wire signal_9301 ;
    wire signal_9302 ;
    wire signal_9303 ;
    wire signal_9304 ;
    wire signal_9305 ;
    wire signal_9306 ;
    wire signal_9307 ;
    wire signal_9308 ;
    wire signal_9309 ;
    wire signal_9310 ;
    wire signal_9311 ;
    wire signal_9312 ;
    wire signal_9313 ;
    wire signal_9314 ;
    wire signal_9315 ;
    wire signal_9316 ;
    wire signal_9317 ;
    wire signal_9318 ;
    wire signal_9319 ;
    wire signal_9320 ;
    wire signal_9321 ;
    wire signal_9322 ;
    wire signal_9323 ;
    wire signal_9324 ;
    wire signal_9325 ;
    wire signal_9326 ;
    wire signal_9327 ;
    wire signal_9328 ;
    wire signal_9329 ;
    wire signal_9330 ;
    wire signal_9331 ;
    wire signal_9332 ;
    wire signal_9333 ;
    wire signal_9334 ;
    wire signal_9335 ;
    wire signal_9336 ;
    wire signal_9337 ;
    wire signal_9338 ;
    wire signal_9339 ;
    wire signal_9340 ;
    wire signal_9341 ;
    wire signal_9342 ;
    wire signal_9343 ;
    wire signal_9344 ;
    wire signal_9345 ;
    wire signal_9346 ;
    wire signal_9347 ;
    wire signal_9348 ;
    wire signal_9349 ;
    wire signal_9350 ;
    wire signal_9351 ;
    wire signal_9352 ;
    wire signal_9353 ;
    wire signal_9354 ;
    wire signal_9355 ;
    wire signal_9356 ;
    wire signal_9357 ;
    wire signal_9358 ;
    wire signal_9359 ;
    wire signal_9360 ;
    wire signal_9361 ;
    wire signal_9362 ;
    wire signal_9363 ;
    wire signal_9364 ;
    wire signal_9365 ;
    wire signal_9366 ;
    wire signal_9367 ;
    wire signal_9368 ;
    wire signal_9369 ;
    wire signal_9370 ;
    wire signal_9371 ;
    wire signal_9372 ;
    wire signal_9373 ;
    wire signal_9374 ;
    wire signal_9375 ;
    wire signal_9376 ;
    wire signal_9377 ;
    wire signal_9378 ;
    wire signal_9379 ;
    wire signal_9380 ;
    wire signal_9381 ;
    wire signal_9382 ;
    wire signal_9383 ;
    wire signal_9384 ;
    wire signal_9385 ;
    wire signal_9386 ;
    wire signal_9387 ;
    wire signal_9388 ;
    wire signal_9389 ;
    wire signal_9390 ;
    wire signal_9391 ;
    wire signal_9392 ;
    wire signal_9393 ;
    wire signal_9394 ;
    wire signal_9395 ;
    wire signal_9396 ;
    wire signal_9397 ;
    wire signal_9398 ;
    wire signal_9399 ;
    wire signal_9400 ;
    wire signal_9401 ;
    wire signal_9402 ;
    wire signal_9403 ;
    wire signal_9404 ;
    wire signal_9405 ;
    wire signal_9406 ;
    wire signal_9407 ;
    wire signal_9408 ;
    wire signal_9409 ;
    wire signal_9410 ;
    wire signal_9411 ;
    wire signal_9412 ;
    wire signal_9413 ;
    wire signal_9414 ;
    wire signal_9415 ;
    wire signal_9416 ;
    wire signal_9417 ;
    wire signal_9418 ;
    wire signal_9419 ;
    wire signal_9420 ;
    wire signal_9421 ;
    wire signal_9422 ;
    wire signal_9423 ;
    wire signal_9424 ;
    wire signal_9425 ;
    wire signal_9426 ;
    wire signal_9427 ;
    wire signal_9428 ;
    wire signal_9429 ;
    wire signal_9430 ;
    wire signal_9431 ;
    wire signal_9432 ;
    wire signal_9433 ;
    wire signal_9434 ;
    wire signal_9435 ;
    wire signal_9436 ;
    wire signal_9437 ;
    wire signal_9438 ;
    wire signal_9439 ;
    wire signal_9440 ;
    wire signal_9441 ;
    wire signal_9442 ;
    wire signal_9443 ;
    wire signal_9444 ;
    wire signal_9445 ;
    wire signal_9446 ;
    wire signal_9447 ;
    wire signal_9448 ;
    wire signal_9449 ;
    wire signal_9450 ;
    wire signal_9451 ;
    wire signal_9452 ;
    wire signal_9453 ;
    wire signal_9454 ;
    wire signal_9455 ;
    wire signal_9456 ;
    wire signal_9457 ;
    wire signal_9458 ;
    wire signal_9459 ;
    wire signal_9460 ;
    wire signal_9461 ;
    wire signal_9462 ;
    wire signal_9463 ;
    wire signal_9464 ;
    wire signal_9465 ;
    wire signal_9466 ;
    wire signal_9467 ;
    wire signal_9468 ;
    wire signal_9469 ;
    wire signal_9470 ;
    wire signal_9471 ;
    wire signal_9472 ;
    wire signal_9473 ;
    wire signal_9474 ;
    wire signal_9475 ;
    wire signal_9476 ;
    wire signal_9477 ;
    wire signal_9478 ;
    wire signal_9479 ;
    wire signal_9480 ;
    wire signal_9481 ;
    wire signal_9482 ;
    wire signal_9483 ;
    wire signal_9484 ;
    wire signal_9485 ;
    wire signal_9486 ;
    wire signal_9487 ;
    wire signal_9488 ;
    wire signal_9489 ;
    wire signal_9490 ;
    wire signal_9491 ;
    wire signal_9492 ;
    wire signal_9493 ;
    wire signal_9494 ;
    wire signal_9495 ;
    wire signal_9496 ;
    wire signal_9497 ;
    wire signal_9498 ;
    wire signal_9499 ;
    wire signal_9500 ;
    wire signal_9501 ;
    wire signal_9502 ;
    wire signal_9503 ;
    wire signal_9504 ;
    wire signal_9505 ;
    wire signal_9506 ;
    wire signal_9507 ;
    wire signal_9508 ;
    wire signal_9509 ;
    wire signal_9510 ;
    wire signal_9511 ;
    wire signal_9512 ;
    wire signal_9513 ;
    wire signal_9514 ;
    wire signal_9515 ;
    wire signal_9516 ;
    wire signal_9517 ;
    wire signal_9518 ;
    wire signal_9519 ;
    wire signal_9520 ;
    wire signal_9521 ;
    wire signal_9522 ;
    wire signal_9523 ;
    wire signal_9524 ;
    wire signal_9525 ;
    wire signal_9526 ;
    wire signal_9527 ;
    wire signal_9528 ;
    wire signal_9529 ;
    wire signal_9530 ;
    wire signal_9531 ;
    wire signal_9532 ;
    wire signal_9533 ;
    wire signal_9534 ;
    wire signal_9535 ;
    wire signal_9536 ;
    wire signal_9537 ;
    wire signal_9538 ;
    wire signal_9539 ;
    wire signal_9540 ;
    wire signal_9541 ;
    wire signal_9542 ;
    wire signal_9543 ;
    wire signal_9544 ;
    wire signal_9545 ;
    wire signal_9546 ;
    wire signal_9547 ;
    wire signal_9548 ;
    wire signal_9549 ;
    wire signal_9550 ;
    wire signal_9551 ;
    wire signal_9552 ;
    wire signal_9553 ;
    wire signal_9554 ;
    wire signal_9555 ;
    wire signal_9556 ;
    wire signal_9557 ;
    wire signal_9558 ;
    wire signal_9559 ;
    wire signal_9560 ;
    wire signal_9561 ;
    wire signal_9562 ;
    wire signal_9563 ;
    wire signal_9564 ;
    wire signal_9565 ;
    wire signal_9566 ;
    wire signal_9567 ;
    wire signal_9568 ;
    wire signal_9569 ;
    wire signal_9570 ;
    wire signal_9571 ;
    wire signal_9572 ;
    wire signal_9573 ;
    wire signal_9574 ;
    wire signal_9575 ;
    wire signal_9576 ;
    wire signal_9577 ;
    wire signal_9578 ;
    wire signal_9579 ;
    wire signal_9580 ;
    wire signal_9581 ;
    wire signal_9582 ;
    wire signal_9583 ;
    wire signal_9584 ;
    wire signal_9585 ;
    wire signal_9586 ;
    wire signal_9587 ;
    wire signal_9588 ;
    wire signal_9589 ;
    wire signal_9590 ;
    wire signal_9591 ;
    wire signal_9592 ;
    wire signal_9593 ;
    wire signal_9594 ;
    wire signal_9595 ;
    wire signal_9596 ;
    wire signal_9597 ;
    wire signal_9598 ;
    wire signal_9599 ;
    wire signal_9600 ;
    wire signal_9601 ;
    wire signal_9602 ;
    wire signal_9603 ;
    wire signal_9604 ;
    wire signal_9605 ;
    wire signal_9606 ;
    wire signal_9607 ;
    wire signal_9608 ;
    wire signal_9609 ;
    wire signal_9610 ;
    wire signal_9611 ;
    wire signal_9612 ;
    wire signal_9613 ;
    wire signal_9614 ;
    wire signal_9615 ;
    wire signal_9616 ;
    wire signal_9617 ;
    wire signal_9618 ;
    wire signal_9619 ;
    wire signal_9620 ;
    wire signal_9621 ;
    wire signal_9622 ;
    wire signal_9623 ;
    wire signal_9624 ;
    wire signal_9625 ;
    wire signal_9626 ;
    wire signal_9627 ;
    wire signal_9628 ;
    wire signal_9629 ;
    wire signal_9630 ;
    wire signal_9631 ;
    wire signal_9632 ;
    wire signal_9633 ;
    wire signal_9634 ;
    wire signal_9635 ;
    wire signal_9636 ;
    wire signal_9637 ;
    wire signal_9638 ;
    wire signal_9639 ;
    wire signal_9640 ;
    wire signal_9641 ;
    wire signal_9642 ;
    wire signal_9643 ;
    wire signal_9644 ;
    wire signal_9645 ;
    wire signal_9646 ;
    wire signal_9647 ;
    wire signal_9648 ;
    wire signal_9649 ;
    wire signal_9650 ;
    wire signal_9651 ;
    wire signal_9652 ;
    wire signal_9653 ;
    wire signal_9654 ;
    wire signal_9655 ;
    wire signal_9656 ;
    wire signal_9657 ;
    wire signal_9658 ;
    wire signal_9659 ;
    wire signal_9660 ;
    wire signal_9661 ;
    wire signal_9662 ;
    wire signal_9663 ;
    wire signal_9664 ;
    wire signal_9665 ;
    wire signal_9666 ;
    wire signal_9667 ;
    wire signal_9668 ;
    wire signal_9669 ;
    wire signal_9670 ;
    wire signal_9671 ;
    wire signal_9672 ;
    wire signal_9673 ;
    wire signal_9674 ;
    wire signal_9675 ;
    wire signal_9676 ;
    wire signal_9677 ;
    wire signal_9678 ;
    wire signal_9679 ;
    wire signal_9680 ;
    wire signal_9681 ;
    wire signal_9682 ;
    wire signal_9683 ;
    wire signal_9684 ;
    wire signal_9685 ;
    wire signal_9686 ;
    wire signal_9687 ;
    wire signal_9688 ;
    wire signal_9689 ;
    wire signal_9690 ;
    wire signal_9691 ;
    wire signal_9692 ;
    wire signal_9693 ;
    wire signal_9694 ;
    wire signal_9695 ;
    wire signal_9696 ;
    wire signal_9697 ;
    wire signal_9698 ;
    wire signal_9699 ;
    wire signal_9700 ;
    wire signal_9701 ;
    wire signal_9702 ;
    wire signal_9703 ;
    wire signal_9704 ;
    wire signal_9705 ;
    wire signal_9706 ;
    wire signal_9707 ;
    wire signal_9708 ;
    wire signal_9709 ;
    wire signal_9710 ;
    wire signal_9711 ;
    wire signal_9712 ;
    wire signal_9713 ;
    wire signal_9714 ;
    wire signal_9715 ;
    wire signal_9716 ;
    wire signal_9717 ;
    wire signal_9718 ;
    wire signal_9719 ;
    wire signal_9720 ;
    wire signal_9721 ;
    wire signal_9722 ;
    wire signal_9723 ;
    wire signal_9724 ;
    wire signal_9725 ;
    wire signal_9726 ;
    wire signal_9727 ;
    wire signal_9728 ;
    wire signal_9729 ;
    wire signal_9730 ;
    wire signal_9731 ;
    wire signal_9732 ;
    wire signal_9733 ;
    wire signal_9734 ;
    wire signal_9735 ;
    wire signal_9736 ;
    wire signal_9737 ;
    wire signal_9738 ;
    wire signal_9739 ;
    wire signal_9740 ;
    wire signal_9741 ;
    wire signal_9742 ;
    wire signal_9743 ;
    wire signal_9744 ;
    wire signal_9745 ;
    wire signal_9746 ;
    wire signal_9747 ;
    wire signal_9748 ;
    wire signal_9749 ;
    wire signal_9750 ;
    wire signal_9751 ;
    wire signal_9752 ;
    wire signal_9753 ;
    wire signal_9754 ;
    wire signal_9755 ;
    wire signal_9756 ;
    wire signal_9757 ;
    wire signal_9758 ;
    wire signal_9759 ;
    wire signal_9760 ;
    wire signal_9761 ;
    wire signal_9762 ;
    wire signal_9763 ;
    wire signal_9764 ;
    wire signal_9765 ;
    wire signal_9766 ;
    wire signal_9767 ;
    wire signal_9768 ;
    wire signal_9769 ;
    wire signal_9770 ;
    wire signal_9771 ;
    wire signal_9772 ;
    wire signal_9773 ;
    wire signal_9774 ;
    wire signal_9775 ;
    wire signal_9776 ;
    wire signal_9777 ;
    wire signal_9778 ;
    wire signal_9779 ;
    wire signal_9780 ;
    wire signal_9781 ;
    wire signal_9782 ;
    wire signal_9783 ;
    wire signal_9784 ;
    wire signal_9785 ;
    wire signal_9786 ;
    wire signal_9787 ;
    wire signal_9788 ;
    wire signal_9789 ;
    wire signal_9790 ;
    wire signal_9791 ;
    wire signal_9792 ;
    wire signal_9793 ;
    wire signal_9794 ;
    wire signal_9795 ;
    wire signal_9796 ;
    wire signal_9797 ;
    wire signal_9798 ;
    wire signal_9799 ;
    wire signal_9800 ;
    wire signal_9801 ;
    wire signal_9802 ;
    wire signal_9803 ;
    wire signal_9804 ;
    wire signal_9805 ;
    wire signal_9806 ;
    wire signal_9807 ;
    wire signal_9808 ;
    wire signal_9809 ;
    wire signal_9810 ;
    wire signal_9811 ;
    wire signal_9812 ;
    wire signal_9813 ;
    wire signal_9814 ;
    wire signal_9815 ;
    wire signal_9816 ;
    wire signal_9817 ;
    wire signal_9818 ;
    wire signal_9819 ;
    wire signal_9820 ;
    wire signal_9821 ;
    wire signal_9822 ;
    wire signal_9823 ;
    wire signal_9824 ;
    wire signal_9825 ;
    wire signal_9826 ;
    wire signal_9827 ;
    wire signal_9828 ;
    wire signal_9829 ;
    wire signal_9830 ;
    wire signal_9831 ;
    wire signal_9832 ;
    wire signal_9833 ;
    wire signal_9834 ;
    wire signal_9835 ;
    wire signal_9836 ;
    wire signal_9837 ;
    wire signal_9838 ;
    wire signal_9839 ;
    wire signal_9840 ;
    wire signal_9841 ;
    wire signal_9842 ;
    wire signal_9843 ;
    wire signal_9844 ;
    wire signal_9845 ;
    wire signal_9846 ;
    wire signal_9847 ;
    wire signal_9848 ;
    wire signal_9849 ;
    wire signal_9850 ;
    wire signal_9851 ;
    wire signal_9852 ;
    wire signal_9853 ;
    wire signal_9854 ;
    wire signal_9855 ;
    wire signal_9856 ;
    wire signal_9857 ;
    wire signal_9858 ;
    wire signal_9859 ;
    wire signal_9860 ;
    wire signal_9861 ;
    wire signal_9862 ;
    wire signal_9863 ;
    wire signal_9864 ;
    wire signal_9865 ;
    wire signal_9866 ;
    wire signal_9867 ;
    wire signal_9868 ;
    wire signal_9869 ;
    wire signal_9870 ;
    wire signal_9871 ;
    wire signal_9872 ;
    wire signal_9873 ;
    wire signal_9874 ;
    wire signal_9875 ;
    wire signal_9876 ;
    wire signal_9877 ;
    wire signal_9878 ;
    wire signal_9879 ;
    wire signal_9880 ;
    wire signal_9881 ;
    wire signal_9882 ;
    wire signal_9883 ;
    wire signal_9884 ;
    wire signal_9885 ;
    wire signal_9886 ;
    wire signal_9887 ;
    wire signal_9888 ;
    wire signal_9889 ;
    wire signal_9890 ;
    wire signal_9891 ;
    wire signal_9892 ;
    wire signal_9893 ;
    wire signal_9894 ;
    wire signal_9895 ;
    wire signal_9896 ;
    wire signal_9897 ;
    wire signal_9898 ;
    wire signal_9899 ;
    wire signal_9900 ;
    wire signal_9901 ;
    wire signal_9902 ;
    wire signal_9903 ;
    wire signal_9904 ;
    wire signal_9905 ;
    wire signal_9906 ;
    wire signal_9907 ;
    wire signal_9908 ;
    wire signal_9909 ;
    wire signal_9910 ;
    wire signal_9911 ;
    wire signal_9912 ;
    wire signal_9913 ;
    wire signal_9914 ;
    wire signal_9915 ;
    wire signal_9916 ;
    wire signal_9917 ;
    wire signal_9918 ;
    wire signal_9919 ;
    wire signal_9920 ;
    wire signal_9921 ;
    wire signal_9922 ;
    wire signal_9923 ;
    wire signal_9924 ;
    wire signal_9925 ;
    wire signal_9926 ;
    wire signal_9927 ;
    wire signal_9928 ;
    wire signal_9929 ;
    wire signal_9930 ;
    wire signal_9931 ;
    wire signal_9932 ;
    wire signal_9933 ;
    wire signal_9934 ;
    wire signal_9935 ;
    wire signal_9936 ;
    wire signal_9937 ;
    wire signal_9938 ;
    wire signal_9939 ;
    wire signal_9940 ;
    wire signal_9941 ;
    wire signal_9942 ;
    wire signal_9943 ;
    wire signal_9944 ;
    wire signal_9945 ;
    wire signal_9946 ;
    wire signal_9947 ;
    wire signal_9948 ;
    wire signal_9949 ;
    wire signal_9950 ;
    wire signal_9951 ;
    wire signal_9952 ;
    wire signal_9953 ;
    wire signal_9954 ;
    wire signal_9955 ;
    wire signal_9956 ;
    wire signal_9957 ;
    wire signal_9958 ;
    wire signal_9959 ;
    wire signal_9960 ;
    wire signal_9961 ;
    wire signal_9962 ;
    wire signal_9963 ;
    wire signal_9964 ;
    wire signal_9965 ;
    wire signal_9966 ;
    wire signal_9967 ;
    wire signal_9968 ;
    wire signal_9969 ;
    wire signal_9970 ;
    wire signal_9971 ;
    wire signal_9972 ;
    wire signal_9973 ;
    wire signal_9974 ;
    wire signal_9975 ;
    wire signal_9976 ;
    wire signal_9977 ;
    wire signal_9978 ;
    wire signal_9979 ;
    wire signal_9980 ;
    wire signal_9981 ;
    wire signal_9982 ;
    wire signal_9983 ;
    wire signal_9984 ;
    wire signal_9985 ;
    wire signal_9986 ;
    wire signal_9987 ;
    wire signal_9988 ;
    wire signal_9989 ;
    wire signal_9990 ;
    wire signal_9991 ;
    wire signal_9992 ;
    wire signal_9993 ;
    wire signal_9994 ;
    wire signal_9995 ;
    wire signal_9996 ;
    wire signal_9997 ;
    wire signal_9998 ;
    wire signal_9999 ;
    wire signal_10000 ;
    wire signal_10001 ;
    wire signal_10002 ;
    wire signal_10003 ;
    wire signal_10004 ;
    wire signal_10005 ;
    wire signal_10006 ;
    wire signal_10007 ;
    wire signal_10008 ;
    wire signal_10009 ;
    wire signal_10010 ;
    wire signal_10011 ;
    wire signal_10012 ;
    wire signal_10013 ;
    wire signal_10014 ;
    wire signal_10015 ;
    wire signal_10016 ;
    wire signal_10017 ;
    wire signal_10018 ;
    wire signal_10019 ;
    wire signal_10020 ;
    wire signal_10021 ;
    wire signal_10022 ;
    wire signal_10023 ;
    wire signal_10024 ;
    wire signal_10025 ;
    wire signal_10026 ;
    wire signal_10027 ;
    wire signal_10028 ;
    wire signal_10029 ;
    wire signal_10030 ;
    wire signal_10031 ;
    wire signal_10032 ;
    wire signal_10033 ;
    wire signal_10034 ;
    wire signal_10035 ;
    wire signal_10036 ;
    wire signal_10037 ;
    wire signal_10038 ;
    wire signal_10039 ;
    wire signal_10040 ;
    wire signal_10041 ;
    wire signal_10042 ;
    wire signal_10043 ;
    wire signal_10044 ;
    wire signal_10045 ;
    wire signal_10046 ;
    wire signal_10047 ;
    wire signal_10048 ;
    wire signal_10049 ;
    wire signal_10050 ;
    wire signal_10051 ;
    wire signal_10052 ;
    wire signal_10053 ;
    wire signal_10054 ;
    wire signal_10055 ;
    wire signal_10056 ;
    wire signal_10057 ;
    wire signal_10058 ;
    wire signal_10059 ;
    wire signal_10060 ;
    wire signal_10061 ;
    wire signal_10062 ;
    wire signal_10063 ;
    wire signal_10064 ;
    wire signal_10065 ;
    wire signal_10066 ;
    wire signal_10067 ;
    wire signal_10068 ;
    wire signal_10069 ;
    wire signal_10070 ;
    wire signal_10071 ;
    wire signal_10072 ;
    wire signal_10073 ;
    wire signal_10074 ;
    wire signal_10075 ;
    wire signal_10076 ;
    wire signal_10077 ;
    wire signal_10078 ;
    wire signal_10079 ;
    wire signal_10080 ;
    wire signal_10081 ;
    wire signal_10082 ;
    wire signal_10083 ;
    wire signal_10084 ;
    wire signal_10085 ;
    wire signal_10086 ;
    wire signal_10087 ;
    wire signal_10088 ;
    wire signal_10089 ;
    wire signal_10090 ;
    wire signal_10091 ;
    wire signal_10092 ;
    wire signal_10093 ;
    wire signal_10094 ;
    wire signal_10095 ;
    wire signal_10096 ;
    wire signal_10097 ;
    wire signal_10098 ;
    wire signal_10099 ;
    wire signal_10100 ;
    wire signal_10101 ;
    wire signal_10102 ;
    wire signal_10103 ;
    wire signal_10104 ;
    wire signal_10105 ;
    wire signal_10106 ;
    wire signal_10107 ;
    wire signal_10108 ;
    wire signal_10109 ;
    wire signal_10110 ;
    wire signal_10111 ;
    wire signal_10112 ;
    wire signal_10113 ;
    wire signal_10114 ;
    wire signal_10115 ;
    wire signal_10116 ;
    wire signal_10117 ;
    wire signal_10118 ;
    wire signal_10119 ;
    wire signal_10120 ;
    wire signal_10121 ;
    wire signal_10122 ;
    wire signal_10123 ;
    wire signal_10124 ;
    wire signal_10125 ;
    wire signal_10126 ;
    wire signal_10127 ;
    wire signal_10128 ;
    wire signal_10129 ;
    wire signal_10130 ;
    wire signal_10131 ;
    wire signal_10132 ;
    wire signal_10133 ;
    wire signal_10134 ;
    wire signal_10135 ;
    wire signal_10136 ;
    wire signal_10137 ;
    wire signal_10138 ;
    wire signal_10139 ;
    wire signal_10140 ;
    wire signal_10141 ;
    wire signal_10142 ;
    wire signal_10143 ;
    wire signal_10144 ;
    wire signal_10145 ;
    wire signal_10146 ;
    wire signal_10147 ;
    wire signal_10148 ;
    wire signal_10149 ;
    wire signal_10150 ;
    wire signal_10151 ;
    wire signal_10152 ;
    wire signal_10153 ;
    wire signal_10154 ;
    wire signal_10155 ;
    wire signal_10156 ;
    wire signal_10157 ;
    wire signal_10158 ;
    wire signal_10159 ;
    wire signal_10160 ;
    wire signal_10161 ;
    wire signal_10162 ;
    wire signal_10163 ;
    wire signal_10164 ;
    wire signal_10165 ;
    wire signal_10166 ;
    wire signal_10167 ;
    wire signal_10168 ;
    wire signal_10169 ;
    wire signal_10170 ;
    wire signal_10171 ;
    wire signal_10172 ;
    wire signal_10173 ;
    wire signal_10174 ;
    wire signal_10175 ;
    wire signal_10176 ;
    wire signal_10177 ;
    wire signal_10178 ;
    wire signal_10179 ;
    wire signal_10180 ;
    wire signal_10181 ;
    wire signal_10182 ;
    wire signal_10183 ;
    wire signal_10184 ;
    wire signal_10185 ;
    wire signal_10186 ;
    wire signal_10187 ;
    wire signal_10188 ;
    wire signal_10189 ;
    wire signal_10190 ;
    wire signal_10191 ;
    wire signal_10192 ;
    wire signal_10193 ;
    wire signal_10194 ;
    wire signal_10195 ;
    wire signal_10196 ;
    wire signal_10197 ;
    wire signal_10198 ;
    wire signal_10199 ;
    wire signal_10200 ;
    wire signal_10201 ;
    wire signal_10202 ;
    wire signal_10203 ;
    wire signal_10204 ;
    wire signal_10205 ;
    wire signal_10206 ;
    wire signal_10207 ;
    wire signal_10208 ;
    wire signal_10209 ;
    wire signal_10210 ;
    wire signal_10211 ;
    wire signal_10212 ;
    wire signal_10213 ;
    wire signal_10214 ;
    wire signal_10215 ;
    wire signal_10216 ;
    wire signal_10217 ;
    wire signal_10218 ;
    wire signal_10219 ;
    wire signal_10220 ;
    wire signal_10221 ;
    wire signal_10222 ;
    wire signal_10223 ;
    wire signal_10224 ;
    wire signal_10225 ;
    wire signal_10226 ;
    wire signal_10227 ;
    wire signal_10228 ;
    wire signal_10229 ;
    wire signal_10230 ;
    wire signal_10231 ;
    wire signal_10232 ;
    wire signal_10233 ;
    wire signal_10234 ;
    wire signal_10235 ;
    wire signal_10236 ;
    wire signal_10237 ;
    wire signal_10238 ;
    wire signal_10239 ;
    wire signal_10240 ;
    wire signal_10241 ;
    wire signal_10242 ;
    wire signal_10243 ;
    wire signal_10244 ;
    wire signal_10245 ;
    wire signal_10246 ;
    wire signal_10247 ;
    wire signal_10248 ;
    wire signal_10249 ;
    wire signal_10250 ;
    wire signal_10251 ;
    wire signal_10252 ;
    wire signal_10253 ;
    wire signal_10254 ;
    wire signal_10255 ;
    wire signal_10256 ;
    wire signal_10257 ;
    wire signal_10258 ;
    wire signal_10259 ;
    wire signal_10260 ;
    wire signal_10261 ;
    wire signal_10262 ;
    wire signal_10263 ;
    wire signal_10264 ;
    wire signal_10265 ;
    wire signal_10266 ;
    wire signal_10267 ;
    wire signal_10268 ;
    wire signal_10269 ;
    wire signal_10270 ;
    wire signal_10271 ;
    wire signal_10272 ;
    wire signal_10273 ;
    wire signal_10274 ;
    wire signal_10275 ;
    wire signal_10276 ;
    wire signal_10277 ;
    wire signal_10278 ;
    wire signal_10279 ;
    wire signal_10280 ;
    wire signal_10281 ;
    wire signal_10282 ;
    wire signal_10283 ;
    wire signal_10284 ;
    wire signal_10285 ;
    wire signal_10286 ;
    wire signal_10287 ;
    wire signal_10288 ;
    wire signal_10289 ;
    wire signal_10290 ;
    wire signal_10291 ;
    wire signal_10292 ;
    wire signal_10293 ;
    wire signal_10294 ;
    wire signal_10295 ;
    wire signal_10296 ;
    wire signal_10297 ;
    wire signal_10298 ;
    wire signal_10299 ;
    wire signal_10300 ;
    wire signal_10301 ;
    wire signal_10302 ;
    wire signal_10303 ;
    wire signal_10304 ;
    wire signal_10305 ;
    wire signal_10306 ;
    wire signal_10307 ;
    wire signal_10308 ;
    wire signal_10309 ;
    wire signal_10310 ;
    wire signal_10311 ;
    wire signal_10312 ;
    wire signal_10313 ;
    wire signal_10314 ;
    wire signal_10315 ;
    wire signal_10316 ;
    wire signal_10317 ;
    wire signal_10318 ;
    wire signal_10319 ;
    wire signal_10320 ;
    wire signal_10321 ;
    wire signal_10322 ;
    wire signal_10323 ;
    wire signal_10324 ;
    wire signal_10325 ;
    wire signal_10326 ;
    wire signal_10327 ;
    wire signal_10328 ;
    wire signal_10329 ;
    wire signal_10330 ;
    wire signal_10331 ;
    wire signal_10332 ;
    wire signal_10333 ;
    wire signal_10334 ;
    wire signal_10335 ;
    wire signal_10336 ;
    wire signal_10337 ;
    wire signal_10338 ;
    wire signal_10339 ;
    wire signal_10340 ;
    wire signal_10341 ;
    wire signal_10342 ;
    wire signal_10343 ;
    wire signal_10344 ;
    wire signal_10345 ;
    wire signal_10346 ;
    wire signal_10347 ;
    wire signal_10348 ;
    wire signal_10349 ;
    wire signal_10350 ;
    wire signal_10351 ;
    wire signal_10352 ;
    wire signal_10353 ;
    wire signal_10354 ;
    wire signal_10355 ;
    wire signal_10356 ;
    wire signal_10357 ;
    wire signal_10358 ;
    wire signal_10359 ;
    wire signal_10360 ;
    wire signal_10361 ;
    wire signal_10362 ;
    wire signal_10363 ;
    wire signal_10364 ;
    wire signal_10365 ;
    wire signal_10366 ;
    wire signal_10367 ;
    wire signal_10368 ;
    wire signal_10369 ;
    wire signal_10370 ;
    wire signal_10371 ;
    wire signal_10372 ;
    wire signal_10373 ;
    wire signal_10374 ;
    wire signal_10375 ;
    wire signal_10376 ;
    wire signal_10377 ;
    wire signal_10378 ;
    wire signal_10379 ;
    wire signal_10380 ;
    wire signal_10381 ;
    wire signal_10382 ;
    wire signal_10383 ;
    wire signal_10384 ;
    wire signal_10385 ;
    wire signal_10386 ;
    wire signal_10387 ;
    wire signal_10388 ;
    wire signal_10389 ;
    wire signal_10390 ;
    wire signal_10391 ;
    wire signal_10392 ;
    wire signal_10393 ;
    wire signal_10394 ;
    wire signal_10395 ;
    wire signal_10396 ;
    wire signal_10397 ;
    wire signal_10398 ;
    wire signal_10399 ;
    wire signal_10400 ;
    wire signal_10401 ;
    wire signal_10402 ;
    wire signal_10403 ;
    wire signal_10404 ;
    wire signal_10405 ;
    wire signal_10406 ;
    wire signal_10407 ;
    wire signal_10408 ;
    wire signal_10409 ;
    wire signal_10410 ;
    wire signal_10411 ;
    wire signal_10412 ;
    wire signal_10413 ;
    wire signal_10414 ;
    wire signal_10415 ;
    wire signal_10416 ;
    wire signal_10417 ;
    wire signal_10418 ;
    wire signal_10419 ;
    wire signal_10420 ;
    wire signal_10421 ;
    wire signal_10422 ;
    wire signal_10423 ;
    wire signal_10424 ;
    wire signal_10425 ;
    wire signal_10426 ;
    wire signal_10427 ;
    wire signal_10428 ;
    wire signal_10429 ;
    wire signal_10430 ;
    wire signal_10431 ;
    wire signal_10432 ;
    wire signal_10433 ;
    wire signal_10434 ;
    wire signal_10435 ;
    wire signal_10436 ;
    wire signal_10437 ;
    wire signal_10438 ;
    wire signal_10439 ;
    wire signal_10440 ;
    wire signal_10441 ;
    wire signal_10442 ;
    wire signal_10443 ;
    wire signal_10444 ;
    wire signal_10445 ;
    wire signal_10446 ;
    wire signal_10447 ;
    wire signal_10448 ;
    wire signal_10449 ;
    wire signal_10450 ;
    wire signal_10451 ;
    wire signal_10452 ;
    wire signal_10453 ;
    wire signal_10454 ;
    wire signal_10455 ;
    wire signal_10456 ;
    wire signal_10457 ;
    wire signal_10458 ;
    wire signal_10459 ;
    wire signal_10460 ;
    wire signal_10461 ;
    wire signal_10462 ;
    wire signal_10463 ;
    wire signal_10464 ;
    wire signal_10465 ;
    wire signal_10466 ;
    wire signal_10467 ;
    wire signal_10468 ;
    wire signal_10469 ;
    wire signal_10470 ;
    wire signal_10471 ;
    wire signal_10472 ;
    wire signal_10473 ;
    wire signal_10474 ;
    wire signal_10475 ;
    wire signal_10476 ;
    wire signal_10477 ;
    wire signal_10478 ;
    wire signal_10479 ;
    wire signal_10480 ;
    wire signal_10481 ;
    wire signal_10482 ;
    wire signal_10483 ;
    wire signal_10484 ;
    wire signal_10485 ;
    wire signal_10486 ;
    wire signal_10487 ;
    wire signal_10488 ;
    wire signal_10489 ;
    wire signal_10490 ;
    wire signal_10491 ;
    wire signal_10492 ;
    wire signal_10493 ;
    wire signal_10494 ;
    wire signal_10495 ;
    wire signal_10496 ;
    wire signal_10497 ;
    wire signal_10498 ;
    wire signal_10499 ;
    wire signal_10500 ;
    wire signal_10501 ;
    wire signal_10502 ;
    wire signal_10503 ;
    wire signal_10504 ;
    wire signal_10505 ;
    wire signal_10506 ;
    wire signal_10507 ;
    wire signal_10508 ;
    wire signal_10509 ;
    wire signal_10510 ;
    wire signal_10511 ;
    wire signal_10512 ;
    wire signal_10513 ;
    wire signal_10514 ;
    wire signal_10515 ;
    wire signal_10516 ;
    wire signal_10517 ;
    wire signal_10518 ;
    wire signal_10519 ;
    wire signal_10520 ;
    wire signal_10521 ;
    wire signal_10522 ;
    wire signal_10523 ;
    wire signal_10524 ;
    wire signal_10525 ;
    wire signal_10526 ;
    wire signal_10527 ;
    wire signal_10528 ;
    wire signal_10529 ;
    wire signal_10530 ;
    wire signal_10531 ;
    wire signal_10532 ;
    wire signal_10533 ;
    wire signal_10534 ;
    wire signal_10535 ;
    wire signal_10536 ;
    wire signal_10537 ;
    wire signal_10538 ;
    wire signal_10539 ;
    wire signal_10540 ;
    wire signal_10541 ;
    wire signal_10542 ;
    wire signal_10543 ;
    wire signal_10544 ;
    wire signal_10545 ;
    wire signal_10546 ;
    wire signal_10547 ;
    wire signal_10548 ;
    wire signal_10549 ;
    wire signal_10550 ;
    wire signal_10551 ;
    wire signal_10552 ;
    wire signal_10553 ;
    wire signal_10554 ;
    wire signal_10555 ;
    wire signal_10556 ;
    wire signal_10557 ;
    wire signal_10558 ;
    wire signal_10559 ;
    wire signal_10560 ;
    wire signal_10561 ;
    wire signal_10562 ;
    wire signal_10563 ;
    wire signal_10564 ;
    wire signal_10565 ;
    wire signal_10566 ;
    wire signal_10567 ;
    wire signal_10568 ;
    wire signal_10569 ;
    wire signal_10570 ;
    wire signal_10571 ;
    wire signal_10572 ;
    wire signal_10573 ;
    wire signal_10574 ;
    wire signal_10575 ;
    wire signal_10576 ;
    wire signal_10577 ;
    wire signal_10578 ;
    wire signal_10579 ;
    wire signal_10580 ;
    wire signal_10581 ;
    wire signal_10582 ;
    wire signal_10583 ;
    wire signal_10584 ;
    wire signal_10585 ;
    wire signal_10586 ;
    wire signal_10587 ;
    wire signal_10588 ;
    wire signal_10589 ;
    wire signal_10590 ;
    wire signal_10591 ;
    wire signal_10592 ;
    wire signal_10593 ;
    wire signal_10594 ;
    wire signal_10595 ;
    wire signal_10596 ;
    wire signal_10597 ;
    wire signal_10598 ;
    wire signal_10599 ;
    wire signal_10600 ;
    wire signal_10601 ;
    wire signal_10602 ;
    wire signal_10603 ;
    wire signal_10604 ;
    wire signal_10605 ;
    wire signal_10606 ;
    wire signal_10607 ;
    wire signal_10608 ;
    wire signal_10609 ;
    wire signal_10610 ;
    wire signal_10611 ;
    wire signal_10612 ;
    wire signal_10613 ;
    wire signal_10614 ;
    wire signal_10615 ;
    wire signal_10616 ;
    wire signal_10617 ;
    wire signal_10618 ;
    wire signal_10619 ;
    wire signal_10620 ;
    wire signal_10621 ;
    wire signal_10622 ;
    wire signal_10623 ;
    wire signal_10624 ;
    wire signal_10625 ;
    wire signal_10626 ;
    wire signal_10627 ;
    wire signal_10628 ;
    wire signal_10629 ;
    wire signal_10630 ;
    wire signal_10631 ;
    wire signal_10632 ;
    wire signal_10633 ;
    wire signal_10634 ;
    wire signal_10635 ;
    wire signal_10636 ;
    wire signal_10637 ;
    wire signal_10638 ;
    wire signal_10639 ;
    wire signal_10640 ;
    wire signal_10641 ;
    wire signal_10642 ;
    wire signal_10643 ;
    wire signal_10644 ;
    wire signal_10645 ;
    wire signal_10646 ;
    wire signal_10647 ;
    wire signal_10648 ;
    wire signal_10649 ;
    wire signal_10650 ;
    wire signal_10651 ;
    wire signal_10652 ;
    wire signal_10653 ;
    wire signal_10654 ;
    wire signal_10655 ;
    wire signal_10656 ;
    wire signal_10657 ;
    wire signal_10658 ;
    wire signal_10659 ;
    wire signal_10660 ;
    wire signal_10661 ;
    wire signal_10662 ;
    wire signal_10663 ;
    wire signal_10664 ;
    wire signal_10665 ;
    wire signal_10666 ;
    wire signal_10667 ;
    wire signal_10668 ;
    wire signal_10669 ;
    wire signal_10670 ;
    wire signal_10671 ;
    wire signal_10672 ;
    wire signal_10673 ;
    wire signal_10674 ;
    wire signal_10675 ;
    wire signal_10676 ;
    wire signal_10677 ;
    wire signal_10678 ;
    wire signal_10679 ;
    wire signal_10680 ;
    wire signal_10681 ;
    wire signal_10682 ;
    wire signal_10683 ;
    wire signal_10684 ;
    wire signal_10685 ;
    wire signal_10686 ;
    wire signal_10687 ;
    wire signal_10688 ;
    wire signal_10689 ;
    wire signal_10690 ;
    wire signal_10691 ;
    wire signal_10692 ;
    wire signal_10693 ;
    wire signal_10694 ;
    wire signal_10695 ;
    wire signal_10696 ;
    wire signal_10697 ;
    wire signal_10698 ;
    wire signal_10699 ;
    wire signal_10700 ;
    wire signal_10701 ;
    wire signal_10702 ;
    wire signal_10703 ;
    wire signal_10704 ;
    wire signal_10705 ;
    wire signal_10706 ;
    wire signal_10707 ;
    wire signal_10708 ;
    wire signal_10709 ;
    wire signal_10710 ;
    wire signal_10711 ;
    wire signal_10712 ;
    wire signal_10713 ;
    wire signal_10714 ;
    wire signal_10715 ;
    wire signal_10716 ;
    wire signal_10717 ;
    wire signal_10718 ;
    wire signal_10719 ;
    wire signal_10720 ;
    wire signal_10721 ;
    wire signal_10722 ;
    wire signal_10723 ;
    wire signal_10724 ;
    wire signal_10725 ;
    wire signal_10726 ;
    wire signal_10727 ;
    wire signal_10728 ;
    wire signal_10729 ;
    wire signal_10730 ;
    wire signal_10731 ;
    wire signal_10732 ;
    wire signal_10733 ;
    wire signal_10734 ;
    wire signal_10735 ;
    wire signal_10736 ;
    wire signal_10737 ;
    wire signal_10738 ;
    wire signal_10739 ;
    wire signal_10740 ;
    wire signal_10741 ;
    wire signal_10742 ;
    wire signal_10743 ;
    wire signal_10744 ;
    wire signal_10745 ;
    wire signal_10746 ;
    wire signal_10747 ;
    wire signal_10748 ;
    wire signal_10749 ;
    wire signal_10750 ;
    wire signal_10751 ;
    wire signal_10752 ;
    wire signal_10753 ;
    wire signal_10754 ;
    wire signal_10755 ;
    wire signal_10756 ;
    wire signal_10757 ;
    wire signal_10758 ;
    wire signal_10759 ;
    wire signal_10760 ;
    wire signal_10761 ;
    wire signal_10762 ;
    wire signal_10763 ;
    wire signal_10764 ;
    wire signal_10765 ;
    wire signal_10766 ;
    wire signal_10767 ;
    wire signal_10768 ;
    wire signal_10769 ;
    wire signal_10770 ;
    wire signal_10771 ;
    wire signal_10772 ;
    wire signal_10773 ;
    wire signal_10774 ;
    wire signal_10775 ;
    wire signal_10776 ;
    wire signal_10777 ;
    wire signal_10778 ;
    wire signal_10779 ;
    wire signal_10780 ;
    wire signal_10781 ;
    wire signal_10782 ;
    wire signal_10783 ;
    wire signal_10784 ;
    wire signal_10785 ;
    wire signal_10786 ;
    wire signal_10787 ;
    wire signal_10788 ;
    wire signal_10789 ;
    wire signal_10790 ;
    wire signal_10791 ;
    wire signal_10792 ;
    wire signal_10793 ;
    wire signal_10794 ;
    wire signal_10795 ;
    wire signal_10796 ;
    wire signal_10797 ;
    wire signal_10798 ;
    wire signal_10799 ;
    wire signal_10800 ;
    wire signal_10801 ;
    wire signal_10802 ;
    wire signal_10803 ;
    wire signal_10804 ;
    wire signal_10805 ;
    wire signal_10806 ;
    wire signal_10807 ;
    wire signal_10808 ;
    wire signal_10809 ;
    wire signal_10810 ;
    wire signal_10811 ;
    wire signal_10812 ;
    wire signal_10813 ;
    wire signal_10814 ;
    wire signal_10815 ;
    wire signal_10816 ;
    wire signal_10817 ;
    wire signal_10818 ;
    wire signal_10819 ;
    wire signal_10820 ;
    wire signal_10821 ;
    wire signal_10822 ;
    wire signal_10823 ;
    wire signal_10824 ;
    wire signal_10825 ;
    wire signal_10826 ;
    wire signal_10827 ;
    wire signal_10828 ;
    wire signal_10829 ;
    wire signal_10830 ;
    wire signal_10831 ;
    wire signal_10832 ;
    wire signal_10833 ;
    wire signal_10834 ;
    wire signal_10835 ;
    wire signal_10836 ;
    wire signal_10837 ;
    wire signal_10838 ;
    wire signal_10839 ;
    wire signal_10840 ;
    wire signal_10841 ;
    wire signal_10842 ;
    wire signal_10843 ;
    wire signal_10844 ;
    wire signal_10845 ;
    wire signal_10846 ;
    wire signal_10847 ;
    wire signal_10848 ;
    wire signal_10849 ;
    wire signal_10850 ;
    wire signal_10851 ;
    wire signal_10852 ;
    wire signal_10853 ;
    wire signal_10854 ;
    wire signal_10855 ;
    wire signal_10856 ;
    wire signal_10857 ;
    wire signal_10858 ;
    wire signal_10859 ;
    wire signal_10860 ;
    wire signal_10861 ;
    wire signal_10862 ;
    wire signal_10863 ;
    wire signal_10864 ;
    wire signal_10865 ;
    wire signal_10866 ;
    wire signal_10867 ;
    wire signal_10868 ;
    wire signal_10869 ;
    wire signal_10870 ;
    wire signal_10871 ;
    wire signal_10872 ;
    wire signal_10873 ;
    wire signal_10874 ;
    wire signal_10875 ;
    wire signal_10876 ;
    wire signal_10877 ;
    wire signal_10878 ;
    wire signal_10879 ;
    wire signal_10880 ;
    wire signal_10881 ;
    wire signal_10882 ;
    wire signal_10883 ;
    wire signal_10884 ;
    wire signal_10885 ;
    wire signal_10886 ;
    wire signal_10887 ;
    wire signal_10888 ;
    wire signal_10889 ;
    wire signal_10890 ;
    wire signal_10891 ;
    wire signal_10892 ;
    wire signal_10893 ;
    wire signal_10894 ;
    wire signal_10895 ;
    wire signal_10896 ;
    wire signal_10897 ;
    wire signal_10898 ;
    wire signal_10899 ;
    wire signal_10900 ;
    wire signal_10901 ;
    wire signal_10902 ;
    wire signal_10903 ;
    wire signal_10904 ;
    wire signal_10905 ;
    wire signal_10906 ;
    wire signal_10907 ;
    wire signal_10908 ;
    wire signal_10909 ;
    wire signal_10910 ;
    wire signal_10911 ;
    wire signal_10912 ;
    wire signal_10913 ;
    wire signal_10914 ;
    wire signal_10915 ;
    wire signal_10916 ;
    wire signal_10917 ;
    wire signal_10918 ;
    wire signal_10919 ;
    wire signal_10920 ;
    wire signal_10921 ;
    wire signal_10922 ;
    wire signal_10923 ;
    wire signal_10924 ;
    wire signal_10925 ;
    wire signal_10926 ;
    wire signal_10927 ;
    wire signal_10928 ;
    wire signal_10929 ;
    wire signal_10930 ;
    wire signal_10931 ;
    wire signal_10932 ;
    wire signal_10933 ;
    wire signal_10934 ;
    wire signal_10935 ;
    wire signal_10936 ;
    wire signal_10937 ;
    wire signal_10938 ;
    wire signal_10939 ;
    wire signal_10940 ;
    wire signal_10941 ;
    wire signal_10942 ;
    wire signal_10943 ;
    wire signal_10944 ;
    wire signal_10945 ;
    wire signal_10946 ;
    wire signal_10947 ;
    wire signal_10948 ;
    wire signal_10949 ;
    wire signal_10950 ;
    wire signal_10951 ;
    wire signal_10952 ;
    wire signal_10953 ;
    wire signal_10954 ;
    wire signal_10955 ;
    wire signal_10956 ;
    wire signal_10957 ;
    wire signal_10958 ;
    wire signal_10959 ;
    wire signal_10960 ;
    wire signal_10961 ;
    wire signal_10962 ;
    wire signal_10963 ;
    wire signal_10964 ;
    wire signal_10965 ;
    wire signal_10966 ;
    wire signal_10967 ;
    wire signal_10968 ;
    wire signal_10969 ;
    wire signal_10970 ;
    wire signal_10971 ;
    wire signal_10972 ;
    wire signal_10973 ;
    wire signal_10974 ;
    wire signal_10975 ;
    wire signal_10976 ;
    wire signal_10977 ;
    wire signal_10978 ;
    wire signal_10979 ;
    wire signal_10980 ;
    wire signal_10981 ;
    wire signal_10982 ;
    wire signal_10983 ;
    wire signal_10984 ;
    wire signal_10985 ;
    wire signal_10986 ;
    wire signal_10987 ;
    wire signal_10988 ;
    wire signal_10989 ;
    wire signal_10990 ;
    wire signal_10991 ;
    wire signal_10992 ;
    wire signal_10993 ;
    wire signal_10994 ;
    wire signal_10995 ;
    wire signal_10996 ;
    wire signal_10997 ;
    wire signal_10998 ;
    wire signal_10999 ;
    wire signal_11000 ;
    wire signal_11001 ;
    wire signal_11002 ;
    wire signal_11003 ;
    wire signal_11004 ;
    wire signal_11005 ;
    wire signal_11006 ;
    wire signal_11007 ;
    wire signal_11008 ;
    wire signal_11009 ;
    wire signal_11010 ;
    wire signal_11011 ;
    wire signal_11012 ;
    wire signal_11013 ;
    wire signal_11014 ;
    wire signal_11015 ;
    wire signal_11016 ;
    wire signal_11017 ;
    wire signal_11018 ;
    wire signal_11019 ;
    wire signal_11020 ;
    wire signal_11021 ;
    wire signal_11022 ;
    wire signal_11023 ;
    wire signal_11024 ;
    wire signal_11025 ;
    wire signal_11026 ;
    wire signal_11027 ;
    wire signal_11028 ;
    wire signal_11029 ;
    wire signal_11030 ;
    wire signal_11031 ;
    wire signal_11032 ;
    wire signal_11033 ;
    wire signal_11034 ;
    wire signal_11035 ;
    wire signal_11036 ;
    wire signal_11037 ;
    wire signal_11038 ;
    wire signal_11039 ;
    wire signal_11040 ;
    wire signal_11041 ;
    wire signal_11042 ;
    wire signal_11043 ;
    wire signal_11044 ;
    wire signal_11045 ;
    wire signal_11046 ;
    wire signal_11047 ;
    wire signal_11048 ;
    wire signal_11049 ;
    wire signal_11050 ;
    wire signal_11051 ;
    wire signal_11052 ;
    wire signal_11053 ;
    wire signal_11054 ;
    wire signal_11055 ;
    wire signal_11056 ;
    wire signal_11057 ;
    wire signal_11058 ;
    wire signal_11059 ;
    wire signal_11060 ;
    wire signal_11061 ;
    wire signal_11062 ;
    wire signal_11063 ;
    wire signal_11064 ;
    wire signal_11065 ;
    wire signal_11066 ;
    wire signal_11067 ;
    wire signal_11068 ;
    wire signal_11069 ;
    wire signal_11070 ;
    wire signal_11071 ;
    wire signal_11072 ;
    wire signal_11073 ;
    wire signal_11074 ;
    wire signal_11075 ;
    wire signal_11076 ;
    wire signal_11077 ;
    wire signal_11078 ;
    wire signal_11079 ;
    wire signal_11080 ;
    wire signal_11081 ;
    wire signal_11082 ;
    wire signal_11083 ;
    wire signal_11084 ;
    wire signal_11085 ;
    wire signal_11086 ;
    wire signal_11087 ;
    wire signal_11088 ;
    wire signal_11089 ;
    wire signal_11090 ;
    wire signal_11091 ;
    wire signal_11092 ;
    wire signal_11093 ;
    wire signal_11094 ;
    wire signal_11095 ;
    wire signal_11096 ;
    wire signal_11097 ;
    wire signal_11098 ;
    wire signal_11099 ;
    wire signal_11100 ;
    wire signal_11101 ;
    wire signal_11102 ;
    wire signal_11103 ;
    wire signal_11104 ;
    wire signal_11105 ;
    wire signal_11106 ;
    wire signal_11107 ;
    wire signal_11108 ;
    wire signal_11109 ;
    wire signal_11110 ;
    wire signal_11111 ;
    wire signal_11112 ;
    wire signal_11113 ;
    wire signal_11114 ;
    wire signal_11115 ;
    wire signal_11116 ;
    wire signal_11117 ;
    wire signal_11118 ;
    wire signal_11119 ;
    wire signal_11120 ;
    wire signal_11121 ;
    wire signal_11122 ;
    wire signal_11123 ;
    wire signal_11124 ;
    wire signal_11125 ;
    wire signal_11126 ;
    wire signal_11127 ;
    wire signal_11128 ;
    wire signal_11129 ;
    wire signal_11130 ;
    wire signal_11131 ;
    wire signal_11132 ;
    wire signal_11133 ;
    wire signal_11134 ;
    wire signal_11135 ;
    wire signal_11136 ;
    wire signal_11137 ;
    wire signal_11138 ;
    wire signal_11139 ;
    wire signal_11140 ;
    wire signal_11141 ;
    wire signal_11142 ;
    wire signal_11143 ;
    wire signal_11144 ;
    wire signal_11145 ;
    wire signal_11146 ;
    wire signal_11147 ;
    wire signal_11148 ;
    wire signal_11149 ;
    wire signal_11150 ;
    wire signal_11151 ;
    wire signal_11152 ;
    wire signal_11153 ;
    wire signal_11154 ;
    wire signal_11155 ;
    wire signal_11156 ;
    wire signal_11157 ;
    wire signal_11158 ;
    wire signal_11159 ;
    wire signal_11160 ;
    wire signal_11161 ;
    wire signal_11162 ;
    wire signal_11163 ;
    wire signal_11164 ;
    wire signal_11165 ;
    wire signal_11166 ;
    wire signal_11167 ;
    wire signal_11168 ;
    wire signal_11169 ;
    wire signal_11170 ;
    wire signal_11171 ;
    wire signal_11172 ;
    wire signal_11173 ;
    wire signal_11174 ;
    wire signal_11175 ;
    wire signal_11176 ;
    wire signal_11177 ;
    wire signal_11178 ;
    wire signal_11179 ;
    wire signal_11180 ;
    wire signal_11181 ;
    wire signal_11182 ;
    wire signal_11183 ;
    wire signal_11184 ;
    wire signal_11185 ;
    wire signal_11186 ;
    wire signal_11187 ;
    wire signal_11188 ;
    wire signal_11189 ;
    wire signal_11190 ;
    wire signal_11191 ;
    wire signal_11192 ;
    wire signal_11193 ;
    wire signal_11194 ;
    wire signal_11195 ;
    wire signal_11196 ;
    wire signal_11197 ;
    wire signal_11198 ;
    wire signal_11199 ;
    wire signal_11200 ;
    wire signal_11201 ;
    wire signal_11202 ;
    wire signal_11203 ;
    wire signal_11204 ;
    wire signal_11205 ;
    wire signal_11206 ;
    wire signal_11207 ;
    wire signal_11208 ;
    wire signal_11209 ;
    wire signal_11210 ;
    wire signal_11211 ;
    wire signal_11212 ;
    wire signal_11213 ;
    wire signal_11214 ;
    wire signal_11215 ;
    wire signal_11216 ;
    wire signal_11217 ;
    wire signal_11218 ;
    wire signal_11219 ;
    wire signal_11220 ;
    wire signal_11221 ;
    wire signal_11222 ;
    wire signal_11223 ;
    wire signal_11224 ;
    wire signal_11225 ;
    wire signal_11226 ;
    wire signal_11227 ;
    wire signal_11228 ;
    wire signal_11229 ;
    wire signal_11230 ;
    wire signal_11231 ;
    wire signal_11232 ;
    wire signal_11233 ;
    wire signal_11234 ;
    wire signal_11235 ;
    wire signal_11236 ;
    wire signal_11237 ;
    wire signal_11238 ;
    wire signal_11239 ;
    wire signal_11240 ;
    wire signal_11241 ;
    wire signal_11242 ;
    wire signal_11243 ;
    wire signal_11244 ;
    wire signal_11245 ;
    wire signal_11246 ;
    wire signal_11247 ;
    wire signal_11248 ;
    wire signal_11249 ;
    wire signal_11250 ;
    wire signal_11251 ;
    wire signal_11252 ;
    wire signal_11253 ;
    wire signal_11254 ;
    wire signal_11255 ;
    wire signal_11256 ;
    wire signal_11257 ;
    wire signal_11258 ;
    wire signal_11259 ;
    wire signal_11260 ;
    wire signal_11261 ;
    wire signal_11262 ;
    wire signal_11263 ;
    wire signal_11264 ;
    wire signal_11265 ;
    wire signal_11266 ;
    wire signal_11267 ;
    wire signal_11268 ;
    wire signal_11269 ;
    wire signal_11270 ;
    wire signal_11271 ;
    wire signal_11272 ;
    wire signal_11273 ;
    wire signal_11274 ;
    wire signal_11275 ;
    wire signal_11276 ;
    wire signal_11277 ;
    wire signal_11278 ;
    wire signal_11279 ;
    wire signal_11280 ;
    wire signal_11281 ;
    wire signal_11282 ;
    wire signal_11283 ;
    wire signal_11284 ;
    wire signal_11285 ;
    wire signal_11286 ;
    wire signal_11287 ;
    wire signal_11288 ;
    wire signal_11289 ;
    wire signal_11290 ;
    wire signal_11291 ;
    wire signal_11292 ;
    wire signal_11293 ;
    wire signal_11294 ;
    wire signal_11295 ;
    wire signal_11296 ;
    wire signal_11297 ;
    wire signal_11298 ;
    wire signal_11299 ;
    wire signal_11300 ;
    wire signal_11301 ;
    wire signal_11302 ;
    wire signal_11303 ;
    wire signal_11304 ;
    wire signal_11305 ;
    wire signal_11306 ;
    wire signal_11307 ;
    wire signal_11308 ;
    wire signal_11309 ;
    wire signal_11310 ;
    wire signal_11311 ;
    wire signal_11312 ;
    wire signal_11313 ;
    wire signal_11314 ;
    wire signal_11315 ;
    wire signal_11316 ;
    wire signal_11317 ;
    wire signal_11318 ;
    wire signal_11319 ;
    wire signal_11320 ;
    wire signal_11321 ;
    wire signal_11322 ;
    wire signal_11323 ;
    wire signal_11324 ;
    wire signal_11325 ;
    wire signal_11326 ;
    wire signal_11327 ;
    wire signal_11328 ;
    wire signal_11329 ;
    wire signal_11330 ;
    wire signal_11331 ;
    wire signal_11332 ;
    wire signal_11333 ;
    wire signal_11334 ;
    wire signal_11335 ;
    wire signal_11336 ;
    wire signal_11337 ;
    wire signal_11338 ;
    wire signal_11339 ;
    wire signal_11340 ;
    wire signal_11341 ;
    wire signal_11342 ;
    wire signal_11343 ;
    wire signal_11344 ;
    wire signal_11345 ;
    wire signal_11346 ;
    wire signal_11347 ;
    wire signal_11348 ;
    wire signal_11349 ;
    wire signal_11350 ;
    wire signal_11351 ;
    wire signal_11352 ;
    wire signal_11353 ;
    wire signal_11354 ;
    wire signal_11355 ;
    wire signal_11356 ;
    wire signal_11357 ;
    wire signal_11358 ;
    wire signal_11359 ;
    wire signal_11360 ;
    wire signal_11361 ;
    wire signal_11362 ;
    wire signal_11363 ;
    wire signal_11364 ;
    wire signal_11365 ;
    wire signal_11366 ;
    wire signal_11367 ;
    wire signal_11368 ;
    wire signal_11369 ;
    wire signal_11370 ;
    wire signal_11371 ;
    wire signal_11372 ;
    wire signal_11373 ;
    wire signal_11374 ;
    wire signal_11375 ;
    wire signal_11376 ;
    wire signal_11377 ;
    wire signal_11378 ;
    wire signal_11379 ;
    wire signal_11380 ;
    wire signal_11381 ;
    wire signal_11382 ;
    wire signal_11383 ;
    wire signal_11384 ;
    wire signal_11385 ;
    wire signal_11386 ;
    wire signal_11387 ;
    wire signal_11388 ;
    wire signal_11389 ;
    wire signal_11390 ;
    wire signal_11391 ;
    wire signal_11392 ;
    wire signal_11393 ;
    wire signal_11394 ;
    wire signal_11395 ;
    wire signal_11396 ;
    wire signal_11397 ;
    wire signal_11398 ;
    wire signal_11399 ;
    wire signal_11400 ;
    wire signal_11401 ;
    wire signal_11402 ;
    wire signal_11403 ;
    wire signal_11404 ;
    wire signal_11405 ;
    wire signal_11406 ;
    wire signal_11407 ;
    wire signal_11408 ;
    wire signal_11409 ;
    wire signal_11410 ;
    wire signal_11411 ;
    wire signal_11412 ;
    wire signal_11413 ;
    wire signal_11414 ;
    wire signal_11415 ;
    wire signal_11416 ;
    wire signal_11417 ;
    wire signal_11418 ;
    wire signal_11419 ;
    wire signal_11420 ;
    wire signal_11421 ;
    wire signal_11422 ;
    wire signal_11423 ;
    wire signal_11424 ;
    wire signal_11425 ;
    wire signal_11426 ;
    wire signal_11427 ;
    wire signal_11428 ;
    wire signal_11429 ;
    wire signal_11430 ;
    wire signal_11431 ;
    wire signal_11432 ;
    wire signal_11433 ;
    wire signal_11434 ;
    wire signal_11435 ;
    wire signal_11436 ;
    wire signal_11437 ;
    wire signal_11438 ;
    wire signal_11439 ;
    wire signal_11440 ;
    wire signal_11441 ;
    wire signal_11442 ;
    wire signal_11443 ;
    wire signal_11444 ;
    wire signal_11445 ;
    wire signal_11446 ;
    wire signal_11447 ;
    wire signal_11448 ;
    wire signal_11449 ;
    wire signal_11450 ;
    wire signal_11451 ;
    wire signal_11452 ;
    wire signal_11453 ;
    wire signal_11454 ;
    wire signal_11455 ;
    wire signal_11456 ;
    wire signal_11457 ;
    wire signal_11458 ;
    wire signal_11459 ;
    wire signal_11460 ;
    wire signal_11461 ;
    wire signal_11462 ;
    wire signal_11463 ;
    wire signal_11464 ;
    wire signal_11465 ;
    wire signal_11466 ;
    wire signal_11467 ;
    wire signal_11468 ;
    wire signal_11469 ;
    wire signal_11470 ;
    wire signal_11471 ;
    wire signal_11472 ;
    wire signal_11473 ;
    wire signal_11474 ;
    wire signal_11475 ;
    wire signal_11476 ;
    wire signal_11477 ;
    wire signal_11478 ;
    wire signal_11479 ;
    wire signal_11480 ;
    wire signal_11481 ;
    wire signal_11482 ;
    wire signal_11483 ;
    wire signal_11484 ;
    wire signal_11485 ;
    wire signal_11486 ;
    wire signal_11487 ;
    wire signal_11488 ;
    wire signal_11489 ;
    wire signal_11490 ;
    wire signal_11491 ;
    wire signal_11492 ;
    wire signal_11493 ;
    wire signal_11494 ;
    wire signal_11495 ;
    wire signal_11496 ;
    wire signal_11497 ;
    wire signal_11498 ;
    wire signal_11499 ;
    wire signal_11500 ;
    wire signal_11501 ;
    wire signal_11502 ;
    wire signal_11503 ;
    wire signal_11504 ;
    wire signal_11505 ;
    wire signal_11506 ;
    wire signal_11507 ;
    wire signal_11508 ;
    wire signal_11509 ;
    wire signal_11510 ;
    wire signal_11511 ;
    wire signal_11512 ;
    wire signal_11513 ;
    wire signal_11514 ;
    wire signal_11515 ;
    wire signal_11516 ;
    wire signal_11517 ;
    wire signal_11518 ;
    wire signal_11519 ;
    wire signal_11520 ;
    wire signal_11521 ;
    wire signal_11522 ;
    wire signal_11523 ;
    wire signal_11524 ;
    wire signal_11525 ;
    wire signal_11526 ;
    wire signal_11527 ;
    wire signal_11528 ;
    wire signal_11529 ;
    wire signal_11530 ;
    wire signal_11531 ;
    wire signal_11532 ;
    wire signal_11533 ;
    wire signal_11534 ;
    wire signal_11535 ;
    wire signal_11536 ;
    wire signal_11537 ;
    wire signal_11538 ;
    wire signal_11539 ;
    wire signal_11540 ;
    wire signal_11541 ;
    wire signal_11542 ;
    wire signal_11543 ;
    wire signal_11544 ;
    wire signal_11545 ;
    wire signal_11546 ;
    wire signal_11547 ;
    wire signal_11548 ;
    wire signal_11549 ;
    wire signal_11550 ;
    wire signal_11551 ;
    wire signal_11552 ;
    wire signal_11553 ;
    wire signal_11554 ;
    wire signal_11555 ;
    wire signal_11556 ;
    wire signal_11557 ;
    wire signal_11558 ;
    wire signal_11559 ;
    wire signal_11560 ;
    wire signal_11561 ;
    wire signal_11562 ;
    wire signal_11563 ;
    wire signal_11564 ;
    wire signal_11565 ;
    wire signal_11566 ;
    wire signal_11567 ;
    wire signal_11568 ;
    wire signal_11569 ;
    wire signal_11570 ;
    wire signal_11571 ;
    wire signal_11572 ;
    wire signal_11573 ;
    wire signal_11574 ;
    wire signal_11575 ;
    wire signal_11576 ;
    wire signal_11577 ;
    wire signal_11578 ;
    wire signal_11579 ;
    wire signal_11580 ;
    wire signal_11581 ;
    wire signal_11582 ;
    wire signal_11583 ;
    wire signal_11584 ;
    wire signal_11585 ;
    wire signal_11586 ;
    wire signal_11587 ;
    wire signal_11588 ;
    wire signal_11589 ;
    wire signal_11590 ;
    wire signal_11591 ;
    wire signal_11592 ;
    wire signal_11593 ;
    wire signal_11594 ;
    wire signal_11595 ;
    wire signal_11596 ;
    wire signal_11597 ;
    wire signal_11598 ;
    wire signal_11599 ;
    wire signal_11600 ;
    wire signal_11601 ;
    wire signal_11602 ;
    wire signal_11603 ;
    wire signal_11604 ;
    wire signal_11605 ;
    wire signal_11606 ;
    wire signal_11607 ;
    wire signal_11608 ;
    wire signal_11609 ;
    wire signal_11610 ;
    wire signal_11611 ;
    wire signal_11612 ;
    wire signal_11613 ;
    wire signal_11614 ;
    wire signal_11615 ;
    wire signal_11616 ;
    wire signal_11617 ;
    wire signal_11618 ;
    wire signal_11619 ;
    wire signal_11620 ;
    wire signal_11621 ;
    wire signal_11622 ;
    wire signal_11623 ;
    wire signal_11624 ;
    wire signal_11625 ;
    wire signal_11626 ;
    wire signal_11627 ;
    wire signal_11628 ;
    wire signal_11629 ;
    wire signal_11630 ;
    wire signal_11631 ;
    wire signal_11632 ;
    wire signal_11633 ;
    wire signal_11634 ;
    wire signal_11635 ;
    wire signal_11636 ;
    wire signal_11637 ;
    wire signal_11638 ;
    wire signal_11639 ;
    wire signal_11640 ;
    wire signal_11641 ;
    wire signal_11642 ;
    wire signal_11643 ;
    wire signal_11644 ;
    wire signal_11645 ;
    wire signal_11646 ;
    wire signal_11647 ;
    wire signal_11648 ;
    wire signal_11649 ;
    wire signal_11650 ;
    wire signal_11651 ;
    wire signal_11652 ;
    wire signal_11653 ;
    wire signal_11654 ;
    wire signal_11655 ;
    wire signal_11656 ;
    wire signal_11657 ;
    wire signal_11658 ;
    wire signal_11659 ;
    wire signal_11660 ;
    wire signal_11661 ;
    wire signal_11662 ;
    wire signal_11663 ;
    wire signal_11664 ;
    wire signal_11665 ;
    wire signal_11666 ;
    wire signal_11667 ;
    wire signal_11668 ;
    wire signal_11669 ;
    wire signal_11670 ;
    wire signal_11671 ;
    wire signal_11672 ;
    wire signal_11673 ;
    wire signal_11674 ;
    wire signal_11675 ;
    wire signal_11676 ;
    wire signal_11677 ;
    wire signal_11678 ;
    wire signal_11679 ;
    wire signal_11680 ;
    wire signal_11681 ;
    wire signal_11682 ;
    wire signal_11683 ;
    wire signal_11684 ;
    wire signal_11685 ;
    wire signal_11686 ;
    wire signal_11687 ;
    wire signal_11688 ;
    wire signal_11689 ;
    wire signal_11690 ;
    wire signal_11691 ;
    wire signal_11692 ;
    wire signal_11693 ;
    wire signal_11694 ;
    wire signal_11695 ;
    wire signal_11696 ;
    wire signal_11697 ;
    wire signal_11698 ;
    wire signal_11699 ;
    wire signal_11700 ;
    wire signal_11701 ;
    wire signal_11702 ;
    wire signal_11703 ;
    wire signal_11704 ;
    wire signal_11705 ;
    wire signal_11706 ;
    wire signal_11707 ;
    wire signal_11708 ;
    wire signal_11709 ;
    wire signal_11710 ;
    wire signal_11711 ;
    wire signal_11712 ;
    wire signal_11713 ;
    wire signal_11714 ;
    wire signal_11715 ;
    wire signal_11716 ;
    wire signal_11717 ;
    wire signal_11718 ;
    wire signal_11719 ;
    wire signal_11720 ;
    wire signal_11721 ;
    wire signal_11722 ;
    wire signal_11723 ;
    wire signal_11724 ;
    wire signal_11725 ;
    wire signal_11726 ;
    wire signal_11727 ;
    wire signal_11728 ;
    wire signal_11729 ;
    wire signal_11730 ;
    wire signal_11731 ;
    wire signal_11732 ;
    wire signal_11733 ;
    wire signal_11734 ;
    wire signal_11735 ;
    wire signal_11736 ;
    wire signal_11737 ;
    wire signal_11738 ;
    wire signal_11739 ;
    wire signal_11740 ;
    wire signal_11741 ;
    wire signal_11742 ;
    wire signal_11743 ;
    wire signal_11744 ;
    wire signal_11745 ;
    wire signal_11746 ;
    wire signal_11747 ;
    wire signal_11748 ;
    wire signal_11749 ;
    wire signal_11750 ;
    wire signal_11751 ;
    wire signal_11752 ;
    wire signal_11753 ;
    wire signal_11754 ;
    wire signal_11755 ;
    wire signal_11756 ;
    wire signal_11757 ;
    wire signal_11758 ;
    wire signal_11759 ;
    wire signal_11760 ;
    wire signal_11761 ;
    wire signal_11762 ;
    wire signal_11763 ;
    wire signal_11764 ;
    wire signal_11765 ;
    wire signal_11766 ;
    wire signal_11767 ;
    wire signal_11768 ;
    wire signal_11769 ;
    wire signal_11770 ;
    wire signal_11771 ;
    wire signal_11772 ;
    wire signal_11773 ;
    wire signal_11774 ;
    wire signal_11775 ;
    wire signal_11776 ;
    wire signal_11777 ;
    wire signal_11778 ;
    wire signal_11779 ;
    wire signal_11780 ;
    wire signal_11781 ;
    wire signal_11782 ;
    wire signal_11783 ;
    wire signal_11784 ;
    wire signal_11785 ;
    wire signal_11786 ;
    wire signal_11787 ;
    wire signal_11788 ;
    wire signal_11789 ;
    wire signal_11790 ;
    wire signal_11791 ;
    wire signal_11792 ;
    wire signal_11793 ;
    wire signal_11794 ;
    wire signal_11795 ;
    wire signal_11796 ;
    wire signal_11797 ;
    wire signal_11798 ;
    wire signal_11799 ;
    wire signal_11800 ;
    wire signal_11801 ;
    wire signal_11802 ;
    wire signal_11803 ;
    wire signal_11804 ;
    wire signal_11805 ;
    wire signal_11806 ;
    wire signal_11807 ;
    wire signal_11808 ;
    wire signal_11809 ;
    wire signal_11810 ;
    wire signal_11811 ;
    wire signal_11812 ;
    wire signal_11813 ;
    wire signal_11814 ;
    wire signal_11815 ;
    wire signal_11816 ;
    wire signal_11817 ;
    wire signal_11818 ;
    wire signal_11819 ;
    wire signal_11820 ;
    wire signal_11821 ;
    wire signal_11822 ;
    wire signal_11823 ;
    wire signal_11824 ;
    wire signal_11825 ;
    wire signal_11826 ;
    wire signal_11827 ;
    wire signal_11828 ;
    wire signal_11829 ;
    wire signal_11830 ;
    wire signal_11831 ;
    wire signal_11832 ;
    wire signal_11833 ;
    wire signal_11834 ;
    wire signal_11835 ;
    wire signal_11836 ;
    wire signal_11837 ;
    wire signal_11838 ;
    wire signal_11839 ;
    wire signal_11840 ;
    wire signal_11841 ;
    wire signal_11842 ;
    wire signal_11843 ;
    wire signal_11844 ;
    wire signal_11845 ;
    wire signal_11846 ;
    wire signal_11847 ;
    wire signal_11848 ;
    wire signal_11849 ;
    wire signal_11850 ;
    wire signal_11851 ;
    wire signal_11852 ;
    wire signal_11853 ;
    wire signal_11854 ;
    wire signal_11855 ;
    wire signal_11856 ;
    wire signal_11857 ;
    wire signal_11858 ;
    wire signal_11859 ;
    wire signal_11860 ;
    wire signal_11861 ;
    wire signal_11862 ;
    wire signal_11863 ;
    wire signal_11864 ;
    wire signal_11865 ;
    wire signal_11866 ;
    wire signal_11867 ;
    wire signal_11868 ;
    wire signal_11869 ;
    wire signal_11870 ;
    wire signal_11871 ;
    wire signal_11872 ;
    wire signal_11873 ;
    wire signal_11874 ;
    wire signal_11875 ;
    wire signal_11876 ;
    wire signal_11877 ;
    wire signal_11878 ;
    wire signal_11879 ;
    wire signal_11880 ;
    wire signal_11881 ;
    wire signal_11882 ;
    wire signal_11883 ;
    wire signal_11884 ;
    wire signal_11885 ;
    wire signal_11886 ;
    wire signal_11887 ;
    wire signal_11888 ;
    wire signal_11889 ;
    wire signal_11890 ;
    wire signal_11891 ;
    wire signal_11892 ;
    wire signal_11893 ;
    wire signal_11894 ;
    wire signal_11895 ;
    wire signal_11896 ;
    wire signal_11897 ;
    wire signal_11898 ;
    wire signal_11899 ;
    wire signal_11900 ;
    wire signal_11901 ;
    wire signal_11902 ;
    wire signal_11903 ;
    wire signal_11904 ;
    wire signal_11905 ;
    wire signal_11906 ;
    wire signal_11907 ;
    wire signal_11908 ;
    wire signal_11909 ;
    wire signal_11910 ;
    wire signal_11911 ;
    wire signal_11912 ;
    wire signal_11913 ;
    wire signal_11914 ;
    wire signal_11915 ;
    wire signal_11916 ;
    wire signal_11917 ;
    wire signal_11918 ;
    wire signal_11919 ;
    wire signal_11920 ;
    wire signal_11921 ;
    wire signal_11922 ;
    wire signal_11923 ;
    wire signal_11924 ;
    wire signal_11925 ;
    wire signal_11926 ;
    wire signal_11927 ;
    wire signal_11928 ;
    wire signal_11929 ;
    wire signal_11930 ;
    wire signal_11931 ;
    wire signal_11932 ;
    wire signal_11933 ;
    wire signal_11934 ;
    wire signal_11935 ;
    wire signal_11936 ;
    wire signal_11937 ;
    wire signal_11938 ;
    wire signal_11939 ;
    wire signal_11940 ;
    wire signal_11941 ;
    wire signal_11942 ;
    wire signal_11943 ;
    wire signal_11944 ;
    wire signal_11945 ;
    wire signal_11946 ;
    wire signal_11947 ;
    wire signal_11948 ;
    wire signal_11949 ;
    wire signal_11950 ;
    wire signal_11951 ;
    wire signal_11952 ;
    wire signal_11953 ;
    wire signal_11954 ;
    wire signal_11955 ;
    wire signal_11956 ;
    wire signal_11957 ;
    wire signal_11958 ;
    wire signal_11959 ;
    wire signal_11960 ;
    wire signal_11961 ;
    wire signal_11962 ;
    wire signal_11963 ;
    wire signal_11964 ;
    wire signal_11965 ;
    wire signal_11966 ;
    wire signal_11967 ;
    wire signal_11968 ;
    wire signal_11969 ;
    wire signal_11970 ;
    wire signal_11971 ;
    wire signal_11972 ;
    wire signal_11973 ;
    wire signal_11974 ;
    wire signal_11975 ;
    wire signal_11976 ;
    wire signal_11977 ;
    wire signal_11978 ;
    wire signal_11979 ;
    wire signal_11980 ;
    wire signal_11981 ;
    wire signal_11982 ;
    wire signal_11983 ;
    wire signal_11984 ;
    wire signal_11985 ;
    wire signal_11986 ;
    wire signal_11987 ;
    wire signal_11988 ;
    wire signal_11989 ;
    wire signal_11990 ;
    wire signal_11991 ;
    wire signal_11992 ;
    wire signal_11993 ;
    wire signal_11994 ;
    wire signal_11995 ;
    wire signal_11996 ;
    wire signal_11997 ;
    wire signal_11998 ;
    wire signal_11999 ;
    wire signal_12000 ;
    wire signal_12001 ;
    wire signal_12002 ;
    wire signal_12003 ;
    wire signal_12004 ;
    wire signal_12005 ;
    wire signal_12006 ;
    wire signal_12007 ;
    wire signal_12008 ;
    wire signal_12009 ;
    wire signal_12010 ;
    wire signal_12011 ;
    wire signal_12012 ;
    wire signal_12013 ;
    wire signal_12014 ;
    wire signal_12015 ;
    wire signal_12016 ;
    wire signal_12017 ;
    wire signal_12018 ;
    wire signal_12019 ;
    wire signal_12020 ;
    wire signal_12021 ;
    wire signal_12022 ;
    wire signal_12023 ;
    wire signal_12024 ;
    wire signal_12025 ;
    wire signal_12026 ;
    wire signal_12027 ;
    wire signal_12028 ;
    wire signal_12029 ;
    wire signal_12030 ;
    wire signal_12031 ;
    wire signal_12032 ;
    wire signal_12033 ;
    wire signal_12034 ;
    wire signal_12035 ;
    wire signal_12036 ;
    wire signal_12037 ;
    wire signal_12038 ;
    wire signal_12039 ;
    wire signal_12040 ;
    wire signal_12041 ;
    wire signal_12042 ;
    wire signal_12043 ;
    wire signal_12044 ;
    wire signal_12045 ;
    wire signal_12046 ;
    wire signal_12047 ;
    wire signal_12048 ;
    wire signal_12049 ;
    wire signal_12050 ;
    wire signal_12051 ;
    wire signal_12052 ;
    wire signal_12053 ;
    wire signal_12054 ;
    wire signal_12055 ;
    wire signal_12056 ;
    wire signal_12057 ;
    wire signal_12058 ;
    wire signal_12059 ;
    wire signal_12060 ;
    wire signal_12061 ;
    wire signal_12062 ;
    wire signal_12063 ;
    wire signal_12064 ;
    wire signal_12065 ;
    wire signal_12066 ;
    wire signal_12067 ;
    wire signal_12068 ;
    wire signal_12069 ;
    wire signal_12070 ;
    wire signal_12071 ;
    wire signal_12072 ;
    wire signal_12073 ;
    wire signal_12074 ;
    wire signal_12075 ;
    wire signal_12076 ;
    wire signal_12077 ;
    wire signal_12078 ;
    wire signal_12079 ;
    wire signal_12080 ;
    wire signal_12081 ;
    wire signal_12082 ;
    wire signal_12083 ;
    wire signal_12084 ;
    wire signal_12085 ;
    wire signal_12086 ;
    wire signal_12087 ;
    wire signal_12088 ;
    wire signal_12089 ;
    wire signal_12090 ;
    wire signal_12091 ;
    wire signal_12092 ;
    wire signal_12093 ;
    wire signal_12094 ;
    wire signal_12095 ;
    wire signal_12096 ;
    wire signal_12097 ;
    wire signal_12098 ;
    wire signal_12099 ;
    wire signal_12100 ;
    wire signal_12101 ;
    wire signal_12102 ;
    wire signal_12103 ;
    wire signal_12104 ;
    wire signal_12105 ;
    wire signal_12106 ;
    wire signal_12107 ;
    wire signal_12108 ;
    wire signal_12109 ;
    wire signal_12110 ;
    wire signal_12111 ;
    wire signal_12112 ;
    wire signal_12113 ;
    wire signal_12114 ;
    wire signal_12115 ;
    wire signal_12116 ;
    wire signal_12117 ;
    wire signal_12118 ;
    wire signal_12119 ;
    wire signal_12120 ;
    wire signal_12121 ;
    wire signal_12122 ;
    wire signal_12123 ;
    wire signal_12124 ;
    wire signal_12125 ;
    wire signal_12126 ;
    wire signal_12127 ;
    wire signal_12128 ;
    wire signal_12129 ;
    wire signal_12130 ;
    wire signal_12131 ;
    wire signal_12132 ;
    wire signal_12133 ;
    wire signal_12134 ;
    wire signal_12135 ;
    wire signal_12136 ;
    wire signal_12137 ;
    wire signal_12138 ;
    wire signal_12139 ;
    wire signal_12140 ;
    wire signal_12141 ;
    wire signal_12142 ;
    wire signal_12143 ;
    wire signal_12144 ;
    wire signal_12145 ;
    wire signal_12146 ;
    wire signal_12147 ;
    wire signal_12148 ;
    wire signal_12149 ;
    wire signal_12150 ;
    wire signal_12151 ;
    wire signal_12152 ;
    wire signal_12153 ;
    wire signal_12154 ;
    wire signal_12155 ;
    wire signal_12156 ;
    wire signal_12157 ;
    wire signal_12158 ;
    wire signal_12159 ;
    wire signal_12160 ;
    wire signal_12161 ;
    wire signal_12162 ;
    wire signal_12163 ;
    wire signal_12164 ;
    wire signal_12165 ;
    wire signal_12166 ;
    wire signal_12167 ;
    wire signal_12168 ;
    wire signal_12169 ;
    wire signal_12170 ;
    wire signal_12171 ;
    wire signal_12172 ;
    wire signal_12173 ;
    wire signal_12174 ;
    wire signal_12175 ;
    wire signal_12176 ;
    wire signal_12177 ;
    wire signal_12178 ;
    wire signal_12179 ;
    wire signal_12180 ;
    wire signal_12181 ;
    wire signal_12182 ;
    wire signal_12183 ;
    wire signal_12184 ;
    wire signal_12185 ;
    wire signal_12186 ;
    wire signal_12187 ;
    wire signal_12188 ;
    wire signal_12189 ;
    wire signal_12190 ;
    wire signal_12191 ;
    wire signal_12192 ;
    wire signal_12193 ;
    wire signal_12194 ;
    wire signal_12195 ;
    wire signal_12196 ;
    wire signal_12197 ;
    wire signal_12198 ;
    wire signal_12199 ;
    wire signal_12200 ;
    wire signal_12201 ;
    wire signal_12202 ;
    wire signal_12203 ;
    wire signal_12204 ;
    wire signal_12205 ;
    wire signal_12206 ;
    wire signal_12207 ;
    wire signal_12208 ;
    wire signal_12209 ;
    wire signal_12210 ;
    wire signal_12211 ;
    wire signal_12212 ;
    wire signal_12213 ;
    wire signal_12214 ;
    wire signal_12215 ;
    wire signal_12216 ;
    wire signal_12217 ;
    wire signal_12218 ;
    wire signal_12219 ;
    wire signal_12220 ;
    wire signal_12221 ;
    wire signal_12222 ;
    wire signal_12223 ;
    wire signal_12224 ;
    wire signal_12225 ;
    wire signal_12226 ;
    wire signal_12227 ;
    wire signal_12228 ;
    wire signal_12229 ;
    wire signal_12230 ;
    wire signal_12231 ;
    wire signal_12232 ;
    wire signal_12233 ;
    wire signal_12234 ;
    wire signal_12235 ;
    wire signal_12236 ;
    wire signal_12237 ;
    wire signal_12238 ;
    wire signal_12239 ;
    wire signal_12240 ;
    wire signal_12241 ;
    wire signal_12242 ;
    wire signal_12243 ;
    wire signal_12244 ;
    wire signal_12245 ;
    wire signal_12246 ;
    wire signal_12247 ;
    wire signal_12248 ;
    wire signal_12249 ;
    wire signal_12250 ;
    wire signal_12251 ;
    wire signal_12252 ;
    wire signal_12253 ;
    wire signal_12254 ;
    wire signal_12255 ;
    wire signal_12256 ;
    wire signal_12257 ;
    wire signal_12258 ;
    wire signal_12259 ;
    wire signal_12260 ;
    wire signal_12261 ;
    wire signal_12262 ;
    wire signal_12263 ;
    wire signal_12264 ;
    wire signal_12265 ;
    wire signal_12266 ;
    wire signal_12267 ;
    wire signal_12268 ;
    wire signal_12269 ;
    wire signal_12270 ;
    wire signal_12271 ;
    wire signal_12272 ;
    wire signal_12273 ;
    wire signal_12274 ;
    wire signal_12275 ;
    wire signal_12276 ;
    wire signal_12277 ;
    wire signal_12278 ;
    wire signal_12279 ;
    wire signal_12280 ;
    wire signal_12281 ;
    wire signal_12282 ;
    wire signal_12283 ;
    wire signal_12284 ;
    wire signal_12285 ;
    wire signal_12286 ;
    wire signal_12287 ;
    wire signal_12288 ;
    wire signal_12289 ;
    wire signal_12290 ;
    wire signal_12291 ;
    wire signal_12292 ;
    wire signal_12293 ;
    wire signal_12294 ;
    wire signal_12295 ;
    wire signal_12296 ;
    wire signal_12297 ;
    wire signal_12298 ;
    wire signal_12299 ;
    wire signal_12300 ;
    wire signal_12301 ;
    wire signal_12302 ;
    wire signal_12303 ;
    wire signal_12304 ;
    wire signal_12305 ;
    wire signal_12306 ;
    wire signal_12307 ;
    wire signal_12308 ;
    wire signal_12309 ;
    wire signal_12310 ;
    wire signal_12311 ;
    wire signal_12312 ;
    wire signal_12313 ;
    wire signal_12314 ;
    wire signal_12315 ;
    wire signal_12316 ;
    wire signal_12317 ;
    wire signal_12318 ;
    wire signal_12319 ;
    wire signal_12320 ;
    wire signal_12321 ;
    wire signal_12322 ;
    wire signal_12323 ;
    wire signal_12324 ;
    wire signal_12325 ;
    wire signal_12326 ;
    wire signal_12327 ;
    wire signal_12328 ;
    wire signal_12329 ;
    wire signal_12330 ;
    wire signal_12331 ;
    wire signal_12332 ;
    wire signal_12333 ;
    wire signal_12334 ;
    wire signal_12335 ;
    wire signal_12336 ;
    wire signal_12337 ;
    wire signal_12338 ;
    wire signal_12339 ;
    wire signal_12340 ;
    wire signal_12341 ;
    wire signal_12342 ;
    wire signal_12343 ;
    wire signal_12344 ;
    wire signal_12345 ;
    wire signal_12346 ;
    wire signal_12347 ;
    wire signal_12348 ;
    wire signal_12349 ;
    wire signal_12350 ;
    wire signal_12351 ;
    wire signal_12352 ;
    wire signal_12353 ;
    wire signal_12354 ;
    wire signal_12355 ;
    wire signal_12356 ;
    wire signal_12357 ;
    wire signal_12358 ;
    wire signal_12359 ;
    wire signal_12360 ;
    wire signal_12361 ;
    wire signal_12362 ;
    wire signal_12363 ;
    wire signal_12364 ;
    wire signal_12365 ;
    wire signal_12366 ;
    wire signal_12367 ;
    wire signal_12368 ;
    wire signal_12369 ;
    wire signal_12370 ;
    wire signal_12371 ;
    wire signal_12372 ;
    wire signal_12373 ;
    wire signal_12374 ;
    wire signal_12375 ;
    wire signal_12376 ;
    wire signal_12377 ;
    wire signal_12378 ;
    wire signal_12379 ;
    wire signal_12380 ;
    wire signal_12381 ;
    wire signal_12382 ;
    wire signal_12383 ;
    wire signal_12384 ;
    wire signal_12385 ;
    wire signal_12386 ;
    wire signal_12387 ;
    wire signal_12388 ;
    wire signal_12389 ;
    wire signal_12390 ;
    wire signal_12391 ;
    wire signal_12392 ;
    wire signal_12393 ;
    wire signal_12394 ;
    wire signal_12395 ;
    wire signal_12396 ;
    wire signal_12397 ;
    wire signal_12398 ;
    wire signal_12399 ;
    wire signal_12400 ;
    wire signal_12401 ;
    wire signal_12402 ;
    wire signal_12403 ;
    wire signal_12404 ;
    wire signal_12405 ;
    wire signal_12406 ;
    wire signal_12407 ;
    wire signal_12408 ;
    wire signal_12409 ;
    wire signal_12410 ;
    wire signal_12411 ;
    wire signal_12412 ;
    wire signal_12413 ;
    wire signal_12414 ;
    wire signal_12415 ;
    wire signal_12416 ;
    wire signal_12417 ;
    wire signal_12418 ;
    wire signal_12419 ;
    wire signal_12420 ;
    wire signal_12421 ;
    wire signal_12422 ;
    wire signal_12423 ;
    wire signal_12424 ;
    wire signal_12425 ;
    wire signal_12426 ;
    wire signal_12427 ;
    wire signal_12428 ;
    wire signal_12429 ;
    wire signal_12430 ;
    wire signal_12431 ;
    wire signal_12432 ;
    wire signal_12433 ;
    wire signal_12434 ;
    wire signal_12435 ;
    wire signal_12436 ;
    wire signal_12437 ;
    wire signal_12438 ;
    wire signal_12439 ;
    wire signal_12440 ;
    wire signal_12441 ;
    wire signal_12442 ;
    wire signal_12443 ;
    wire signal_12444 ;
    wire signal_12445 ;
    wire signal_12446 ;
    wire signal_12447 ;
    wire signal_12448 ;
    wire signal_12449 ;
    wire signal_12450 ;
    wire signal_12451 ;
    wire signal_12452 ;
    wire signal_12453 ;
    wire signal_12454 ;
    wire signal_12455 ;
    wire signal_12456 ;
    wire signal_12457 ;
    wire signal_12458 ;
    wire signal_12459 ;
    wire signal_12460 ;
    wire signal_12461 ;
    wire signal_12462 ;
    wire signal_12463 ;
    wire signal_12464 ;
    wire signal_12465 ;
    wire signal_12466 ;
    wire signal_12467 ;
    wire signal_12468 ;
    wire signal_12469 ;
    wire signal_12470 ;
    wire signal_12471 ;
    wire signal_12472 ;
    wire signal_12473 ;
    wire signal_12474 ;
    wire signal_12475 ;
    wire signal_12476 ;
    wire signal_12477 ;
    wire signal_12478 ;
    wire signal_12479 ;
    wire signal_12480 ;
    wire signal_12481 ;
    wire signal_12482 ;
    wire signal_12483 ;
    wire signal_12484 ;
    wire signal_12485 ;
    wire signal_12486 ;
    wire signal_12487 ;
    wire signal_12488 ;
    wire signal_12489 ;
    wire signal_12490 ;
    wire signal_12491 ;
    wire signal_12492 ;
    wire signal_12493 ;
    wire signal_12494 ;
    wire signal_12495 ;
    wire signal_12496 ;
    wire signal_12497 ;
    wire signal_12498 ;
    wire signal_12499 ;
    wire signal_12500 ;
    wire signal_12501 ;
    wire signal_12502 ;
    wire signal_12503 ;
    wire signal_12504 ;
    wire signal_12505 ;
    wire signal_12506 ;
    wire signal_12507 ;
    wire signal_12508 ;
    wire signal_12509 ;
    wire signal_12510 ;
    wire signal_12511 ;
    wire signal_12512 ;
    wire signal_12513 ;
    wire signal_12514 ;
    wire signal_12515 ;
    wire signal_12516 ;
    wire signal_12517 ;
    wire signal_12518 ;
    wire signal_12519 ;
    wire signal_12520 ;
    wire signal_12521 ;
    wire signal_12522 ;
    wire signal_12523 ;
    wire signal_12524 ;
    wire signal_12525 ;
    wire signal_12526 ;
    wire signal_12527 ;
    wire signal_12528 ;
    wire signal_12529 ;
    wire signal_12530 ;
    wire signal_12531 ;
    wire signal_12532 ;
    wire signal_12533 ;
    wire signal_12534 ;
    wire signal_12535 ;
    wire signal_12536 ;
    wire signal_12537 ;
    wire signal_12538 ;
    wire signal_12539 ;
    wire signal_12540 ;
    wire signal_12541 ;
    wire signal_12542 ;
    wire signal_12543 ;
    wire signal_12544 ;
    wire signal_12545 ;
    wire signal_12546 ;
    wire signal_12547 ;
    wire signal_12548 ;
    wire signal_12549 ;
    wire signal_12550 ;
    wire signal_12551 ;
    wire signal_12552 ;
    wire signal_12553 ;
    wire signal_12554 ;
    wire signal_12555 ;
    wire signal_12556 ;
    wire signal_12557 ;
    wire signal_12558 ;
    wire signal_12559 ;
    wire signal_12560 ;
    wire signal_12561 ;
    wire signal_12562 ;
    wire signal_12563 ;
    wire signal_12564 ;
    wire signal_12565 ;
    wire signal_12566 ;
    wire signal_12567 ;
    wire signal_12568 ;
    wire signal_12569 ;
    wire signal_12570 ;
    wire signal_12571 ;
    wire signal_12572 ;
    wire signal_12573 ;
    wire signal_12574 ;
    wire signal_12575 ;
    wire signal_12576 ;
    wire signal_12577 ;
    wire signal_12578 ;
    wire signal_12579 ;
    wire signal_12580 ;
    wire signal_12581 ;
    wire signal_12582 ;
    wire signal_12583 ;
    wire signal_12584 ;
    wire signal_12585 ;
    wire signal_12586 ;
    wire signal_12587 ;
    wire signal_12588 ;
    wire signal_12589 ;
    wire signal_12590 ;
    wire signal_12591 ;
    wire signal_12592 ;
    wire signal_12593 ;
    wire signal_12594 ;
    wire signal_12595 ;
    wire signal_12596 ;
    wire signal_12597 ;
    wire signal_12598 ;
    wire signal_12599 ;
    wire signal_12600 ;
    wire signal_12601 ;
    wire signal_12602 ;
    wire signal_12603 ;
    wire signal_12604 ;
    wire signal_12605 ;
    wire signal_12606 ;
    wire signal_12607 ;
    wire signal_12608 ;
    wire signal_12609 ;
    wire signal_12610 ;
    wire signal_12611 ;
    wire signal_12612 ;
    wire signal_12613 ;
    wire signal_12614 ;
    wire signal_12615 ;
    wire signal_12616 ;
    wire signal_12617 ;
    wire signal_12618 ;
    wire signal_12619 ;
    wire signal_12620 ;
    wire signal_12621 ;
    wire signal_12622 ;
    wire signal_12623 ;
    wire signal_12624 ;
    wire signal_12625 ;
    wire signal_12626 ;
    wire signal_12627 ;
    wire signal_12628 ;
    wire signal_12629 ;
    wire signal_12630 ;
    wire signal_12631 ;
    wire signal_12632 ;
    wire signal_12633 ;
    wire signal_12634 ;
    wire signal_12635 ;
    wire signal_12636 ;
    wire signal_12637 ;
    wire signal_12638 ;
    wire signal_12639 ;
    wire signal_12640 ;
    wire signal_12641 ;
    wire signal_12642 ;
    wire signal_12643 ;
    wire signal_12644 ;
    wire signal_12645 ;
    wire signal_12646 ;
    wire signal_12647 ;
    wire signal_12648 ;
    wire signal_12649 ;
    wire signal_12650 ;
    wire signal_12651 ;
    wire signal_12652 ;
    wire signal_12653 ;
    wire signal_12654 ;
    wire signal_12655 ;
    wire signal_12656 ;
    wire signal_12657 ;
    wire signal_12658 ;
    wire signal_12659 ;
    wire signal_12660 ;
    wire signal_12661 ;
    wire signal_12662 ;
    wire signal_12663 ;
    wire signal_12664 ;
    wire signal_12665 ;
    wire signal_12666 ;
    wire signal_12667 ;
    wire signal_12668 ;
    wire signal_12669 ;
    wire signal_12670 ;
    wire signal_12671 ;
    wire signal_12672 ;
    wire signal_12673 ;
    wire signal_12674 ;
    wire signal_12675 ;
    wire signal_12676 ;
    wire signal_12677 ;
    wire signal_12678 ;
    wire signal_12679 ;
    wire signal_12680 ;
    wire signal_12681 ;
    wire signal_12682 ;
    wire signal_12683 ;
    wire signal_12684 ;
    wire signal_12685 ;
    wire signal_12686 ;
    wire signal_12687 ;
    wire signal_12688 ;
    wire signal_12689 ;
    wire signal_12690 ;
    wire signal_12691 ;
    wire signal_12692 ;
    wire signal_12693 ;
    wire signal_12694 ;
    wire signal_12695 ;
    wire signal_12696 ;
    wire signal_12697 ;
    wire signal_12698 ;
    wire signal_12699 ;
    wire signal_12700 ;
    wire signal_12701 ;
    wire signal_12702 ;
    wire signal_12703 ;
    wire signal_12704 ;
    wire signal_12705 ;
    wire signal_12706 ;
    wire signal_12707 ;
    wire signal_12708 ;
    wire signal_12709 ;
    wire signal_12710 ;
    wire signal_12711 ;
    wire signal_12712 ;
    wire signal_12713 ;
    wire signal_12714 ;
    wire signal_12715 ;
    wire signal_12716 ;
    wire signal_12717 ;
    wire signal_12718 ;
    wire signal_12719 ;
    wire signal_12720 ;
    wire signal_12721 ;
    wire signal_12722 ;
    wire signal_12723 ;
    wire signal_12724 ;
    wire signal_12725 ;
    wire signal_12726 ;
    wire signal_12727 ;
    wire signal_12728 ;
    wire signal_12729 ;
    wire signal_12730 ;
    wire signal_12731 ;
    wire signal_12732 ;
    wire signal_12733 ;
    wire signal_12734 ;
    wire signal_12735 ;
    wire signal_12736 ;
    wire signal_12737 ;
    wire signal_12738 ;
    wire signal_12739 ;
    wire signal_12740 ;
    wire signal_12741 ;
    wire signal_12742 ;
    wire signal_12743 ;
    wire signal_12744 ;
    wire signal_12745 ;
    wire signal_12746 ;
    wire signal_12747 ;
    wire signal_12748 ;
    wire signal_12749 ;
    wire signal_12750 ;
    wire signal_12751 ;
    wire signal_12752 ;
    wire signal_12753 ;
    wire signal_12754 ;
    wire signal_12755 ;
    wire signal_12756 ;
    wire signal_12757 ;
    wire signal_12758 ;
    wire signal_12759 ;
    wire signal_12760 ;
    wire signal_12761 ;
    wire signal_12762 ;
    wire signal_12763 ;
    wire signal_12764 ;
    wire signal_12765 ;
    wire signal_12766 ;
    wire signal_12767 ;
    wire signal_12768 ;
    wire signal_12769 ;
    wire signal_12770 ;
    wire signal_12771 ;
    wire signal_12772 ;
    wire signal_12773 ;
    wire signal_12774 ;
    wire signal_12775 ;
    wire signal_12776 ;
    wire signal_12777 ;
    wire signal_12778 ;
    wire signal_12779 ;
    wire signal_12780 ;
    wire signal_12781 ;
    wire signal_12782 ;
    wire signal_12783 ;
    wire signal_12784 ;
    wire signal_12785 ;
    wire signal_12786 ;
    wire signal_12787 ;
    wire signal_12788 ;
    wire signal_12789 ;
    wire signal_12790 ;
    wire signal_12791 ;
    wire signal_12792 ;
    wire signal_12793 ;
    wire signal_12794 ;
    wire signal_12795 ;
    wire signal_12796 ;
    wire signal_12797 ;
    wire signal_12798 ;
    wire signal_12799 ;
    wire signal_12800 ;
    wire signal_12801 ;
    wire signal_12802 ;
    wire signal_12803 ;
    wire signal_12804 ;
    wire signal_12805 ;
    wire signal_12806 ;
    wire signal_12807 ;
    wire signal_12808 ;
    wire signal_12809 ;
    wire signal_12810 ;
    wire signal_12811 ;
    wire signal_12812 ;
    wire signal_12813 ;
    wire signal_12814 ;
    wire signal_12815 ;
    wire signal_12816 ;
    wire signal_12817 ;
    wire signal_12818 ;
    wire signal_12819 ;
    wire signal_12820 ;
    wire signal_12821 ;
    wire signal_12822 ;
    wire signal_12823 ;
    wire signal_12824 ;
    wire signal_12825 ;
    wire signal_12826 ;
    wire signal_12827 ;
    wire signal_12828 ;
    wire signal_12829 ;
    wire signal_12830 ;
    wire signal_12831 ;
    wire signal_12832 ;
    wire signal_12833 ;
    wire signal_12834 ;
    wire signal_12835 ;
    wire signal_12836 ;
    wire signal_12837 ;
    wire signal_12838 ;
    wire signal_12839 ;
    wire signal_12840 ;
    wire signal_12841 ;
    wire signal_12842 ;
    wire signal_12843 ;
    wire signal_12844 ;
    wire signal_12845 ;
    wire signal_12846 ;
    wire signal_12847 ;
    wire signal_12848 ;
    wire signal_12849 ;
    wire signal_12850 ;
    wire signal_12851 ;
    wire signal_12852 ;
    wire signal_12853 ;
    wire signal_12854 ;
    wire signal_12855 ;
    wire signal_12856 ;
    wire signal_12857 ;
    wire signal_12858 ;
    wire signal_12859 ;
    wire signal_12860 ;
    wire signal_12861 ;
    wire signal_12862 ;
    wire signal_12863 ;
    wire signal_12864 ;
    wire signal_12865 ;
    wire signal_12866 ;
    wire signal_12867 ;
    wire signal_12868 ;
    wire signal_12869 ;
    wire signal_12870 ;
    wire signal_12871 ;
    wire signal_12872 ;
    wire signal_12873 ;
    wire signal_12874 ;
    wire signal_12875 ;
    wire signal_12876 ;
    wire signal_12877 ;
    wire signal_12878 ;
    wire signal_12879 ;
    wire signal_12880 ;
    wire signal_12881 ;
    wire signal_12882 ;
    wire signal_12883 ;
    wire signal_12884 ;
    wire signal_12885 ;
    wire signal_12886 ;
    wire signal_12887 ;
    wire signal_12888 ;
    wire signal_12889 ;
    wire signal_12890 ;
    wire signal_12891 ;
    wire signal_12892 ;
    wire signal_12893 ;
    wire signal_12894 ;
    wire signal_12895 ;
    wire signal_12896 ;
    wire signal_12897 ;
    wire signal_12898 ;
    wire signal_12899 ;
    wire signal_12900 ;
    wire signal_12901 ;
    wire signal_12902 ;
    wire signal_12903 ;
    wire signal_12904 ;
    wire signal_12905 ;
    wire signal_12906 ;
    wire signal_12907 ;
    wire signal_12908 ;
    wire signal_12909 ;
    wire signal_12910 ;
    wire signal_12911 ;
    wire signal_12912 ;
    wire signal_12913 ;
    wire signal_12914 ;
    wire signal_12915 ;
    wire signal_12916 ;
    wire signal_12917 ;
    wire signal_12918 ;
    wire signal_12919 ;
    wire signal_12920 ;
    wire signal_12921 ;
    wire signal_12922 ;
    wire signal_12923 ;
    wire signal_12924 ;
    wire signal_12925 ;
    wire signal_12926 ;
    wire signal_12927 ;
    wire signal_12928 ;
    wire signal_12929 ;
    wire signal_12930 ;
    wire signal_12931 ;
    wire signal_12932 ;
    wire signal_12933 ;
    wire signal_12934 ;
    wire signal_12935 ;
    wire signal_12936 ;
    wire signal_12937 ;
    wire signal_12938 ;
    wire signal_12939 ;
    wire signal_12940 ;
    wire signal_12941 ;
    wire signal_12942 ;
    wire signal_12943 ;
    wire signal_12944 ;
    wire signal_12945 ;
    wire signal_12946 ;
    wire signal_12947 ;
    wire signal_12948 ;
    wire signal_12949 ;
    wire signal_12950 ;
    wire signal_12951 ;
    wire signal_12952 ;
    wire signal_12953 ;
    wire signal_12954 ;
    wire signal_12955 ;
    wire signal_12956 ;
    wire signal_12957 ;
    wire signal_12958 ;
    wire signal_12959 ;
    wire signal_12960 ;
    wire signal_12961 ;
    wire signal_12962 ;
    wire signal_12963 ;
    wire signal_12964 ;
    wire signal_12965 ;
    wire signal_12966 ;
    wire signal_12967 ;
    wire signal_12968 ;
    wire signal_12969 ;
    wire signal_12970 ;
    wire signal_12971 ;
    wire signal_12972 ;
    wire signal_12973 ;
    wire signal_12974 ;
    wire signal_12975 ;
    wire signal_12976 ;
    wire signal_12977 ;
    wire signal_12978 ;
    wire signal_12979 ;
    wire signal_12980 ;
    wire signal_12981 ;
    wire signal_12982 ;
    wire signal_12983 ;
    wire signal_12984 ;
    wire signal_12985 ;
    wire signal_12986 ;
    wire signal_12987 ;
    wire signal_12988 ;
    wire signal_12989 ;
    wire signal_12990 ;
    wire signal_12991 ;
    wire signal_12992 ;
    wire signal_12993 ;
    wire signal_12994 ;
    wire signal_12995 ;
    wire signal_12996 ;
    wire signal_12997 ;
    wire signal_12998 ;
    wire signal_12999 ;
    wire signal_13000 ;
    wire signal_13001 ;
    wire signal_13002 ;
    wire signal_13003 ;
    wire signal_13004 ;
    wire signal_13005 ;
    wire signal_13006 ;
    wire signal_13007 ;
    wire signal_13008 ;
    wire signal_13009 ;
    wire signal_13010 ;
    wire signal_13011 ;
    wire signal_13012 ;
    wire signal_13013 ;
    wire signal_13014 ;
    wire signal_13015 ;
    wire signal_13016 ;
    wire signal_13017 ;
    wire signal_13018 ;
    wire signal_13019 ;
    wire signal_13020 ;
    wire signal_13021 ;
    wire signal_13022 ;
    wire signal_13023 ;
    wire signal_13024 ;
    wire signal_13025 ;
    wire signal_13026 ;
    wire signal_13027 ;
    wire signal_13028 ;
    wire signal_13029 ;
    wire signal_13030 ;
    wire signal_13031 ;
    wire signal_13032 ;
    wire signal_13033 ;
    wire signal_13034 ;
    wire signal_13035 ;
    wire signal_13036 ;
    wire signal_13037 ;
    wire signal_13038 ;
    wire signal_13039 ;
    wire signal_13040 ;
    wire signal_13041 ;
    wire signal_13042 ;
    wire signal_13043 ;
    wire signal_13044 ;
    wire signal_13045 ;
    wire signal_13046 ;
    wire signal_13047 ;
    wire signal_13048 ;
    wire signal_13049 ;
    wire signal_13050 ;
    wire signal_13051 ;
    wire signal_13052 ;
    wire signal_13053 ;
    wire signal_13054 ;
    wire signal_13055 ;
    wire signal_13056 ;
    wire signal_13057 ;
    wire signal_13058 ;
    wire signal_13059 ;
    wire signal_13060 ;
    wire signal_13061 ;
    wire signal_13062 ;
    wire signal_13063 ;
    wire signal_13064 ;
    wire signal_13065 ;
    wire signal_13066 ;
    wire signal_13067 ;
    wire signal_13068 ;
    wire signal_13069 ;
    wire signal_13070 ;
    wire signal_13071 ;
    wire signal_13072 ;
    wire signal_13073 ;
    wire signal_13074 ;
    wire signal_13075 ;
    wire signal_13076 ;
    wire signal_13077 ;
    wire signal_13078 ;
    wire signal_13079 ;
    wire signal_13080 ;
    wire signal_13081 ;
    wire signal_13082 ;
    wire signal_13083 ;
    wire signal_13084 ;
    wire signal_13085 ;
    wire signal_13086 ;
    wire signal_13087 ;
    wire signal_13088 ;
    wire signal_13089 ;
    wire signal_13090 ;
    wire signal_13091 ;
    wire signal_13092 ;
    wire signal_13093 ;
    wire signal_13094 ;
    wire signal_13095 ;
    wire signal_13096 ;
    wire signal_13097 ;
    wire signal_13098 ;
    wire signal_13099 ;
    wire signal_13100 ;
    wire signal_13101 ;
    wire signal_13102 ;
    wire signal_13103 ;
    wire signal_13104 ;
    wire signal_13105 ;
    wire signal_13106 ;
    wire signal_13107 ;
    wire signal_13108 ;
    wire signal_13109 ;
    wire signal_13110 ;
    wire signal_13111 ;
    wire signal_13112 ;
    wire signal_13113 ;
    wire signal_13114 ;
    wire signal_13115 ;
    wire signal_13116 ;
    wire signal_13117 ;
    wire signal_13118 ;
    wire signal_13119 ;
    wire signal_13120 ;
    wire signal_13121 ;
    wire signal_13122 ;
    wire signal_13123 ;
    wire signal_13124 ;
    wire signal_13125 ;
    wire signal_13126 ;
    wire signal_13127 ;
    wire signal_13128 ;
    wire signal_13129 ;
    wire signal_13130 ;
    wire signal_13131 ;
    wire signal_13132 ;
    wire signal_13133 ;
    wire signal_13134 ;
    wire signal_13135 ;
    wire signal_13136 ;
    wire signal_13137 ;
    wire signal_13138 ;
    wire signal_13139 ;
    wire signal_13140 ;
    wire signal_13141 ;
    wire signal_13142 ;
    wire signal_13143 ;
    wire signal_13144 ;
    wire signal_13145 ;
    wire signal_13146 ;
    wire signal_13147 ;
    wire signal_13148 ;
    wire signal_13149 ;
    wire signal_13150 ;
    wire signal_13151 ;
    wire signal_13152 ;
    wire signal_13153 ;
    wire signal_13154 ;
    wire signal_13155 ;
    wire signal_13156 ;
    wire signal_13157 ;
    wire signal_13158 ;
    wire signal_13159 ;
    wire signal_13160 ;
    wire signal_13161 ;
    wire signal_13162 ;
    wire signal_13163 ;
    wire signal_13164 ;
    wire signal_13165 ;
    wire signal_13166 ;
    wire signal_13167 ;
    wire signal_13168 ;
    wire signal_13169 ;
    wire signal_13170 ;
    wire signal_13171 ;
    wire signal_13172 ;
    wire signal_13173 ;
    wire signal_13174 ;
    wire signal_13175 ;
    wire signal_13176 ;
    wire signal_13177 ;
    wire signal_13178 ;
    wire signal_13179 ;
    wire signal_13180 ;
    wire signal_13181 ;
    wire signal_13182 ;
    wire signal_13183 ;
    wire signal_13184 ;
    wire signal_13185 ;
    wire signal_13186 ;
    wire signal_13187 ;
    wire signal_13188 ;
    wire signal_13189 ;
    wire signal_13190 ;
    wire signal_13191 ;
    wire signal_13192 ;
    wire signal_13193 ;
    wire signal_13194 ;
    wire signal_13195 ;
    wire signal_13196 ;
    wire signal_13197 ;
    wire signal_13198 ;
    wire signal_13199 ;
    wire signal_13200 ;
    wire signal_13201 ;
    wire signal_13202 ;
    wire signal_13203 ;
    wire signal_13204 ;
    wire signal_13205 ;
    wire signal_13206 ;
    wire signal_13207 ;
    wire signal_13208 ;
    wire signal_13209 ;
    wire signal_13210 ;
    wire signal_13211 ;
    wire signal_13212 ;
    wire signal_13213 ;
    wire signal_13214 ;
    wire signal_13215 ;
    wire signal_13216 ;
    wire signal_13217 ;
    wire signal_13218 ;
    wire signal_13219 ;
    wire signal_13220 ;
    wire signal_13221 ;
    wire signal_13222 ;
    wire signal_13223 ;
    wire signal_13224 ;
    wire signal_13225 ;
    wire signal_13226 ;
    wire signal_13227 ;
    wire signal_13228 ;
    wire signal_13229 ;
    wire signal_13230 ;
    wire signal_13231 ;
    wire signal_13232 ;
    wire signal_13233 ;
    wire signal_13234 ;
    wire signal_13235 ;
    wire signal_13236 ;
    wire signal_13237 ;
    wire signal_13238 ;
    wire signal_13239 ;
    wire signal_13240 ;
    wire signal_13241 ;
    wire signal_13242 ;
    wire signal_13243 ;
    wire signal_13244 ;
    wire signal_13245 ;
    wire signal_13246 ;
    wire signal_13247 ;
    wire signal_13248 ;
    wire signal_13249 ;
    wire signal_13250 ;
    wire signal_13251 ;
    wire signal_13252 ;
    wire signal_13253 ;
    wire signal_13254 ;
    wire signal_13255 ;
    wire signal_13256 ;
    wire signal_13257 ;
    wire signal_13258 ;
    wire signal_13259 ;
    wire signal_13260 ;
    wire signal_13261 ;
    wire signal_13262 ;
    wire signal_13263 ;
    wire signal_13264 ;
    wire signal_13265 ;
    wire signal_13266 ;
    wire signal_13267 ;
    wire signal_13268 ;
    wire signal_13269 ;
    wire signal_13270 ;
    wire signal_13271 ;
    wire signal_13272 ;
    wire signal_13273 ;
    wire signal_13274 ;
    wire signal_13275 ;
    wire signal_13276 ;
    wire signal_13277 ;
    wire signal_13278 ;
    wire signal_13279 ;
    wire signal_13280 ;
    wire signal_13281 ;
    wire signal_13282 ;
    wire signal_13283 ;
    wire signal_13284 ;
    wire signal_13285 ;
    wire signal_13286 ;
    wire signal_13287 ;
    wire signal_13288 ;
    wire signal_13289 ;
    wire signal_13290 ;
    wire signal_13291 ;
    wire signal_13292 ;
    wire signal_13293 ;
    wire signal_13294 ;
    wire signal_13295 ;
    wire signal_13296 ;
    wire signal_13297 ;
    wire signal_13298 ;
    wire signal_13299 ;
    wire signal_13300 ;
    wire signal_13301 ;
    wire signal_13302 ;
    wire signal_13303 ;
    wire signal_13304 ;
    wire signal_13305 ;
    wire signal_13306 ;
    wire signal_13307 ;
    wire signal_13308 ;
    wire signal_13309 ;
    wire signal_13310 ;
    wire signal_13311 ;
    wire signal_13312 ;
    wire signal_13313 ;
    wire signal_13314 ;
    wire signal_13315 ;
    wire signal_13316 ;
    wire signal_13317 ;
    wire signal_13318 ;
    wire signal_13319 ;
    wire signal_13320 ;
    wire signal_13321 ;
    wire signal_13322 ;
    wire signal_13323 ;
    wire signal_13324 ;
    wire signal_13325 ;
    wire signal_13326 ;
    wire signal_13327 ;
    wire signal_13328 ;
    wire signal_13329 ;
    wire signal_13330 ;
    wire signal_13331 ;
    wire signal_13332 ;
    wire signal_13333 ;
    wire signal_13334 ;
    wire signal_13335 ;
    wire signal_13336 ;
    wire signal_13337 ;
    wire signal_13338 ;
    wire signal_13339 ;
    wire signal_13340 ;
    wire signal_13341 ;
    wire signal_13342 ;
    wire signal_13343 ;
    wire signal_13344 ;
    wire signal_13345 ;
    wire signal_13346 ;
    wire signal_13347 ;
    wire signal_13348 ;
    wire signal_13349 ;
    wire signal_13350 ;
    wire signal_13351 ;
    wire signal_13352 ;
    wire signal_13353 ;
    wire signal_13354 ;
    wire signal_13355 ;
    wire signal_13356 ;
    wire signal_13357 ;
    wire signal_13358 ;
    wire signal_13359 ;
    wire signal_13360 ;
    wire signal_13361 ;
    wire signal_13362 ;
    wire signal_13363 ;
    wire signal_13364 ;
    wire signal_13365 ;
    wire signal_13366 ;
    wire signal_13367 ;
    wire signal_13368 ;
    wire signal_13369 ;
    wire signal_13370 ;
    wire signal_13371 ;
    wire signal_13372 ;
    wire signal_13373 ;
    wire signal_13374 ;
    wire signal_13375 ;
    wire signal_13376 ;
    wire signal_13377 ;
    wire signal_13378 ;
    wire signal_13379 ;
    wire signal_13380 ;
    wire signal_13381 ;
    wire signal_13382 ;
    wire signal_13383 ;
    wire signal_13384 ;
    wire signal_13385 ;
    wire signal_13386 ;
    wire signal_13387 ;
    wire signal_13388 ;
    wire signal_13389 ;
    wire signal_13390 ;
    wire signal_13391 ;
    wire signal_13392 ;
    wire signal_13393 ;
    wire signal_13394 ;
    wire signal_13395 ;
    wire signal_13396 ;
    wire signal_13397 ;
    wire signal_13398 ;
    wire signal_13399 ;
    wire signal_13400 ;
    wire signal_13401 ;
    wire signal_13402 ;
    wire signal_13403 ;
    wire signal_13404 ;
    wire signal_13405 ;
    wire signal_13406 ;
    wire signal_13407 ;
    wire signal_13408 ;
    wire signal_13409 ;
    wire signal_13410 ;
    wire signal_13411 ;
    wire signal_13412 ;
    wire signal_13413 ;
    wire signal_13414 ;
    wire signal_13415 ;
    wire signal_13416 ;
    wire signal_13417 ;
    wire signal_13418 ;
    wire signal_13419 ;
    wire signal_13420 ;
    wire signal_13421 ;
    wire signal_13422 ;
    wire signal_13423 ;
    wire signal_13424 ;
    wire signal_13425 ;
    wire signal_13426 ;
    wire signal_13427 ;
    wire signal_13428 ;
    wire signal_13429 ;
    wire signal_13430 ;
    wire signal_13431 ;
    wire signal_13432 ;
    wire signal_13433 ;
    wire signal_13434 ;
    wire signal_13435 ;
    wire signal_13436 ;
    wire signal_13437 ;
    wire signal_13438 ;
    wire signal_13439 ;
    wire signal_13440 ;
    wire signal_13441 ;
    wire signal_13442 ;
    wire signal_13443 ;
    wire signal_13444 ;
    wire signal_13445 ;
    wire signal_13446 ;
    wire signal_13447 ;
    wire signal_13448 ;
    wire signal_13449 ;
    wire signal_13450 ;
    wire signal_13451 ;
    wire signal_13452 ;
    wire signal_13453 ;
    wire signal_13454 ;
    wire signal_13455 ;
    wire signal_13456 ;
    wire signal_13457 ;
    wire signal_13458 ;
    wire signal_13459 ;
    wire signal_13460 ;
    wire signal_13461 ;
    wire signal_13462 ;
    wire signal_13463 ;
    wire signal_13464 ;
    wire signal_13465 ;
    wire signal_13466 ;
    wire signal_13467 ;
    wire signal_13468 ;
    wire signal_13469 ;
    wire signal_13470 ;
    wire signal_13471 ;
    wire signal_13472 ;
    wire signal_13473 ;
    wire signal_13474 ;
    wire signal_13475 ;
    wire signal_13476 ;
    wire signal_13477 ;
    wire signal_13478 ;
    wire signal_13479 ;
    wire signal_13480 ;
    wire signal_13481 ;
    wire signal_13482 ;
    wire signal_13483 ;
    wire signal_13484 ;
    wire signal_13485 ;
    wire signal_13486 ;
    wire signal_13487 ;
    wire signal_13488 ;
    wire signal_13489 ;
    wire signal_13490 ;
    wire signal_13491 ;
    wire signal_13492 ;
    wire signal_13493 ;
    wire signal_13494 ;
    wire signal_13495 ;
    wire signal_13496 ;
    wire signal_13497 ;
    wire signal_13498 ;
    wire signal_13499 ;
    wire signal_13500 ;
    wire signal_13501 ;
    wire signal_13502 ;
    wire signal_13503 ;
    wire signal_13504 ;
    wire signal_13505 ;
    wire signal_13506 ;
    wire signal_13507 ;
    wire signal_13508 ;
    wire signal_13509 ;
    wire signal_13510 ;
    wire signal_13511 ;
    wire signal_13512 ;
    wire signal_13513 ;
    wire signal_13514 ;
    wire signal_13515 ;
    wire signal_13516 ;
    wire signal_13517 ;
    wire signal_13518 ;
    wire signal_13519 ;
    wire signal_13520 ;
    wire signal_13521 ;
    wire signal_13522 ;
    wire signal_13523 ;
    wire signal_13524 ;
    wire signal_13525 ;
    wire signal_13526 ;
    wire signal_13527 ;
    wire signal_13528 ;
    wire signal_13529 ;
    wire signal_13530 ;
    wire signal_13531 ;
    wire signal_13532 ;
    wire signal_13533 ;
    wire signal_13534 ;
    wire signal_13535 ;
    wire signal_13536 ;
    wire signal_13537 ;
    wire signal_13538 ;
    wire signal_13539 ;
    wire signal_13540 ;
    wire signal_13541 ;
    wire signal_13542 ;
    wire signal_13543 ;
    wire signal_13544 ;
    wire signal_13545 ;
    wire signal_13546 ;
    wire signal_13547 ;
    wire signal_13548 ;
    wire signal_13549 ;
    wire signal_13550 ;
    wire signal_13551 ;
    wire signal_13552 ;
    wire signal_13553 ;
    wire signal_13554 ;
    wire signal_13555 ;
    wire signal_13556 ;
    wire signal_13557 ;
    wire signal_13558 ;
    wire signal_13559 ;
    wire signal_13560 ;
    wire signal_13561 ;
    wire signal_13562 ;
    wire signal_13563 ;
    wire signal_13564 ;
    wire signal_13565 ;
    wire signal_13566 ;
    wire signal_13567 ;
    wire signal_13568 ;
    wire signal_13569 ;
    wire signal_13570 ;
    wire signal_13571 ;
    wire signal_13572 ;
    wire signal_13573 ;
    wire signal_13574 ;
    wire signal_13575 ;
    wire signal_13576 ;
    wire signal_13577 ;
    wire signal_13578 ;
    wire signal_13579 ;
    wire signal_13580 ;
    wire signal_13581 ;
    wire signal_13582 ;
    wire signal_13583 ;
    wire signal_13584 ;
    wire signal_13585 ;
    wire signal_13586 ;
    wire signal_13587 ;
    wire signal_13588 ;
    wire signal_13589 ;
    wire signal_13590 ;
    wire signal_13591 ;
    wire signal_13592 ;
    wire signal_13593 ;
    wire signal_13594 ;
    wire signal_13595 ;
    wire signal_13596 ;
    wire signal_13597 ;
    wire signal_13598 ;
    wire signal_13599 ;
    wire signal_13600 ;
    wire signal_13601 ;
    wire signal_13602 ;
    wire signal_13603 ;
    wire signal_13604 ;
    wire signal_13605 ;
    wire signal_13606 ;
    wire signal_13607 ;
    wire signal_13608 ;
    wire signal_13609 ;
    wire signal_13610 ;
    wire signal_13611 ;
    wire signal_13612 ;
    wire signal_13613 ;
    wire signal_13614 ;
    wire signal_13615 ;
    wire signal_13616 ;
    wire signal_13617 ;
    wire signal_13618 ;
    wire signal_13619 ;
    wire signal_13620 ;
    wire signal_13621 ;
    wire signal_13622 ;
    wire signal_13623 ;
    wire signal_13624 ;
    wire signal_13625 ;
    wire signal_13626 ;
    wire signal_13627 ;
    wire signal_13628 ;
    wire signal_13629 ;
    wire signal_13630 ;
    wire signal_13631 ;
    wire signal_13632 ;
    wire signal_13633 ;
    wire signal_13634 ;
    wire signal_13635 ;
    wire signal_13636 ;
    wire signal_13637 ;
    wire signal_13638 ;
    wire signal_13639 ;
    wire signal_13640 ;
    wire signal_13641 ;
    wire signal_13642 ;
    wire signal_13643 ;
    wire signal_13644 ;
    wire signal_13645 ;
    wire signal_13646 ;
    wire signal_13647 ;
    wire signal_13648 ;
    wire signal_13649 ;
    wire signal_13650 ;
    wire signal_13651 ;
    wire signal_13652 ;
    wire signal_13653 ;
    wire signal_13654 ;
    wire signal_13655 ;
    wire signal_13656 ;
    wire signal_13657 ;
    wire signal_13658 ;
    wire signal_13659 ;
    wire signal_13660 ;
    wire signal_13661 ;
    wire signal_13662 ;
    wire signal_13663 ;
    wire signal_13664 ;
    wire signal_13665 ;
    wire signal_13666 ;
    wire signal_13667 ;
    wire signal_13668 ;
    wire signal_13669 ;
    wire signal_13670 ;
    wire signal_13671 ;
    wire signal_13672 ;
    wire signal_13673 ;
    wire signal_13674 ;
    wire signal_13675 ;
    wire signal_13676 ;
    wire signal_13677 ;
    wire signal_13678 ;
    wire signal_13679 ;
    wire signal_13680 ;
    wire signal_13681 ;
    wire signal_13682 ;
    wire signal_13683 ;
    wire signal_13684 ;
    wire signal_13685 ;
    wire signal_13686 ;
    wire signal_13687 ;
    wire signal_13688 ;
    wire signal_13689 ;
    wire signal_13690 ;
    wire signal_13691 ;
    wire signal_13692 ;
    wire signal_13693 ;
    wire signal_13694 ;
    wire signal_13695 ;
    wire signal_13696 ;
    wire signal_13697 ;
    wire signal_13698 ;
    wire signal_13699 ;
    wire signal_13700 ;
    wire signal_13701 ;
    wire signal_13702 ;
    wire signal_13703 ;
    wire signal_13704 ;
    wire signal_13705 ;
    wire signal_13706 ;
    wire signal_13707 ;
    wire signal_13708 ;
    wire signal_13709 ;
    wire signal_13710 ;
    wire signal_13711 ;
    wire signal_13712 ;
    wire signal_13713 ;
    wire signal_13714 ;
    wire signal_13715 ;
    wire signal_13716 ;
    wire signal_13717 ;
    wire signal_13718 ;
    wire signal_13719 ;
    wire signal_13720 ;
    wire signal_13721 ;
    wire signal_13722 ;
    wire signal_13723 ;
    wire signal_13724 ;
    wire signal_13725 ;
    wire signal_13726 ;
    wire signal_13727 ;
    wire signal_13728 ;
    wire signal_13729 ;
    wire signal_13730 ;
    wire signal_13731 ;
    wire signal_13732 ;
    wire signal_13733 ;
    wire signal_13734 ;
    wire signal_13735 ;
    wire signal_13736 ;
    wire signal_13737 ;
    wire signal_13738 ;
    wire signal_13739 ;
    wire signal_13740 ;
    wire signal_13741 ;
    wire signal_13742 ;
    wire signal_13743 ;
    wire signal_13744 ;
    wire signal_13745 ;
    wire signal_13746 ;
    wire signal_13747 ;
    wire signal_13748 ;
    wire signal_13749 ;
    wire signal_13750 ;
    wire signal_13751 ;
    wire signal_13752 ;
    wire signal_13753 ;
    wire signal_13754 ;
    wire signal_13755 ;
    wire signal_13756 ;
    wire signal_13757 ;
    wire signal_13758 ;
    wire signal_13759 ;
    wire signal_13760 ;
    wire signal_13761 ;
    wire signal_13762 ;
    wire signal_13763 ;
    wire signal_13764 ;
    wire signal_13765 ;
    wire signal_13766 ;
    wire signal_13767 ;
    wire signal_13768 ;
    wire signal_13769 ;
    wire signal_13770 ;
    wire signal_13771 ;
    wire signal_13772 ;
    wire signal_13773 ;
    wire signal_13774 ;
    wire signal_13775 ;
    wire signal_13776 ;
    wire signal_13777 ;
    wire signal_13778 ;
    wire signal_13779 ;
    wire signal_13780 ;
    wire signal_13781 ;
    wire signal_13782 ;
    wire signal_13783 ;
    wire signal_13784 ;
    wire signal_13785 ;
    wire signal_13786 ;
    wire signal_13787 ;
    wire signal_13788 ;
    wire signal_13789 ;
    wire signal_13790 ;
    wire signal_13791 ;
    wire signal_13792 ;
    wire signal_13793 ;
    wire signal_13794 ;
    wire signal_13795 ;
    wire signal_13796 ;
    wire signal_13797 ;
    wire signal_13798 ;
    wire signal_13799 ;
    wire signal_13800 ;
    wire signal_13801 ;
    wire signal_13802 ;
    wire signal_13803 ;
    wire signal_13804 ;
    wire signal_13805 ;
    wire signal_13806 ;
    wire signal_13807 ;
    wire signal_13808 ;
    wire signal_13809 ;
    wire signal_13810 ;
    wire signal_13811 ;
    wire signal_13812 ;
    wire signal_13813 ;
    wire signal_13814 ;
    wire signal_13815 ;
    wire signal_13816 ;
    wire signal_13817 ;
    wire signal_13818 ;
    wire signal_13819 ;
    wire signal_13820 ;
    wire signal_13821 ;
    wire signal_13822 ;
    wire signal_13823 ;
    wire signal_13824 ;
    wire signal_13825 ;
    wire signal_13826 ;
    wire signal_13827 ;
    wire signal_13828 ;
    wire signal_13829 ;
    wire signal_13830 ;
    wire signal_13831 ;
    wire signal_13832 ;
    wire signal_13833 ;
    wire signal_13834 ;
    wire signal_13835 ;
    wire signal_13836 ;
    wire signal_13837 ;
    wire signal_13838 ;
    wire signal_13839 ;
    wire signal_13840 ;
    wire signal_13841 ;
    wire signal_13842 ;
    wire signal_13843 ;
    wire signal_13844 ;
    wire signal_13845 ;
    wire signal_13846 ;
    wire signal_13847 ;
    wire signal_13848 ;
    wire signal_13849 ;
    wire signal_13850 ;
    wire signal_13851 ;
    wire signal_13852 ;
    wire signal_13853 ;
    wire signal_13854 ;
    wire signal_13855 ;
    wire signal_13856 ;
    wire signal_13857 ;
    wire signal_13858 ;
    wire signal_13859 ;
    wire signal_13860 ;
    wire signal_13861 ;
    wire signal_13862 ;
    wire signal_13863 ;
    wire signal_13864 ;
    wire signal_13865 ;
    wire signal_13866 ;
    wire signal_13867 ;
    wire signal_13868 ;
    wire signal_13869 ;
    wire signal_13870 ;
    wire signal_13871 ;
    wire signal_13872 ;
    wire signal_13873 ;
    wire signal_13874 ;
    wire signal_13875 ;
    wire signal_13876 ;
    wire signal_13877 ;
    wire signal_13878 ;
    wire signal_13879 ;
    wire signal_13880 ;
    wire signal_13881 ;
    wire signal_13882 ;
    wire signal_13883 ;
    wire signal_13884 ;
    wire signal_13885 ;
    wire signal_13886 ;
    wire signal_13887 ;
    wire signal_13888 ;
    wire signal_13889 ;
    wire signal_13890 ;
    wire signal_13891 ;
    wire signal_13892 ;
    wire signal_13893 ;
    wire signal_13894 ;
    wire signal_13895 ;
    wire signal_13896 ;
    wire signal_13897 ;
    wire signal_13898 ;
    wire signal_13899 ;
    wire signal_13900 ;
    wire signal_13901 ;
    wire signal_13902 ;
    wire signal_13903 ;
    wire signal_13904 ;
    wire signal_13905 ;
    wire signal_13906 ;
    wire signal_13907 ;
    wire signal_13908 ;
    wire signal_13909 ;
    wire signal_13910 ;
    wire signal_13911 ;
    wire signal_13912 ;
    wire signal_13913 ;
    wire signal_13914 ;
    wire signal_13915 ;
    wire signal_13916 ;
    wire signal_13917 ;
    wire signal_13918 ;
    wire signal_13919 ;
    wire signal_13920 ;
    wire signal_13921 ;
    wire signal_13922 ;
    wire signal_13923 ;
    wire signal_13924 ;
    wire signal_13925 ;
    wire signal_13926 ;
    wire signal_13927 ;
    wire signal_13928 ;
    wire signal_13929 ;
    wire signal_13930 ;
    wire signal_13931 ;
    wire signal_13932 ;
    wire signal_13933 ;
    wire signal_13934 ;
    wire signal_13935 ;
    wire signal_13936 ;
    wire signal_13937 ;
    wire signal_13938 ;
    wire signal_13939 ;
    wire signal_13940 ;
    wire signal_13941 ;
    wire signal_13942 ;
    wire signal_13943 ;
    wire signal_13944 ;
    wire signal_13945 ;
    wire signal_13946 ;
    wire signal_13947 ;
    wire signal_13948 ;
    wire signal_13949 ;
    wire signal_13950 ;
    wire signal_13951 ;
    wire signal_13952 ;
    wire signal_13953 ;
    wire signal_13954 ;
    wire signal_13955 ;
    wire signal_13956 ;
    wire signal_13957 ;
    wire signal_13958 ;
    wire signal_13959 ;
    wire signal_13960 ;
    wire signal_13961 ;
    wire signal_13962 ;
    wire signal_13963 ;
    wire signal_13964 ;
    wire signal_13965 ;
    wire signal_13966 ;
    wire signal_13967 ;
    wire signal_13968 ;
    wire signal_13969 ;
    wire signal_13970 ;
    wire signal_13971 ;
    wire signal_13972 ;
    wire signal_13973 ;
    wire signal_13974 ;
    wire signal_13975 ;
    wire signal_13976 ;
    wire signal_13977 ;
    wire signal_13978 ;
    wire signal_13979 ;
    wire signal_13980 ;
    wire signal_13981 ;
    wire signal_13982 ;
    wire signal_13983 ;
    wire signal_13984 ;
    wire signal_13985 ;
    wire signal_13986 ;
    wire signal_13987 ;
    wire signal_13988 ;
    wire signal_13989 ;
    wire signal_13990 ;
    wire signal_13991 ;
    wire signal_13992 ;
    wire signal_13993 ;
    wire signal_13994 ;
    wire signal_13995 ;
    wire signal_13996 ;
    wire signal_13997 ;
    wire signal_13998 ;
    wire signal_13999 ;
    wire signal_14000 ;
    wire signal_14001 ;
    wire signal_14002 ;
    wire signal_14003 ;
    wire signal_14004 ;
    wire signal_14005 ;
    wire signal_14006 ;
    wire signal_14007 ;
    wire signal_14008 ;
    wire signal_14009 ;
    wire signal_14010 ;
    wire signal_14011 ;
    wire signal_14012 ;
    wire signal_14013 ;
    wire signal_14014 ;
    wire signal_14015 ;
    wire signal_14016 ;
    wire signal_14017 ;
    wire signal_14018 ;
    wire signal_14019 ;
    wire signal_14020 ;
    wire signal_14021 ;
    wire signal_14022 ;
    wire signal_14023 ;
    wire signal_14024 ;
    wire signal_14025 ;
    wire signal_14026 ;
    wire signal_14027 ;
    wire signal_14028 ;
    wire signal_14029 ;
    wire signal_14030 ;
    wire signal_14031 ;
    wire signal_14032 ;
    wire signal_14033 ;
    wire signal_14034 ;
    wire signal_14035 ;
    wire signal_14036 ;
    wire signal_14037 ;
    wire signal_14038 ;
    wire signal_14039 ;
    wire signal_14040 ;
    wire signal_14041 ;
    wire signal_14042 ;
    wire signal_14043 ;
    wire signal_14044 ;
    wire signal_14045 ;
    wire signal_14046 ;
    wire signal_14047 ;
    wire signal_14048 ;
    wire signal_14049 ;
    wire signal_14050 ;
    wire signal_14051 ;
    wire signal_14052 ;
    wire signal_14053 ;
    wire signal_14054 ;
    wire signal_14055 ;
    wire signal_14056 ;
    wire signal_14057 ;
    wire signal_14058 ;
    wire signal_14059 ;
    wire signal_14060 ;
    wire signal_14061 ;
    wire signal_14062 ;
    wire signal_14063 ;
    wire signal_14064 ;
    wire signal_14065 ;
    wire signal_14066 ;
    wire signal_14067 ;
    wire signal_14068 ;
    wire signal_14069 ;
    wire signal_14070 ;
    wire signal_14071 ;
    wire signal_14072 ;
    wire signal_14073 ;
    wire signal_14074 ;
    wire signal_14075 ;
    wire signal_14076 ;
    wire signal_14077 ;
    wire signal_14078 ;
    wire signal_14079 ;
    wire signal_14080 ;
    wire signal_14081 ;
    wire signal_14082 ;
    wire signal_14083 ;
    wire signal_14084 ;
    wire signal_14085 ;
    wire signal_14086 ;
    wire signal_14087 ;
    wire signal_14088 ;
    wire signal_14089 ;
    wire signal_14090 ;
    wire signal_14091 ;
    wire signal_14092 ;
    wire signal_14093 ;
    wire signal_14094 ;
    wire signal_14095 ;
    wire signal_14096 ;
    wire signal_14097 ;
    wire signal_14098 ;
    wire signal_14099 ;
    wire signal_14100 ;
    wire signal_14101 ;
    wire signal_14102 ;
    wire signal_14103 ;
    wire signal_14104 ;
    wire signal_14105 ;
    wire signal_14106 ;
    wire signal_14107 ;
    wire signal_14108 ;
    wire signal_14109 ;
    wire signal_14110 ;
    wire signal_14111 ;
    wire signal_14112 ;
    wire signal_14113 ;
    wire signal_14114 ;
    wire signal_14115 ;
    wire signal_14116 ;
    wire signal_14117 ;
    wire signal_14118 ;
    wire signal_14119 ;
    wire signal_14120 ;
    wire signal_14121 ;
    wire signal_14122 ;
    wire signal_14123 ;
    wire signal_14124 ;
    wire signal_14125 ;
    wire signal_14126 ;
    wire signal_14127 ;
    wire signal_14128 ;
    wire signal_14129 ;
    wire signal_14130 ;
    wire signal_14131 ;
    wire signal_14132 ;
    wire signal_14133 ;
    wire signal_14134 ;
    wire signal_14135 ;
    wire signal_14136 ;
    wire signal_14137 ;
    wire signal_14138 ;
    wire signal_14139 ;
    wire signal_14140 ;
    wire signal_14141 ;
    wire signal_14142 ;
    wire signal_14143 ;
    wire signal_14144 ;
    wire signal_14145 ;
    wire signal_14146 ;
    wire signal_14147 ;
    wire signal_14148 ;
    wire signal_14149 ;
    wire signal_14150 ;
    wire signal_14151 ;
    wire signal_14152 ;
    wire signal_14153 ;
    wire signal_14154 ;
    wire signal_14155 ;
    wire signal_14156 ;
    wire signal_14157 ;
    wire signal_14158 ;
    wire signal_14159 ;
    wire signal_14160 ;
    wire signal_14161 ;
    wire signal_14162 ;
    wire signal_14163 ;
    wire signal_14164 ;
    wire signal_14165 ;
    wire signal_14166 ;
    wire signal_14167 ;
    wire signal_14168 ;
    wire signal_14169 ;
    wire signal_14170 ;
    wire signal_14171 ;
    wire signal_14172 ;
    wire signal_14173 ;
    wire signal_14174 ;
    wire signal_14175 ;
    wire signal_14176 ;
    wire signal_14177 ;
    wire signal_14178 ;
    wire signal_14179 ;
    wire signal_14180 ;
    wire signal_14181 ;
    wire signal_14182 ;
    wire signal_14183 ;
    wire signal_14184 ;
    wire signal_14185 ;
    wire signal_14186 ;
    wire signal_14187 ;
    wire signal_14188 ;
    wire signal_14189 ;
    wire signal_14190 ;
    wire signal_14191 ;
    wire signal_14192 ;
    wire signal_14193 ;
    wire signal_14194 ;
    wire signal_14195 ;
    wire signal_14196 ;
    wire signal_14197 ;
    wire signal_14198 ;
    wire signal_14199 ;
    wire signal_14200 ;
    wire signal_14201 ;
    wire signal_14202 ;
    wire signal_14203 ;
    wire signal_14204 ;
    wire signal_14205 ;
    wire signal_14206 ;
    wire signal_14207 ;
    wire signal_14208 ;
    wire signal_14209 ;
    wire signal_14210 ;
    wire signal_14211 ;
    wire signal_14212 ;
    wire signal_14213 ;
    wire signal_14214 ;
    wire signal_14215 ;
    wire signal_14216 ;
    wire signal_14217 ;
    wire signal_14218 ;
    wire signal_14219 ;
    wire signal_14220 ;
    wire signal_14221 ;
    wire signal_14222 ;
    wire signal_14223 ;
    wire signal_14224 ;
    wire signal_14225 ;
    wire signal_14226 ;
    wire signal_14227 ;
    wire signal_14228 ;
    wire signal_14229 ;
    wire signal_14230 ;
    wire signal_14231 ;
    wire signal_14232 ;
    wire signal_14233 ;
    wire signal_14234 ;
    wire signal_14235 ;
    wire signal_14236 ;
    wire signal_14237 ;
    wire signal_14238 ;
    wire signal_14239 ;
    wire signal_14240 ;
    wire signal_14241 ;
    wire signal_14242 ;
    wire signal_14243 ;
    wire signal_14244 ;
    wire signal_14245 ;
    wire signal_14246 ;
    wire signal_14247 ;
    wire signal_14248 ;
    wire signal_14249 ;
    wire signal_14250 ;
    wire signal_14251 ;
    wire signal_14252 ;
    wire signal_14253 ;
    wire signal_14254 ;
    wire signal_14255 ;
    wire signal_14256 ;
    wire signal_14257 ;
    wire signal_14258 ;
    wire signal_14259 ;
    wire signal_14260 ;
    wire signal_14261 ;
    wire signal_14262 ;
    wire signal_14263 ;
    wire signal_14264 ;
    wire signal_14265 ;
    wire signal_14266 ;
    wire signal_14267 ;
    wire signal_14268 ;
    wire signal_14269 ;
    wire signal_14270 ;
    wire signal_14271 ;
    wire signal_14272 ;
    wire signal_14273 ;
    wire signal_14274 ;
    wire signal_14275 ;
    wire signal_14276 ;
    wire signal_14277 ;
    wire signal_14278 ;
    wire signal_14279 ;
    wire signal_14280 ;
    wire signal_14281 ;
    wire signal_14282 ;
    wire signal_14283 ;
    wire signal_14284 ;
    wire signal_14285 ;
    wire signal_14286 ;
    wire signal_14287 ;
    wire signal_14288 ;
    wire signal_14289 ;
    wire signal_14290 ;
    wire signal_14291 ;
    wire signal_14292 ;
    wire signal_14293 ;
    wire signal_14294 ;
    wire signal_14295 ;
    wire signal_14296 ;
    wire signal_14297 ;
    wire signal_14298 ;
    wire signal_14299 ;
    wire signal_14300 ;
    wire signal_14301 ;
    wire signal_14302 ;
    wire signal_14303 ;
    wire signal_14304 ;
    wire signal_14305 ;
    wire signal_14306 ;
    wire signal_14307 ;
    wire signal_14308 ;
    wire signal_14309 ;
    wire signal_14310 ;
    wire signal_14311 ;
    wire signal_14312 ;
    wire signal_14313 ;
    wire signal_14314 ;
    wire signal_14315 ;
    wire signal_14316 ;
    wire signal_14317 ;
    wire signal_14318 ;
    wire signal_14319 ;
    wire signal_14320 ;
    wire signal_14321 ;
    wire signal_14322 ;
    wire signal_14323 ;
    wire signal_14324 ;
    wire signal_14325 ;
    wire signal_14326 ;
    wire signal_14327 ;
    wire signal_14328 ;
    wire signal_14329 ;
    wire signal_14330 ;
    wire signal_14331 ;
    wire signal_14332 ;
    wire signal_14333 ;
    wire signal_14334 ;
    wire signal_14335 ;
    wire signal_14336 ;
    wire signal_14337 ;
    wire signal_14338 ;
    wire signal_14339 ;
    wire signal_14340 ;
    wire signal_14341 ;
    wire signal_14342 ;
    wire signal_14343 ;
    wire signal_14344 ;
    wire signal_14345 ;
    wire signal_14346 ;
    wire signal_14347 ;
    wire signal_14348 ;
    wire signal_14349 ;
    wire signal_14350 ;
    wire signal_14351 ;
    wire signal_14352 ;
    wire signal_14353 ;
    wire signal_14354 ;
    wire signal_14355 ;
    wire signal_14356 ;
    wire signal_14357 ;
    wire signal_14358 ;
    wire signal_14359 ;
    wire signal_14360 ;
    wire signal_14361 ;
    wire signal_14362 ;
    wire signal_14363 ;
    wire signal_14364 ;
    wire signal_14365 ;
    wire signal_14366 ;
    wire signal_14367 ;
    wire signal_14368 ;
    wire signal_14369 ;
    wire signal_14370 ;
    wire signal_14371 ;
    wire signal_14372 ;
    wire signal_14373 ;
    wire signal_14374 ;
    wire signal_14375 ;
    wire signal_14376 ;
    wire signal_14377 ;
    wire signal_14378 ;
    wire signal_14379 ;
    wire signal_14380 ;
    wire signal_14381 ;
    wire signal_14382 ;
    wire signal_14383 ;
    wire signal_14384 ;
    wire signal_14385 ;
    wire signal_14386 ;
    wire signal_14387 ;
    wire signal_14388 ;
    wire signal_14389 ;
    wire signal_14390 ;
    wire signal_14391 ;
    wire signal_14392 ;
    wire signal_14393 ;
    wire signal_14394 ;
    wire signal_14395 ;
    wire signal_14396 ;
    wire signal_14397 ;
    wire signal_14398 ;
    wire signal_14399 ;
    wire signal_14400 ;
    wire signal_14401 ;
    wire signal_14402 ;
    wire signal_14403 ;
    wire signal_14404 ;
    wire signal_14405 ;
    wire signal_14406 ;
    wire signal_14407 ;
    wire signal_14408 ;
    wire signal_14409 ;
    wire signal_14410 ;
    wire signal_14411 ;
    wire signal_14412 ;
    wire signal_14413 ;
    wire signal_14414 ;
    wire signal_14415 ;
    wire signal_14416 ;
    wire signal_14417 ;
    wire signal_14418 ;
    wire signal_14419 ;
    wire signal_14420 ;
    wire signal_14421 ;
    wire signal_14422 ;
    wire signal_14423 ;
    wire signal_14424 ;
    wire signal_14425 ;
    wire signal_14426 ;
    wire signal_14427 ;
    wire signal_14428 ;
    wire signal_14429 ;
    wire signal_14430 ;
    wire signal_14431 ;
    wire signal_14432 ;
    wire signal_14433 ;
    wire signal_14434 ;
    wire signal_14435 ;
    wire signal_14436 ;
    wire signal_14437 ;
    wire signal_14438 ;
    wire signal_14439 ;
    wire signal_14440 ;
    wire signal_14441 ;
    wire signal_14442 ;
    wire signal_14443 ;
    wire signal_14444 ;
    wire signal_14445 ;
    wire signal_14446 ;
    wire signal_14447 ;
    wire signal_14448 ;
    wire signal_14449 ;
    wire signal_14450 ;
    wire signal_14451 ;
    wire signal_14452 ;
    wire signal_14453 ;
    wire signal_14454 ;
    wire signal_14455 ;
    wire signal_14456 ;
    wire signal_14457 ;
    wire signal_14458 ;
    wire signal_14459 ;
    wire signal_14460 ;
    wire signal_14461 ;
    wire signal_14462 ;
    wire signal_14463 ;
    wire signal_14464 ;
    wire signal_14465 ;
    wire signal_14466 ;
    wire signal_14467 ;
    wire signal_14468 ;
    wire signal_14469 ;
    wire signal_14470 ;
    wire signal_14471 ;
    wire signal_14472 ;
    wire signal_14473 ;
    wire signal_14474 ;
    wire signal_14475 ;
    wire signal_14476 ;
    wire signal_14477 ;
    wire signal_14478 ;
    wire signal_14479 ;
    wire signal_14480 ;
    wire signal_14481 ;
    wire signal_14482 ;
    wire signal_14483 ;
    wire signal_14484 ;
    wire signal_14485 ;
    wire signal_14486 ;
    wire signal_14487 ;
    wire signal_14488 ;
    wire signal_14489 ;
    wire signal_14490 ;
    wire signal_14491 ;
    wire signal_14492 ;
    wire signal_14493 ;
    wire signal_14494 ;
    wire signal_14495 ;
    wire signal_14496 ;
    wire signal_14497 ;
    wire signal_14498 ;
    wire signal_14499 ;
    wire signal_14500 ;
    wire signal_14501 ;
    wire signal_14502 ;
    wire signal_14503 ;
    wire signal_14504 ;
    wire signal_14505 ;
    wire signal_14506 ;
    wire signal_14507 ;
    wire signal_14508 ;
    wire signal_14509 ;
    wire signal_14510 ;
    wire signal_14511 ;
    wire signal_14512 ;
    wire signal_14513 ;
    wire signal_14514 ;
    wire signal_14515 ;
    wire signal_14516 ;
    wire signal_14517 ;
    wire signal_14518 ;
    wire signal_14519 ;
    wire signal_14520 ;
    wire signal_14521 ;
    wire signal_14522 ;
    wire signal_14523 ;
    wire signal_14524 ;
    wire signal_14525 ;
    wire signal_14526 ;
    wire signal_14527 ;
    wire signal_14528 ;
    wire signal_14529 ;
    wire signal_14530 ;
    wire signal_14531 ;
    wire signal_14532 ;
    wire signal_14533 ;
    wire signal_14534 ;
    wire signal_14535 ;
    wire signal_14536 ;
    wire signal_14537 ;
    wire signal_14538 ;
    wire signal_14539 ;
    wire signal_14540 ;
    wire signal_14541 ;
    wire signal_14542 ;
    wire signal_14543 ;
    wire signal_14544 ;
    wire signal_14545 ;
    wire signal_14546 ;
    wire signal_14547 ;
    wire signal_14548 ;
    wire signal_14549 ;
    wire signal_14550 ;
    wire signal_14551 ;
    wire signal_14552 ;
    wire signal_14553 ;
    wire signal_14554 ;
    wire signal_14555 ;
    wire signal_14556 ;
    wire signal_14557 ;
    wire signal_14558 ;
    wire signal_14559 ;
    wire signal_14560 ;
    wire signal_14561 ;
    wire signal_14562 ;
    wire signal_14563 ;
    wire signal_14564 ;
    wire signal_14565 ;
    wire signal_14566 ;
    wire signal_14567 ;
    wire signal_14568 ;
    wire signal_14569 ;
    wire signal_14570 ;
    wire signal_14571 ;
    wire signal_14572 ;
    wire signal_14573 ;
    wire signal_14574 ;
    wire signal_14575 ;
    wire signal_14576 ;
    wire signal_14577 ;
    wire signal_14578 ;
    wire signal_14579 ;
    wire signal_14580 ;
    wire signal_14581 ;
    wire signal_14582 ;
    wire signal_14583 ;
    wire signal_14584 ;
    wire signal_14585 ;
    wire signal_14586 ;
    wire signal_14587 ;
    wire signal_14588 ;
    wire signal_14589 ;
    wire signal_14590 ;
    wire signal_14591 ;
    wire signal_14592 ;
    wire signal_14593 ;
    wire signal_14594 ;
    wire signal_14595 ;
    wire signal_14596 ;
    wire signal_14597 ;
    wire signal_14598 ;
    wire signal_14599 ;
    wire signal_14600 ;
    wire signal_14601 ;
    wire signal_14602 ;
    wire signal_14603 ;
    wire signal_14604 ;
    wire signal_14605 ;
    wire signal_14606 ;
    wire signal_14607 ;
    wire signal_14608 ;
    wire signal_14609 ;
    wire signal_14610 ;
    wire signal_14611 ;
    wire signal_14612 ;
    wire signal_14613 ;
    wire signal_14614 ;
    wire signal_14615 ;
    wire signal_14616 ;
    wire signal_14617 ;
    wire signal_14618 ;
    wire signal_14619 ;
    wire signal_14620 ;
    wire signal_14621 ;
    wire signal_14622 ;
    wire signal_14623 ;
    wire signal_14624 ;
    wire signal_14625 ;
    wire signal_14626 ;
    wire signal_14627 ;
    wire signal_14628 ;
    wire signal_14629 ;
    wire signal_14630 ;
    wire signal_14631 ;
    wire signal_14632 ;
    wire signal_14633 ;
    wire signal_14634 ;
    wire signal_14635 ;
    wire signal_14636 ;
    wire signal_14637 ;
    wire signal_14638 ;
    wire signal_14639 ;
    wire signal_14640 ;
    wire signal_14641 ;
    wire signal_14642 ;
    wire signal_14643 ;
    wire signal_14644 ;
    wire signal_14645 ;
    wire signal_14646 ;
    wire signal_14647 ;
    wire signal_14648 ;
    wire signal_14649 ;
    wire signal_14650 ;
    wire signal_14651 ;
    wire signal_14652 ;
    wire signal_14653 ;
    wire signal_14654 ;
    wire signal_14655 ;
    wire signal_14656 ;
    wire signal_14657 ;
    wire signal_14658 ;
    wire signal_14659 ;
    wire signal_14660 ;
    wire signal_14661 ;
    wire signal_14662 ;
    wire signal_14663 ;
    wire signal_14664 ;
    wire signal_14665 ;
    wire signal_14666 ;
    wire signal_14667 ;
    wire signal_14668 ;
    wire signal_14669 ;
    wire signal_14670 ;
    wire signal_14671 ;
    wire signal_14672 ;
    wire signal_14673 ;
    wire signal_14674 ;
    wire signal_14675 ;
    wire signal_14676 ;
    wire signal_14677 ;
    wire signal_14678 ;
    wire signal_14679 ;
    wire signal_14680 ;
    wire signal_14681 ;
    wire signal_14682 ;
    wire signal_14683 ;
    wire signal_14684 ;
    wire signal_14685 ;
    wire signal_14686 ;
    wire signal_14687 ;
    wire signal_14688 ;
    wire signal_14689 ;
    wire signal_14690 ;
    wire signal_14691 ;
    wire signal_14692 ;
    wire signal_14693 ;
    wire signal_14694 ;
    wire signal_14695 ;
    wire signal_14696 ;
    wire signal_14697 ;
    wire signal_14698 ;
    wire signal_14699 ;
    wire signal_14700 ;
    wire signal_14701 ;
    wire signal_14702 ;
    wire signal_14703 ;
    wire signal_14704 ;
    wire signal_14705 ;
    wire signal_14706 ;
    wire signal_14707 ;
    wire signal_14708 ;
    wire signal_14709 ;
    wire signal_14710 ;
    wire signal_14711 ;
    wire signal_14712 ;
    wire signal_14713 ;
    wire signal_14714 ;
    wire signal_14715 ;
    wire signal_14716 ;
    wire signal_14717 ;
    wire signal_14718 ;
    wire signal_14719 ;
    wire signal_14720 ;
    wire signal_14721 ;
    wire signal_14722 ;
    wire signal_14723 ;
    wire signal_14724 ;
    wire signal_14725 ;
    wire signal_14726 ;
    wire signal_14727 ;
    wire signal_14728 ;
    wire signal_14729 ;
    wire signal_14730 ;
    wire signal_14731 ;
    wire signal_14732 ;
    wire signal_14733 ;
    wire signal_14734 ;
    wire signal_14735 ;
    wire signal_14736 ;
    wire signal_14737 ;
    wire signal_14738 ;
    wire signal_14739 ;
    wire signal_14740 ;
    wire signal_14741 ;
    wire signal_14742 ;
    wire signal_14743 ;
    wire signal_14744 ;
    wire signal_14745 ;
    wire signal_14746 ;
    wire signal_14747 ;
    wire signal_14748 ;
    wire signal_14749 ;
    wire signal_14750 ;
    wire signal_14751 ;
    wire signal_14752 ;
    wire signal_14753 ;
    wire signal_14754 ;
    wire signal_14755 ;
    wire signal_14756 ;
    wire signal_14757 ;
    wire signal_14758 ;
    wire signal_14759 ;
    wire signal_14760 ;
    wire signal_14761 ;
    wire signal_14762 ;
    wire signal_14763 ;
    wire signal_14764 ;
    wire signal_14765 ;
    wire signal_14766 ;
    wire signal_14767 ;
    wire signal_14768 ;
    wire signal_14769 ;
    wire signal_14770 ;
    wire signal_14771 ;
    wire signal_14772 ;
    wire signal_14773 ;
    wire signal_14774 ;
    wire signal_14775 ;
    wire signal_14776 ;
    wire signal_14777 ;
    wire signal_14778 ;
    wire signal_14779 ;
    wire signal_14780 ;
    wire signal_14781 ;
    wire signal_14782 ;
    wire signal_14783 ;
    wire signal_14784 ;
    wire signal_14785 ;
    wire signal_14786 ;
    wire signal_14787 ;
    wire signal_14788 ;
    wire signal_14789 ;
    wire signal_14790 ;
    wire signal_14791 ;
    wire signal_14792 ;
    wire signal_14793 ;
    wire signal_14794 ;
    wire signal_14795 ;
    wire signal_14796 ;
    wire signal_14797 ;
    wire signal_14798 ;
    wire signal_14799 ;
    wire signal_14800 ;
    wire signal_14801 ;
    wire signal_14802 ;
    wire signal_14803 ;
    wire signal_14804 ;
    wire signal_14805 ;
    wire signal_14806 ;
    wire signal_14807 ;
    wire signal_14808 ;
    wire signal_14809 ;
    wire signal_14810 ;
    wire signal_14811 ;
    wire signal_14812 ;
    wire signal_14813 ;
    wire signal_14814 ;
    wire signal_14815 ;
    wire signal_14816 ;
    wire signal_14817 ;
    wire signal_14818 ;
    wire signal_14819 ;
    wire signal_14820 ;
    wire signal_14821 ;
    wire signal_14822 ;
    wire signal_14823 ;
    wire signal_14824 ;
    wire signal_14825 ;
    wire signal_14826 ;
    wire signal_14827 ;
    wire signal_14828 ;
    wire signal_14829 ;
    wire signal_14830 ;
    wire signal_14831 ;
    wire signal_14832 ;
    wire signal_14833 ;
    wire signal_14834 ;
    wire signal_14835 ;
    wire signal_14836 ;
    wire signal_14837 ;
    wire signal_14838 ;
    wire signal_14839 ;
    wire signal_14840 ;
    wire signal_14841 ;
    wire signal_14842 ;
    wire signal_14843 ;
    wire signal_14844 ;
    wire signal_14845 ;
    wire signal_14846 ;
    wire signal_14847 ;
    wire signal_14848 ;
    wire signal_14849 ;
    wire signal_14850 ;
    wire signal_14851 ;
    wire signal_14852 ;
    wire signal_14853 ;
    wire signal_14854 ;
    wire signal_14855 ;
    wire signal_14856 ;
    wire signal_14857 ;
    wire signal_14858 ;
    wire signal_14859 ;
    wire signal_14860 ;
    wire signal_14861 ;
    wire signal_14862 ;
    wire signal_14863 ;
    wire signal_14864 ;
    wire signal_14865 ;
    wire signal_14866 ;
    wire signal_14867 ;
    wire signal_14868 ;
    wire signal_14869 ;
    wire signal_14870 ;
    wire signal_14871 ;
    wire signal_14872 ;
    wire signal_14873 ;
    wire signal_14874 ;
    wire signal_14875 ;
    wire signal_14876 ;
    wire signal_14877 ;
    wire signal_14878 ;
    wire signal_14879 ;
    wire signal_14880 ;
    wire signal_14881 ;
    wire signal_14882 ;
    wire signal_14883 ;
    wire signal_14884 ;
    wire signal_14885 ;
    wire signal_14886 ;
    wire signal_14887 ;
    wire signal_14888 ;
    wire signal_14889 ;
    wire signal_14890 ;
    wire signal_14891 ;
    wire signal_14892 ;
    wire signal_14893 ;
    wire signal_14894 ;
    wire signal_14895 ;
    wire signal_14896 ;
    wire signal_14897 ;
    wire signal_14898 ;
    wire signal_14899 ;
    wire signal_14900 ;
    wire signal_14901 ;
    wire signal_14902 ;
    wire signal_14903 ;
    wire signal_14904 ;
    wire signal_14905 ;
    wire signal_14906 ;
    wire signal_14907 ;
    wire signal_14908 ;
    wire signal_14909 ;
    wire signal_14910 ;
    wire signal_14911 ;
    wire signal_14912 ;
    wire signal_14913 ;
    wire signal_14914 ;
    wire signal_14915 ;
    wire signal_14916 ;
    wire signal_14917 ;
    wire signal_14918 ;
    wire signal_14919 ;
    wire signal_14920 ;
    wire signal_14921 ;
    wire signal_14922 ;
    wire signal_14923 ;
    wire signal_14924 ;
    wire signal_14925 ;
    wire signal_14926 ;
    wire signal_14927 ;
    wire signal_14928 ;
    wire signal_14929 ;
    wire signal_14930 ;
    wire signal_14931 ;
    wire signal_14932 ;
    wire signal_14933 ;
    wire signal_14934 ;
    wire signal_14935 ;
    wire signal_14936 ;
    wire signal_14937 ;
    wire signal_14938 ;
    wire signal_14939 ;
    wire signal_14940 ;
    wire signal_14941 ;
    wire signal_14942 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_404) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_2406, signal_1493}), .c ({signal_2407, signal_1413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_2 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2409, signal_1492}), .c ({signal_2410, signal_1412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_3 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_2412, signal_1491}), .c ({signal_2413, signal_1411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_4 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2415, signal_1490}), .c ({signal_2416, signal_1410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_5 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2418, signal_1489}), .c ({signal_2419, signal_1409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_6 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2421, signal_1488}), .c ({signal_2422, signal_1408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_7 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2424, signal_1487}), .c ({signal_2425, signal_1407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_8 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2427, signal_1486}), .c ({signal_2428, signal_1406}) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_399), .A2 (signal_398), .ZN (signal_405) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_402), .A2 (signal_405), .ZN (done) ) ;
    AND2_X1 cell_11 ( .A1 (signal_401), .A2 (signal_396), .ZN (signal_400) ) ;
    INV_X1 cell_12 ( .A (start), .ZN (signal_403) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_406), .A2 (signal_415), .ZN (signal_422) ) ;
    XNOR2_X1 cell_14 ( .A (signal_424), .B (signal_425), .ZN (signal_423) ) ;
    NOR2_X1 cell_15 ( .A1 (signal_407), .A2 (signal_408), .ZN (signal_398) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_421), .A2 (signal_416), .ZN (signal_408) ) ;
    INV_X1 cell_17 ( .A (signal_406), .ZN (signal_407) ) ;
    INV_X1 cell_18 ( .A (signal_420), .ZN (signal_416) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_409), .A2 (signal_410), .ZN (signal_419) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_396), .A2 (signal_418), .ZN (signal_409) ) ;
    NOR2_X1 cell_21 ( .A1 (signal_427), .A2 (signal_424), .ZN (signal_413) ) ;
    NOR2_X1 cell_22 ( .A1 (signal_425), .A2 (signal_428), .ZN (signal_412) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_415), .A2 (signal_414), .ZN (signal_396) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_420), .A2 (signal_421), .ZN (signal_414) ) ;
    INV_X1 cell_25 ( .A (signal_393), .ZN (signal_415) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_412), .A2 (signal_413), .ZN (signal_411) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_426), .A2 (signal_411), .ZN (signal_406) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_393), .A2 (signal_406), .ZN (signal_410) ) ;
    INV_X1 cell_29 ( .A (signal_410), .ZN (signal_395) ) ;
    NOR2_X1 cell_30 ( .A1 (signal_417), .A2 (signal_415), .ZN (signal_394) ) ;
    MUX2_X1 cell_31 ( .S (signal_393), .A (1'b1), .B (signal_423), .Z (signal_429) ) ;
    MUX2_X1 cell_34 ( .S (signal_393), .A (1'b0), .B (signal_425), .Z (signal_431) ) ;
    MUX2_X1 cell_37 ( .S (signal_393), .A (1'b1), .B (signal_426), .Z (signal_433) ) ;
    MUX2_X1 cell_40 ( .S (signal_393), .A (1'b0), .B (signal_427), .Z (signal_435) ) ;
    MUX2_X1 cell_43 ( .S (signal_393), .A (1'b1), .B (signal_428), .Z (signal_437) ) ;
    MUX2_X1 cell_46 ( .S (signal_422), .A (1'b1), .B (signal_416), .Z (signal_439) ) ;
    MUX2_X1 cell_49 ( .S (signal_422), .A (1'b0), .B (signal_421), .Z (signal_441) ) ;
    INV_X1 cell_52 ( .A (signal_418), .ZN (signal_417) ) ;
    INV_X1 cell_64 ( .A (signal_394), .ZN (signal_453) ) ;
    INV_X1 cell_65 ( .A (signal_453), .ZN (signal_455) ) ;
    INV_X1 cell_66 ( .A (signal_393), .ZN (signal_444) ) ;
    INV_X1 cell_67 ( .A (signal_444), .ZN (signal_452) ) ;
    INV_X1 cell_68 ( .A (signal_456), .ZN (signal_464) ) ;
    INV_X1 cell_69 ( .A (signal_453), .ZN (signal_454) ) ;
    INV_X1 cell_70 ( .A (signal_444), .ZN (signal_448) ) ;
    INV_X1 cell_71 ( .A (signal_456), .ZN (signal_460) ) ;
    INV_X1 cell_72 ( .A (signal_444), .ZN (signal_446) ) ;
    INV_X1 cell_73 ( .A (signal_456), .ZN (signal_458) ) ;
    INV_X1 cell_74 ( .A (signal_444), .ZN (signal_450) ) ;
    INV_X1 cell_75 ( .A (signal_456), .ZN (signal_462) ) ;
    INV_X1 cell_76 ( .A (signal_444), .ZN (signal_445) ) ;
    INV_X1 cell_77 ( .A (signal_456), .ZN (signal_457) ) ;
    INV_X1 cell_78 ( .A (signal_444), .ZN (signal_447) ) ;
    INV_X1 cell_79 ( .A (signal_456), .ZN (signal_459) ) ;
    INV_X1 cell_80 ( .A (signal_444), .ZN (signal_449) ) ;
    INV_X1 cell_81 ( .A (signal_456), .ZN (signal_461) ) ;
    INV_X1 cell_82 ( .A (signal_444), .ZN (signal_451) ) ;
    INV_X1 cell_83 ( .A (signal_456), .ZN (signal_463) ) ;
    INV_X1 cell_84 ( .A (signal_395), .ZN (signal_456) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_85 ( .s (signal_457), .b ({signal_2579, signal_1677}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_3820, signal_465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_88 ( .s (signal_457), .b ({signal_2582, signal_1676}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_3821, signal_467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_91 ( .s (signal_457), .b ({signal_2585, signal_1675}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_3822, signal_469}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_94 ( .s (signal_457), .b ({signal_2588, signal_1674}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_3823, signal_471}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_97 ( .s (signal_457), .b ({signal_2591, signal_1673}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_3824, signal_473}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_100 ( .s (signal_457), .b ({signal_2594, signal_1672}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_3825, signal_475}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_103 ( .s (signal_457), .b ({signal_2597, signal_1671}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_3826, signal_477}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_106 ( .s (signal_457), .b ({signal_2600, signal_1670}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_3827, signal_479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_109 ( .s (signal_457), .b ({signal_2603, signal_1669}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({signal_3828, signal_481}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_112 ( .s (signal_457), .b ({signal_2606, signal_1668}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_3829, signal_483}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_115 ( .s (signal_457), .b ({signal_2609, signal_1667}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({signal_3830, signal_485}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_118 ( .s (signal_457), .b ({signal_2612, signal_1666}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_3831, signal_487}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_121 ( .s (signal_457), .b ({signal_2615, signal_1665}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_3832, signal_489}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_124 ( .s (signal_457), .b ({signal_2618, signal_1664}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_3833, signal_491}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_127 ( .s (signal_457), .b ({signal_2621, signal_1663}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_3834, signal_493}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_130 ( .s (signal_457), .b ({signal_2624, signal_1662}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_3835, signal_495}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_133 ( .s (signal_458), .b ({signal_2627, signal_1661}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({signal_3836, signal_497}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_136 ( .s (signal_458), .b ({signal_2630, signal_1660}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_3837, signal_499}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_139 ( .s (signal_458), .b ({signal_2633, signal_1659}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({signal_3838, signal_501}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_142 ( .s (signal_458), .b ({signal_2636, signal_1658}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_3839, signal_503}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_145 ( .s (signal_458), .b ({signal_2639, signal_1657}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_3840, signal_505}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_148 ( .s (signal_458), .b ({signal_2642, signal_1656}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_3841, signal_507}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_151 ( .s (signal_458), .b ({signal_2645, signal_1655}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_3842, signal_509}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_154 ( .s (signal_458), .b ({signal_2648, signal_1654}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_3843, signal_511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_157 ( .s (signal_458), .b ({signal_3628, signal_1653}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_3844, signal_513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_160 ( .s (signal_458), .b ({signal_3630, signal_1652}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_3845, signal_515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_163 ( .s (signal_458), .b ({signal_3632, signal_1651}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_3846, signal_517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_166 ( .s (signal_458), .b ({signal_3634, signal_1650}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_3847, signal_519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_169 ( .s (signal_458), .b ({signal_3636, signal_1649}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({signal_3848, signal_521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_172 ( .s (signal_458), .b ({signal_3638, signal_1648}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({signal_3849, signal_523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_175 ( .s (signal_458), .b ({signal_3640, signal_1647}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_3850, signal_525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_178 ( .s (signal_458), .b ({signal_3642, signal_1646}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_3851, signal_527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_181 ( .s (signal_459), .b ({signal_2651, signal_1645}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({signal_3852, signal_529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_184 ( .s (signal_459), .b ({signal_2654, signal_1644}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_3853, signal_531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_187 ( .s (signal_459), .b ({signal_2657, signal_1643}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({signal_3854, signal_533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_190 ( .s (signal_459), .b ({signal_2660, signal_1642}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_3855, signal_535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_193 ( .s (signal_459), .b ({signal_2663, signal_1641}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_3856, signal_537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_196 ( .s (signal_459), .b ({signal_2666, signal_1640}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_3857, signal_539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_199 ( .s (signal_459), .b ({signal_2669, signal_1639}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_3858, signal_541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_202 ( .s (signal_459), .b ({signal_2672, signal_1638}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_3859, signal_543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_205 ( .s (signal_459), .b ({signal_2675, signal_1637}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({signal_3860, signal_545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_208 ( .s (signal_459), .b ({signal_2678, signal_1636}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_3861, signal_547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_211 ( .s (signal_459), .b ({signal_2681, signal_1635}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({signal_3862, signal_549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_214 ( .s (signal_459), .b ({signal_2684, signal_1634}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_3863, signal_551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_217 ( .s (signal_459), .b ({signal_2687, signal_1633}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_3864, signal_553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_220 ( .s (signal_459), .b ({signal_2690, signal_1632}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_3865, signal_555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_223 ( .s (signal_459), .b ({signal_2693, signal_1631}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_3866, signal_557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_226 ( .s (signal_459), .b ({signal_2696, signal_1630}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_3867, signal_559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_229 ( .s (signal_460), .b ({signal_2699, signal_1629}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({signal_3868, signal_561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_232 ( .s (signal_460), .b ({signal_2702, signal_1628}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_3869, signal_563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_235 ( .s (signal_460), .b ({signal_2705, signal_1627}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({signal_3870, signal_565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_238 ( .s (signal_460), .b ({signal_2708, signal_1626}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_3871, signal_567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_241 ( .s (signal_460), .b ({signal_2711, signal_1625}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_3872, signal_569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_244 ( .s (signal_460), .b ({signal_2714, signal_1624}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_3873, signal_571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_247 ( .s (signal_460), .b ({signal_2717, signal_1623}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_3874, signal_573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_250 ( .s (signal_460), .b ({signal_2720, signal_1622}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_3875, signal_575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_253 ( .s (signal_460), .b ({signal_3644, signal_1621}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_3876, signal_577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_256 ( .s (signal_460), .b ({signal_3646, signal_1620}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_3877, signal_579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_259 ( .s (signal_460), .b ({signal_3648, signal_1619}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_3878, signal_581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_262 ( .s (signal_460), .b ({signal_3650, signal_1618}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_3879, signal_583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_265 ( .s (signal_460), .b ({signal_3652, signal_1617}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_3880, signal_585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_268 ( .s (signal_460), .b ({signal_3654, signal_1616}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_3881, signal_587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_271 ( .s (signal_460), .b ({signal_3656, signal_1615}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_3882, signal_589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_274 ( .s (signal_460), .b ({signal_3658, signal_1614}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_3883, signal_591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_277 ( .s (signal_461), .b ({signal_2723, signal_1613}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({signal_3884, signal_593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_280 ( .s (signal_461), .b ({signal_2726, signal_1612}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_3885, signal_595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_283 ( .s (signal_461), .b ({signal_2729, signal_1611}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({signal_3886, signal_597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_286 ( .s (signal_461), .b ({signal_2732, signal_1610}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_3887, signal_599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_289 ( .s (signal_461), .b ({signal_2735, signal_1609}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_3888, signal_601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_292 ( .s (signal_461), .b ({signal_2738, signal_1608}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_3889, signal_603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_295 ( .s (signal_461), .b ({signal_2741, signal_1607}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_3890, signal_605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_298 ( .s (signal_461), .b ({signal_2744, signal_1606}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_3891, signal_607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_301 ( .s (signal_461), .b ({signal_2747, signal_1605}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({signal_3892, signal_609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_304 ( .s (signal_461), .b ({signal_2750, signal_1604}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_3893, signal_611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_307 ( .s (signal_461), .b ({signal_2753, signal_1603}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({signal_3894, signal_613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_310 ( .s (signal_461), .b ({signal_2756, signal_1602}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_3895, signal_615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_313 ( .s (signal_461), .b ({signal_2759, signal_1601}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_3896, signal_617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_316 ( .s (signal_461), .b ({signal_2762, signal_1600}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_3897, signal_619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_319 ( .s (signal_461), .b ({signal_2765, signal_1599}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_3898, signal_621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_322 ( .s (signal_461), .b ({signal_2768, signal_1598}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_3899, signal_623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_325 ( .s (signal_462), .b ({signal_2771, signal_1597}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_3900, signal_625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_328 ( .s (signal_462), .b ({signal_2774, signal_1596}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_3901, signal_627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_331 ( .s (signal_462), .b ({signal_2777, signal_1595}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_3902, signal_629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_334 ( .s (signal_462), .b ({signal_2780, signal_1594}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_3903, signal_631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_337 ( .s (signal_462), .b ({signal_2783, signal_1593}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_3904, signal_633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_340 ( .s (signal_462), .b ({signal_2786, signal_1592}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_3905, signal_635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_343 ( .s (signal_462), .b ({signal_2789, signal_1591}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_3906, signal_637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_346 ( .s (signal_462), .b ({signal_2792, signal_1590}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_3907, signal_639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_349 ( .s (signal_462), .b ({signal_3660, signal_1589}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({signal_3908, signal_641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_352 ( .s (signal_462), .b ({signal_3662, signal_1588}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_3909, signal_643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_355 ( .s (signal_462), .b ({signal_3664, signal_1587}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({signal_3910, signal_645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_358 ( .s (signal_462), .b ({signal_3666, signal_1586}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_3911, signal_647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_361 ( .s (signal_462), .b ({signal_3668, signal_1585}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_3912, signal_649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_364 ( .s (signal_462), .b ({signal_3670, signal_1584}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_3913, signal_651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_367 ( .s (signal_462), .b ({signal_3672, signal_1583}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_3914, signal_653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_370 ( .s (signal_462), .b ({signal_3674, signal_1582}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_3915, signal_655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_373 ( .s (signal_463), .b ({signal_2795, signal_1581}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({signal_3916, signal_657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_376 ( .s (signal_463), .b ({signal_2798, signal_1580}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_3917, signal_659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_379 ( .s (signal_463), .b ({signal_2801, signal_1579}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({signal_3918, signal_661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_382 ( .s (signal_463), .b ({signal_2804, signal_1578}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_3919, signal_663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_385 ( .s (signal_463), .b ({signal_2807, signal_1577}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_3920, signal_665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_388 ( .s (signal_463), .b ({signal_2810, signal_1576}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_3921, signal_667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_391 ( .s (signal_463), .b ({signal_2813, signal_1575}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_3922, signal_669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_394 ( .s (signal_463), .b ({signal_2816, signal_1574}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_3923, signal_671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_397 ( .s (signal_463), .b ({signal_2819, signal_1573}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_3924, signal_673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_400 ( .s (signal_463), .b ({signal_2822, signal_1572}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_3925, signal_675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_403 ( .s (signal_463), .b ({signal_2825, signal_1571}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_3926, signal_677}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_406 ( .s (signal_463), .b ({signal_2828, signal_1570}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_3927, signal_679}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_409 ( .s (signal_463), .b ({signal_2831, signal_1569}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_3928, signal_681}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_412 ( .s (signal_463), .b ({signal_2834, signal_1568}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_3929, signal_683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_415 ( .s (signal_463), .b ({signal_2837, signal_1567}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_3930, signal_685}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_418 ( .s (signal_463), .b ({signal_2840, signal_1566}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_3931, signal_687}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_421 ( .s (signal_464), .b ({signal_2843, signal_1565}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({signal_3932, signal_689}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_424 ( .s (signal_464), .b ({signal_2846, signal_1564}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_3933, signal_691}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_427 ( .s (signal_464), .b ({signal_2849, signal_1563}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({signal_3934, signal_693}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_430 ( .s (signal_464), .b ({signal_2852, signal_1562}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_3935, signal_695}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_433 ( .s (signal_464), .b ({signal_2855, signal_1561}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_3936, signal_697}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_436 ( .s (signal_464), .b ({signal_2858, signal_1560}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_3937, signal_699}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_439 ( .s (signal_464), .b ({signal_2861, signal_1559}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_3938, signal_701}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_442 ( .s (signal_464), .b ({signal_2864, signal_1558}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_3939, signal_703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_469 ( .s (signal_445), .b ({plaintext_s1[120], plaintext_s0[120]}), .a ({ciphertext_s1[112], ciphertext_s0[112]}), .c ({signal_2579, signal_1677}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_470 ( .s (signal_445), .b ({plaintext_s1[121], plaintext_s0[121]}), .a ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_2582, signal_1676}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_471 ( .s (signal_445), .b ({plaintext_s1[122], plaintext_s0[122]}), .a ({ciphertext_s1[114], ciphertext_s0[114]}), .c ({signal_2585, signal_1675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_472 ( .s (signal_445), .b ({plaintext_s1[123], plaintext_s0[123]}), .a ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_2588, signal_1674}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_473 ( .s (signal_445), .b ({plaintext_s1[124], plaintext_s0[124]}), .a ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_2591, signal_1673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_474 ( .s (signal_445), .b ({plaintext_s1[125], plaintext_s0[125]}), .a ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_2594, signal_1672}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_475 ( .s (signal_445), .b ({plaintext_s1[126], plaintext_s0[126]}), .a ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_2597, signal_1671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_476 ( .s (signal_445), .b ({plaintext_s1[127], plaintext_s0[127]}), .a ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_2600, signal_1670}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_477 ( .s (signal_445), .b ({plaintext_s1[112], plaintext_s0[112]}), .a ({ciphertext_s1[104], ciphertext_s0[104]}), .c ({signal_2603, signal_1669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_478 ( .s (signal_445), .b ({plaintext_s1[113], plaintext_s0[113]}), .a ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_2606, signal_1668}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_479 ( .s (signal_445), .b ({plaintext_s1[114], plaintext_s0[114]}), .a ({ciphertext_s1[106], ciphertext_s0[106]}), .c ({signal_2609, signal_1667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_480 ( .s (signal_445), .b ({plaintext_s1[115], plaintext_s0[115]}), .a ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_2612, signal_1666}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_481 ( .s (signal_445), .b ({plaintext_s1[116], plaintext_s0[116]}), .a ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_2615, signal_1665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_482 ( .s (signal_445), .b ({plaintext_s1[117], plaintext_s0[117]}), .a ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_2618, signal_1664}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_483 ( .s (signal_445), .b ({plaintext_s1[118], plaintext_s0[118]}), .a ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_2621, signal_1663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_484 ( .s (signal_445), .b ({plaintext_s1[119], plaintext_s0[119]}), .a ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_2624, signal_1662}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_485 ( .s (signal_446), .b ({plaintext_s1[104], plaintext_s0[104]}), .a ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_2627, signal_1661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_486 ( .s (signal_446), .b ({plaintext_s1[105], plaintext_s0[105]}), .a ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_2630, signal_1660}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_487 ( .s (signal_446), .b ({plaintext_s1[106], plaintext_s0[106]}), .a ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_2633, signal_1659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_488 ( .s (signal_446), .b ({plaintext_s1[107], plaintext_s0[107]}), .a ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_2636, signal_1658}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_489 ( .s (signal_446), .b ({plaintext_s1[108], plaintext_s0[108]}), .a ({ciphertext_s1[100], ciphertext_s0[100]}), .c ({signal_2639, signal_1657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_490 ( .s (signal_446), .b ({plaintext_s1[109], plaintext_s0[109]}), .a ({ciphertext_s1[101], ciphertext_s0[101]}), .c ({signal_2642, signal_1656}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_491 ( .s (signal_446), .b ({plaintext_s1[110], plaintext_s0[110]}), .a ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_2645, signal_1655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_492 ( .s (signal_446), .b ({plaintext_s1[111], plaintext_s0[111]}), .a ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_2648, signal_1654}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_493 ( .s (signal_454), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_3298, signal_1429}), .c ({signal_3452, signal_1549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_494 ( .s (signal_454), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_3299, signal_1428}), .c ({signal_3453, signal_1548}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_495 ( .s (signal_454), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_3300, signal_1427}), .c ({signal_3454, signal_1547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_496 ( .s (signal_454), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_3301, signal_1426}), .c ({signal_3455, signal_1546}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_497 ( .s (signal_454), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_3302, signal_1425}), .c ({signal_3456, signal_1545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_498 ( .s (signal_454), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_3303, signal_1424}), .c ({signal_3457, signal_1544}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_499 ( .s (signal_454), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_3304, signal_1423}), .c ({signal_3458, signal_1543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_500 ( .s (signal_454), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_3305, signal_1422}), .c ({signal_3459, signal_1542}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_501 ( .s (signal_446), .b ({plaintext_s1[96], plaintext_s0[96]}), .a ({signal_3452, signal_1549}), .c ({signal_3628, signal_1653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_502 ( .s (signal_446), .b ({plaintext_s1[97], plaintext_s0[97]}), .a ({signal_3453, signal_1548}), .c ({signal_3630, signal_1652}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_503 ( .s (signal_446), .b ({plaintext_s1[98], plaintext_s0[98]}), .a ({signal_3454, signal_1547}), .c ({signal_3632, signal_1651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_504 ( .s (signal_446), .b ({plaintext_s1[99], plaintext_s0[99]}), .a ({signal_3455, signal_1546}), .c ({signal_3634, signal_1650}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_505 ( .s (signal_446), .b ({plaintext_s1[100], plaintext_s0[100]}), .a ({signal_3456, signal_1545}), .c ({signal_3636, signal_1649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_506 ( .s (signal_446), .b ({plaintext_s1[101], plaintext_s0[101]}), .a ({signal_3457, signal_1544}), .c ({signal_3638, signal_1648}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_507 ( .s (signal_446), .b ({plaintext_s1[102], plaintext_s0[102]}), .a ({signal_3458, signal_1543}), .c ({signal_3640, signal_1647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_508 ( .s (signal_446), .b ({plaintext_s1[103], plaintext_s0[103]}), .a ({signal_3459, signal_1542}), .c ({signal_3642, signal_1646}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_509 ( .s (signal_447), .b ({plaintext_s1[88], plaintext_s0[88]}), .a ({ciphertext_s1[80], ciphertext_s0[80]}), .c ({signal_2651, signal_1645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_510 ( .s (signal_447), .b ({plaintext_s1[89], plaintext_s0[89]}), .a ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_2654, signal_1644}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_511 ( .s (signal_447), .b ({plaintext_s1[90], plaintext_s0[90]}), .a ({ciphertext_s1[82], ciphertext_s0[82]}), .c ({signal_2657, signal_1643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_512 ( .s (signal_447), .b ({plaintext_s1[91], plaintext_s0[91]}), .a ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_2660, signal_1642}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_513 ( .s (signal_447), .b ({plaintext_s1[92], plaintext_s0[92]}), .a ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_2663, signal_1641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_514 ( .s (signal_447), .b ({plaintext_s1[93], plaintext_s0[93]}), .a ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_2666, signal_1640}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_515 ( .s (signal_447), .b ({plaintext_s1[94], plaintext_s0[94]}), .a ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_2669, signal_1639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_516 ( .s (signal_447), .b ({plaintext_s1[95], plaintext_s0[95]}), .a ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_2672, signal_1638}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_517 ( .s (signal_447), .b ({plaintext_s1[80], plaintext_s0[80]}), .a ({ciphertext_s1[72], ciphertext_s0[72]}), .c ({signal_2675, signal_1637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_518 ( .s (signal_447), .b ({plaintext_s1[81], plaintext_s0[81]}), .a ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_2678, signal_1636}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_519 ( .s (signal_447), .b ({plaintext_s1[82], plaintext_s0[82]}), .a ({ciphertext_s1[74], ciphertext_s0[74]}), .c ({signal_2681, signal_1635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_520 ( .s (signal_447), .b ({plaintext_s1[83], plaintext_s0[83]}), .a ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_2684, signal_1634}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_521 ( .s (signal_447), .b ({plaintext_s1[84], plaintext_s0[84]}), .a ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_2687, signal_1633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_522 ( .s (signal_447), .b ({plaintext_s1[85], plaintext_s0[85]}), .a ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_2690, signal_1632}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_523 ( .s (signal_447), .b ({plaintext_s1[86], plaintext_s0[86]}), .a ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_2693, signal_1631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_524 ( .s (signal_447), .b ({plaintext_s1[87], plaintext_s0[87]}), .a ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_2696, signal_1630}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_525 ( .s (signal_448), .b ({plaintext_s1[72], plaintext_s0[72]}), .a ({ciphertext_s1[64], ciphertext_s0[64]}), .c ({signal_2699, signal_1629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_526 ( .s (signal_448), .b ({plaintext_s1[73], plaintext_s0[73]}), .a ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_2702, signal_1628}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_527 ( .s (signal_448), .b ({plaintext_s1[74], plaintext_s0[74]}), .a ({ciphertext_s1[66], ciphertext_s0[66]}), .c ({signal_2705, signal_1627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_528 ( .s (signal_448), .b ({plaintext_s1[75], plaintext_s0[75]}), .a ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_2708, signal_1626}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_529 ( .s (signal_448), .b ({plaintext_s1[76], plaintext_s0[76]}), .a ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_2711, signal_1625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_530 ( .s (signal_448), .b ({plaintext_s1[77], plaintext_s0[77]}), .a ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_2714, signal_1624}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_531 ( .s (signal_448), .b ({plaintext_s1[78], plaintext_s0[78]}), .a ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_2717, signal_1623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_532 ( .s (signal_448), .b ({plaintext_s1[79], plaintext_s0[79]}), .a ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_2720, signal_1622}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_533 ( .s (signal_454), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_3290, signal_1437}), .c ({signal_3460, signal_1541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_534 ( .s (signal_454), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_3291, signal_1436}), .c ({signal_3461, signal_1540}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_535 ( .s (signal_454), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_3292, signal_1435}), .c ({signal_3462, signal_1539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_536 ( .s (signal_454), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_3293, signal_1434}), .c ({signal_3463, signal_1538}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_537 ( .s (signal_454), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_3294, signal_1433}), .c ({signal_3464, signal_1537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_538 ( .s (signal_454), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_3295, signal_1432}), .c ({signal_3465, signal_1536}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_539 ( .s (signal_454), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_3296, signal_1431}), .c ({signal_3466, signal_1535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_540 ( .s (signal_454), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_3297, signal_1430}), .c ({signal_3467, signal_1534}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_541 ( .s (signal_448), .b ({plaintext_s1[64], plaintext_s0[64]}), .a ({signal_3460, signal_1541}), .c ({signal_3644, signal_1621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_542 ( .s (signal_448), .b ({plaintext_s1[65], plaintext_s0[65]}), .a ({signal_3461, signal_1540}), .c ({signal_3646, signal_1620}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_543 ( .s (signal_448), .b ({plaintext_s1[66], plaintext_s0[66]}), .a ({signal_3462, signal_1539}), .c ({signal_3648, signal_1619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_544 ( .s (signal_448), .b ({plaintext_s1[67], plaintext_s0[67]}), .a ({signal_3463, signal_1538}), .c ({signal_3650, signal_1618}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_545 ( .s (signal_448), .b ({plaintext_s1[68], plaintext_s0[68]}), .a ({signal_3464, signal_1537}), .c ({signal_3652, signal_1617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_546 ( .s (signal_448), .b ({plaintext_s1[69], plaintext_s0[69]}), .a ({signal_3465, signal_1536}), .c ({signal_3654, signal_1616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_547 ( .s (signal_448), .b ({plaintext_s1[70], plaintext_s0[70]}), .a ({signal_3466, signal_1535}), .c ({signal_3656, signal_1615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_548 ( .s (signal_448), .b ({plaintext_s1[71], plaintext_s0[71]}), .a ({signal_3467, signal_1534}), .c ({signal_3658, signal_1614}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_549 ( .s (signal_449), .b ({plaintext_s1[56], plaintext_s0[56]}), .a ({ciphertext_s1[48], ciphertext_s0[48]}), .c ({signal_2723, signal_1613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_550 ( .s (signal_449), .b ({plaintext_s1[57], plaintext_s0[57]}), .a ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_2726, signal_1612}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_551 ( .s (signal_449), .b ({plaintext_s1[58], plaintext_s0[58]}), .a ({ciphertext_s1[50], ciphertext_s0[50]}), .c ({signal_2729, signal_1611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_552 ( .s (signal_449), .b ({plaintext_s1[59], plaintext_s0[59]}), .a ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_2732, signal_1610}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_553 ( .s (signal_449), .b ({plaintext_s1[60], plaintext_s0[60]}), .a ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_2735, signal_1609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_554 ( .s (signal_449), .b ({plaintext_s1[61], plaintext_s0[61]}), .a ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_2738, signal_1608}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_555 ( .s (signal_449), .b ({plaintext_s1[62], plaintext_s0[62]}), .a ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_2741, signal_1607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_556 ( .s (signal_449), .b ({plaintext_s1[63], plaintext_s0[63]}), .a ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_2744, signal_1606}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_557 ( .s (signal_449), .b ({plaintext_s1[48], plaintext_s0[48]}), .a ({ciphertext_s1[40], ciphertext_s0[40]}), .c ({signal_2747, signal_1605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_558 ( .s (signal_449), .b ({plaintext_s1[49], plaintext_s0[49]}), .a ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_2750, signal_1604}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_559 ( .s (signal_449), .b ({plaintext_s1[50], plaintext_s0[50]}), .a ({ciphertext_s1[42], ciphertext_s0[42]}), .c ({signal_2753, signal_1603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_560 ( .s (signal_449), .b ({plaintext_s1[51], plaintext_s0[51]}), .a ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_2756, signal_1602}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_561 ( .s (signal_449), .b ({plaintext_s1[52], plaintext_s0[52]}), .a ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_2759, signal_1601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_562 ( .s (signal_449), .b ({plaintext_s1[53], plaintext_s0[53]}), .a ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_2762, signal_1600}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_563 ( .s (signal_449), .b ({plaintext_s1[54], plaintext_s0[54]}), .a ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_2765, signal_1599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_564 ( .s (signal_449), .b ({plaintext_s1[55], plaintext_s0[55]}), .a ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_2768, signal_1598}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_565 ( .s (signal_450), .b ({plaintext_s1[40], plaintext_s0[40]}), .a ({ciphertext_s1[32], ciphertext_s0[32]}), .c ({signal_2771, signal_1597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_566 ( .s (signal_450), .b ({plaintext_s1[41], plaintext_s0[41]}), .a ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_2774, signal_1596}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_567 ( .s (signal_450), .b ({plaintext_s1[42], plaintext_s0[42]}), .a ({ciphertext_s1[34], ciphertext_s0[34]}), .c ({signal_2777, signal_1595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_568 ( .s (signal_450), .b ({plaintext_s1[43], plaintext_s0[43]}), .a ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_2780, signal_1594}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_569 ( .s (signal_450), .b ({plaintext_s1[44], plaintext_s0[44]}), .a ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_2783, signal_1593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_570 ( .s (signal_450), .b ({plaintext_s1[45], plaintext_s0[45]}), .a ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_2786, signal_1592}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_571 ( .s (signal_450), .b ({plaintext_s1[46], plaintext_s0[46]}), .a ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_2789, signal_1591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_572 ( .s (signal_450), .b ({plaintext_s1[47], plaintext_s0[47]}), .a ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_2792, signal_1590}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_573 ( .s (signal_455), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_3282, signal_1445}), .c ({signal_3468, signal_1533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_574 ( .s (signal_455), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_3283, signal_1444}), .c ({signal_3469, signal_1532}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_575 ( .s (signal_455), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_3284, signal_1443}), .c ({signal_3470, signal_1531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_576 ( .s (signal_455), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_3285, signal_1442}), .c ({signal_3471, signal_1530}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_577 ( .s (signal_455), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_3286, signal_1441}), .c ({signal_3472, signal_1529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_578 ( .s (signal_455), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_3287, signal_1440}), .c ({signal_3473, signal_1528}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_579 ( .s (signal_455), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_3288, signal_1439}), .c ({signal_3474, signal_1527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_580 ( .s (signal_455), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_3289, signal_1438}), .c ({signal_3475, signal_1526}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_581 ( .s (signal_450), .b ({plaintext_s1[32], plaintext_s0[32]}), .a ({signal_3468, signal_1533}), .c ({signal_3660, signal_1589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_582 ( .s (signal_450), .b ({plaintext_s1[33], plaintext_s0[33]}), .a ({signal_3469, signal_1532}), .c ({signal_3662, signal_1588}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_583 ( .s (signal_450), .b ({plaintext_s1[34], plaintext_s0[34]}), .a ({signal_3470, signal_1531}), .c ({signal_3664, signal_1587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_584 ( .s (signal_450), .b ({plaintext_s1[35], plaintext_s0[35]}), .a ({signal_3471, signal_1530}), .c ({signal_3666, signal_1586}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_585 ( .s (signal_450), .b ({plaintext_s1[36], plaintext_s0[36]}), .a ({signal_3472, signal_1529}), .c ({signal_3668, signal_1585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_586 ( .s (signal_450), .b ({plaintext_s1[37], plaintext_s0[37]}), .a ({signal_3473, signal_1528}), .c ({signal_3670, signal_1584}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_587 ( .s (signal_450), .b ({plaintext_s1[38], plaintext_s0[38]}), .a ({signal_3474, signal_1527}), .c ({signal_3672, signal_1583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_588 ( .s (signal_450), .b ({plaintext_s1[39], plaintext_s0[39]}), .a ({signal_3475, signal_1526}), .c ({signal_3674, signal_1582}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_589 ( .s (signal_451), .b ({plaintext_s1[24], plaintext_s0[24]}), .a ({ciphertext_s1[16], ciphertext_s0[16]}), .c ({signal_2795, signal_1581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_590 ( .s (signal_451), .b ({plaintext_s1[25], plaintext_s0[25]}), .a ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_2798, signal_1580}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_591 ( .s (signal_451), .b ({plaintext_s1[26], plaintext_s0[26]}), .a ({ciphertext_s1[18], ciphertext_s0[18]}), .c ({signal_2801, signal_1579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_592 ( .s (signal_451), .b ({plaintext_s1[27], plaintext_s0[27]}), .a ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_2804, signal_1578}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_593 ( .s (signal_451), .b ({plaintext_s1[28], plaintext_s0[28]}), .a ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_2807, signal_1577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_594 ( .s (signal_451), .b ({plaintext_s1[29], plaintext_s0[29]}), .a ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_2810, signal_1576}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_595 ( .s (signal_451), .b ({plaintext_s1[30], plaintext_s0[30]}), .a ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_2813, signal_1575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_596 ( .s (signal_451), .b ({plaintext_s1[31], plaintext_s0[31]}), .a ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_2816, signal_1574}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_597 ( .s (signal_451), .b ({plaintext_s1[16], plaintext_s0[16]}), .a ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({signal_2819, signal_1573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_598 ( .s (signal_451), .b ({plaintext_s1[17], plaintext_s0[17]}), .a ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_2822, signal_1572}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_599 ( .s (signal_451), .b ({plaintext_s1[18], plaintext_s0[18]}), .a ({ciphertext_s1[10], ciphertext_s0[10]}), .c ({signal_2825, signal_1571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_600 ( .s (signal_451), .b ({plaintext_s1[19], plaintext_s0[19]}), .a ({ciphertext_s1[11], ciphertext_s0[11]}), .c ({signal_2828, signal_1570}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_601 ( .s (signal_451), .b ({plaintext_s1[20], plaintext_s0[20]}), .a ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({signal_2831, signal_1569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_602 ( .s (signal_451), .b ({plaintext_s1[21], plaintext_s0[21]}), .a ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({signal_2834, signal_1568}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_603 ( .s (signal_451), .b ({plaintext_s1[22], plaintext_s0[22]}), .a ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_2837, signal_1567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_604 ( .s (signal_451), .b ({plaintext_s1[23], plaintext_s0[23]}), .a ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_2840, signal_1566}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_605 ( .s (signal_452), .b ({plaintext_s1[8], plaintext_s0[8]}), .a ({ciphertext_s1[0], ciphertext_s0[0]}), .c ({signal_2843, signal_1565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_606 ( .s (signal_452), .b ({plaintext_s1[9], plaintext_s0[9]}), .a ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_2846, signal_1564}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_607 ( .s (signal_452), .b ({plaintext_s1[10], plaintext_s0[10]}), .a ({ciphertext_s1[2], ciphertext_s0[2]}), .c ({signal_2849, signal_1563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_608 ( .s (signal_452), .b ({plaintext_s1[11], plaintext_s0[11]}), .a ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_2852, signal_1562}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_609 ( .s (signal_452), .b ({plaintext_s1[12], plaintext_s0[12]}), .a ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_2855, signal_1561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_610 ( .s (signal_452), .b ({plaintext_s1[13], plaintext_s0[13]}), .a ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_2858, signal_1560}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_611 ( .s (signal_452), .b ({plaintext_s1[14], plaintext_s0[14]}), .a ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_2861, signal_1559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_612 ( .s (signal_452), .b ({plaintext_s1[15], plaintext_s0[15]}), .a ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_2864, signal_1558}) ) ;
    INV_X1 cell_629 ( .A (signal_399), .ZN (signal_721) ) ;
    INV_X1 cell_630 ( .A (signal_721), .ZN (signal_722) ) ;
    INV_X1 cell_631 ( .A (signal_721), .ZN (signal_723) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_632 ( .s (signal_723), .b ({signal_3248, signal_1485}), .a ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_3278, signal_1453}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_633 ( .s (signal_722), .b ({signal_3272, signal_1484}), .a ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_3279, signal_1452}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_634 ( .s (signal_399), .b ({signal_3246, signal_1483}), .a ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_3257, signal_1451}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_635 ( .s (signal_399), .b ({signal_3271, signal_1482}), .a ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_3280, signal_1450}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_636 ( .s (signal_399), .b ({signal_3270, signal_1481}), .a ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_3281, signal_1449}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_637 ( .s (signal_399), .b ({signal_3243, signal_1480}), .a ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_3258, signal_1448}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_638 ( .s (signal_399), .b ({signal_3242, signal_1479}), .a ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_3259, signal_1447}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_639 ( .s (signal_399), .b ({signal_3241, signal_1478}), .a ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_3260, signal_1446}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_640 ( .s (signal_722), .b ({signal_3240, signal_1477}), .a ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_3282, signal_1445}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_641 ( .s (signal_722), .b ({signal_3269, signal_1476}), .a ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_3283, signal_1444}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_642 ( .s (signal_722), .b ({signal_3238, signal_1475}), .a ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_3284, signal_1443}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_643 ( .s (signal_722), .b ({signal_3268, signal_1474}), .a ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_3285, signal_1442}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_644 ( .s (signal_722), .b ({signal_3267, signal_1473}), .a ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_3286, signal_1441}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_645 ( .s (signal_722), .b ({signal_3235, signal_1472}), .a ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_3287, signal_1440}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_646 ( .s (signal_722), .b ({signal_3234, signal_1471}), .a ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_3288, signal_1439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_647 ( .s (signal_722), .b ({signal_3233, signal_1470}), .a ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_3289, signal_1438}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_648 ( .s (signal_722), .b ({signal_3232, signal_1469}), .a ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_3290, signal_1437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_649 ( .s (signal_722), .b ({signal_3266, signal_1468}), .a ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_3291, signal_1436}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_650 ( .s (signal_722), .b ({signal_3230, signal_1467}), .a ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_3292, signal_1435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_651 ( .s (signal_722), .b ({signal_3265, signal_1466}), .a ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_3293, signal_1434}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_652 ( .s (signal_723), .b ({signal_3264, signal_1465}), .a ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_3294, signal_1433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_653 ( .s (signal_723), .b ({signal_3227, signal_1464}), .a ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_3295, signal_1432}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_654 ( .s (signal_723), .b ({signal_3226, signal_1463}), .a ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_3296, signal_1431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_655 ( .s (signal_723), .b ({signal_3225, signal_1462}), .a ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_3297, signal_1430}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_656 ( .s (signal_723), .b ({signal_3224, signal_1461}), .a ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_3298, signal_1429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_657 ( .s (signal_723), .b ({signal_3263, signal_1460}), .a ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_3299, signal_1428}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_658 ( .s (signal_723), .b ({signal_3222, signal_1459}), .a ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_3300, signal_1427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_659 ( .s (signal_723), .b ({signal_3262, signal_1458}), .a ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_3301, signal_1426}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_660 ( .s (signal_723), .b ({signal_3261, signal_1457}), .a ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_3302, signal_1425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_661 ( .s (signal_723), .b ({signal_3219, signal_1456}), .a ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_3303, signal_1424}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_662 ( .s (signal_723), .b ({signal_3218, signal_1455}), .a ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_3304, signal_1423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_663 ( .s (signal_723), .b ({signal_3217, signal_1454}), .a ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_3305, signal_1422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_664 ( .a ({signal_2429, signal_765}), .b ({signal_2427, signal_1486}), .c ({signal_2430, signal_1686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_665 ( .a ({signal_2431, signal_764}), .b ({signal_2424, signal_1487}), .c ({signal_2432, signal_1687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_666 ( .a ({signal_2433, signal_763}), .b ({signal_2421, signal_1488}), .c ({signal_2434, signal_1688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_667 ( .a ({signal_2435, signal_762}), .b ({signal_2418, signal_1489}), .c ({signal_2436, signal_1689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_668 ( .a ({signal_2437, signal_761}), .b ({signal_2415, signal_1490}), .c ({signal_2438, signal_1690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_669 ( .a ({signal_2439, signal_760}), .b ({signal_2412, signal_1491}), .c ({signal_2440, signal_1691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_670 ( .a ({signal_2441, signal_759}), .b ({signal_2409, signal_1492}), .c ({signal_2442, signal_1692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_671 ( .a ({signal_2443, signal_758}), .b ({signal_2406, signal_1493}), .c ({signal_2444, signal_1693}) ) ;
    INV_X1 cell_688 ( .A (signal_732), .ZN (signal_733) ) ;
    INV_X1 cell_689 ( .A (signal_732), .ZN (signal_734) ) ;
    INV_X1 cell_690 ( .A (signal_732), .ZN (signal_735) ) ;
    INV_X1 cell_691 ( .A (signal_732), .ZN (signal_736) ) ;
    INV_X1 cell_692 ( .A (signal_732), .ZN (signal_737) ) ;
    INV_X1 cell_693 ( .A (signal_732), .ZN (signal_738) ) ;
    INV_X1 cell_694 ( .A (signal_732), .ZN (signal_739) ) ;
    INV_X1 cell_695 ( .A (signal_732), .ZN (signal_740) ) ;
    INV_X1 cell_696 ( .A (signal_393), .ZN (signal_732) ) ;
    INV_X1 cell_697 ( .A (signal_741), .ZN (signal_748) ) ;
    INV_X1 cell_698 ( .A (signal_750), .ZN (signal_756) ) ;
    INV_X1 cell_699 ( .A (signal_741), .ZN (signal_742) ) ;
    INV_X1 cell_700 ( .A (signal_750), .ZN (signal_751) ) ;
    INV_X1 cell_701 ( .A (signal_741), .ZN (signal_743) ) ;
    INV_X1 cell_702 ( .A (signal_750), .ZN (signal_752) ) ;
    INV_X1 cell_703 ( .A (signal_741), .ZN (signal_744) ) ;
    INV_X1 cell_704 ( .A (signal_750), .ZN (signal_753) ) ;
    INV_X1 cell_705 ( .A (signal_741), .ZN (signal_747) ) ;
    INV_X1 cell_706 ( .A (signal_750), .ZN (signal_755) ) ;
    INV_X1 cell_707 ( .A (signal_741), .ZN (signal_746) ) ;
    INV_X1 cell_708 ( .A (signal_750), .ZN (signal_754) ) ;
    INV_X1 cell_709 ( .A (signal_741), .ZN (signal_749) ) ;
    INV_X1 cell_710 ( .A (signal_750), .ZN (signal_757) ) ;
    INV_X1 cell_711 ( .A (signal_741), .ZN (signal_745) ) ;
    INV_X1 cell_712 ( .A (signal_394), .ZN (signal_741) ) ;
    INV_X1 cell_713 ( .A (signal_404), .ZN (signal_750) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_714 ( .s (signal_751), .b ({signal_2406, signal_1493}), .a ({signal_4020, signal_767}), .c ({signal_4156, signal_766}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_715 ( .s (signal_742), .b ({signal_3941, signal_1933}), .a ({signal_2914, signal_1877}), .c ({signal_4020, signal_767}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_718 ( .s (signal_751), .b ({signal_2409, signal_1492}), .a ({signal_4021, signal_770}), .c ({signal_4157, signal_769}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_719 ( .s (signal_742), .b ({signal_3943, signal_1932}), .a ({signal_2917, signal_1876}), .c ({signal_4021, signal_770}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_722 ( .s (signal_751), .b ({signal_2412, signal_1491}), .a ({signal_4022, signal_773}), .c ({signal_4158, signal_772}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_723 ( .s (signal_742), .b ({signal_3945, signal_1931}), .a ({signal_2920, signal_1875}), .c ({signal_4022, signal_773}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_726 ( .s (signal_751), .b ({signal_2415, signal_1490}), .a ({signal_4023, signal_776}), .c ({signal_4159, signal_775}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_727 ( .s (signal_742), .b ({signal_3947, signal_1930}), .a ({signal_2923, signal_1874}), .c ({signal_4023, signal_776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_730 ( .s (signal_751), .b ({signal_2418, signal_1489}), .a ({signal_4024, signal_779}), .c ({signal_4160, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_731 ( .s (signal_742), .b ({signal_3949, signal_1929}), .a ({signal_2926, signal_1873}), .c ({signal_4024, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_734 ( .s (signal_751), .b ({signal_2421, signal_1488}), .a ({signal_4025, signal_782}), .c ({signal_4161, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_735 ( .s (signal_742), .b ({signal_3951, signal_1928}), .a ({signal_2929, signal_1872}), .c ({signal_4025, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_738 ( .s (signal_751), .b ({signal_2424, signal_1487}), .a ({signal_4026, signal_785}), .c ({signal_4162, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_739 ( .s (signal_742), .b ({signal_3953, signal_1927}), .a ({signal_2932, signal_1871}), .c ({signal_4026, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_742 ( .s (signal_751), .b ({signal_2427, signal_1486}), .a ({signal_4027, signal_788}), .c ({signal_4163, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_743 ( .s (signal_742), .b ({signal_3955, signal_1926}), .a ({signal_2935, signal_1870}), .c ({signal_4027, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_746 ( .s (signal_751), .b ({signal_2443, signal_758}), .a ({signal_3306, signal_791}), .c ({signal_4028, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_747 ( .s (signal_742), .b ({signal_2867, signal_1925}), .a ({signal_2938, signal_1861}), .c ({signal_3306, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_750 ( .s (signal_751), .b ({signal_2441, signal_759}), .a ({signal_3307, signal_794}), .c ({signal_4029, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_751 ( .s (signal_742), .b ({signal_2870, signal_1924}), .a ({signal_2941, signal_1860}), .c ({signal_3307, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_754 ( .s (signal_751), .b ({signal_2439, signal_760}), .a ({signal_3308, signal_797}), .c ({signal_4030, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_755 ( .s (signal_742), .b ({signal_2873, signal_1923}), .a ({signal_2944, signal_1859}), .c ({signal_3308, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_758 ( .s (signal_751), .b ({signal_2437, signal_761}), .a ({signal_3309, signal_800}), .c ({signal_4031, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_759 ( .s (signal_742), .b ({signal_2876, signal_1922}), .a ({signal_2947, signal_1858}), .c ({signal_3309, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_762 ( .s (signal_751), .b ({signal_2435, signal_762}), .a ({signal_3310, signal_803}), .c ({signal_4032, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_763 ( .s (signal_742), .b ({signal_2879, signal_1921}), .a ({signal_2950, signal_1857}), .c ({signal_3310, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_766 ( .s (signal_751), .b ({signal_2433, signal_763}), .a ({signal_3311, signal_806}), .c ({signal_4033, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_767 ( .s (signal_742), .b ({signal_2882, signal_1920}), .a ({signal_2953, signal_1856}), .c ({signal_3311, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_770 ( .s (signal_751), .b ({signal_2431, signal_764}), .a ({signal_3312, signal_809}), .c ({signal_4034, signal_808}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_771 ( .s (signal_742), .b ({signal_2885, signal_1919}), .a ({signal_2956, signal_1855}), .c ({signal_3312, signal_809}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_774 ( .s (signal_751), .b ({signal_2429, signal_765}), .a ({signal_3313, signal_812}), .c ({signal_4035, signal_811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_775 ( .s (signal_742), .b ({signal_2888, signal_1918}), .a ({signal_2959, signal_1854}), .c ({signal_3313, signal_812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_778 ( .s (signal_752), .b ({signal_2866, signal_1909}), .a ({signal_3314, signal_815}), .c ({signal_4036, signal_814}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_779 ( .s (signal_743), .b ({signal_2891, signal_1917}), .a ({signal_2962, signal_1845}), .c ({signal_3314, signal_815}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_782 ( .s (signal_752), .b ({signal_2869, signal_1908}), .a ({signal_3315, signal_818}), .c ({signal_4037, signal_817}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_783 ( .s (signal_743), .b ({signal_2894, signal_1916}), .a ({signal_2965, signal_1844}), .c ({signal_3315, signal_818}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_786 ( .s (signal_752), .b ({signal_2872, signal_1907}), .a ({signal_3316, signal_821}), .c ({signal_4038, signal_820}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_787 ( .s (signal_743), .b ({signal_2897, signal_1915}), .a ({signal_2968, signal_1843}), .c ({signal_3316, signal_821}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_790 ( .s (signal_752), .b ({signal_2875, signal_1906}), .a ({signal_3317, signal_824}), .c ({signal_4039, signal_823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_791 ( .s (signal_743), .b ({signal_2900, signal_1914}), .a ({signal_2971, signal_1842}), .c ({signal_3317, signal_824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_794 ( .s (signal_752), .b ({signal_2878, signal_1905}), .a ({signal_3318, signal_827}), .c ({signal_4040, signal_826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_795 ( .s (signal_743), .b ({signal_2903, signal_1913}), .a ({signal_2974, signal_1841}), .c ({signal_3318, signal_827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_798 ( .s (signal_752), .b ({signal_2881, signal_1904}), .a ({signal_3319, signal_830}), .c ({signal_4041, signal_829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_799 ( .s (signal_743), .b ({signal_2906, signal_1912}), .a ({signal_2977, signal_1840}), .c ({signal_3319, signal_830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_802 ( .s (signal_752), .b ({signal_2884, signal_1903}), .a ({signal_3320, signal_833}), .c ({signal_4042, signal_832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_803 ( .s (signal_743), .b ({signal_2909, signal_1911}), .a ({signal_2980, signal_1839}), .c ({signal_3320, signal_833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_806 ( .s (signal_752), .b ({signal_2887, signal_1902}), .a ({signal_3321, signal_836}), .c ({signal_4043, signal_835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_807 ( .s (signal_743), .b ({signal_2912, signal_1910}), .a ({signal_2983, signal_1838}), .c ({signal_3321, signal_836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_810 ( .s (signal_752), .b ({signal_2890, signal_1893}), .a ({signal_3322, signal_839}), .c ({signal_4044, signal_838}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_811 ( .s (signal_743), .b ({signal_2915, signal_1901}), .a ({signal_2986, signal_1509}), .c ({signal_3322, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_814 ( .s (signal_752), .b ({signal_2893, signal_1892}), .a ({signal_3323, signal_842}), .c ({signal_4045, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_815 ( .s (signal_743), .b ({signal_2918, signal_1900}), .a ({signal_2989, signal_1508}), .c ({signal_3323, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_818 ( .s (signal_752), .b ({signal_2896, signal_1891}), .a ({signal_3324, signal_845}), .c ({signal_4046, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_819 ( .s (signal_743), .b ({signal_2921, signal_1899}), .a ({signal_2992, signal_1507}), .c ({signal_3324, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_822 ( .s (signal_752), .b ({signal_2899, signal_1890}), .a ({signal_3325, signal_848}), .c ({signal_4047, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_823 ( .s (signal_743), .b ({signal_2924, signal_1898}), .a ({signal_2995, signal_1506}), .c ({signal_3325, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_826 ( .s (signal_752), .b ({signal_2902, signal_1889}), .a ({signal_3326, signal_851}), .c ({signal_4048, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_827 ( .s (signal_743), .b ({signal_2927, signal_1897}), .a ({signal_2998, signal_1505}), .c ({signal_3326, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_830 ( .s (signal_752), .b ({signal_2905, signal_1888}), .a ({signal_3327, signal_854}), .c ({signal_4049, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_831 ( .s (signal_743), .b ({signal_2930, signal_1896}), .a ({signal_3001, signal_1504}), .c ({signal_3327, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_834 ( .s (signal_752), .b ({signal_2908, signal_1887}), .a ({signal_3328, signal_857}), .c ({signal_4050, signal_856}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_835 ( .s (signal_743), .b ({signal_2933, signal_1895}), .a ({signal_3004, signal_1503}), .c ({signal_3328, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_838 ( .s (signal_752), .b ({signal_2911, signal_1886}), .a ({signal_3329, signal_860}), .c ({signal_4051, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_839 ( .s (signal_743), .b ({signal_2936, signal_1894}), .a ({signal_3007, signal_1502}), .c ({signal_3329, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_842 ( .s (signal_753), .b ({signal_2914, signal_1877}), .a ({signal_3330, signal_863}), .c ({signal_4052, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_843 ( .s (signal_744), .b ({signal_2939, signal_1885}), .a ({signal_3010, signal_1821}), .c ({signal_3330, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_846 ( .s (signal_753), .b ({signal_2917, signal_1876}), .a ({signal_3331, signal_866}), .c ({signal_4053, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_847 ( .s (signal_744), .b ({signal_2942, signal_1884}), .a ({signal_3013, signal_1820}), .c ({signal_3331, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_850 ( .s (signal_753), .b ({signal_2920, signal_1875}), .a ({signal_3332, signal_869}), .c ({signal_4054, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_851 ( .s (signal_744), .b ({signal_2945, signal_1883}), .a ({signal_3016, signal_1819}), .c ({signal_3332, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_854 ( .s (signal_753), .b ({signal_2923, signal_1874}), .a ({signal_3333, signal_872}), .c ({signal_4055, signal_871}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_855 ( .s (signal_744), .b ({signal_2948, signal_1882}), .a ({signal_3019, signal_1818}), .c ({signal_3333, signal_872}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_858 ( .s (signal_753), .b ({signal_2926, signal_1873}), .a ({signal_3334, signal_875}), .c ({signal_4056, signal_874}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_859 ( .s (signal_744), .b ({signal_2951, signal_1881}), .a ({signal_3022, signal_1817}), .c ({signal_3334, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_862 ( .s (signal_753), .b ({signal_2929, signal_1872}), .a ({signal_3335, signal_878}), .c ({signal_4057, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_863 ( .s (signal_744), .b ({signal_2954, signal_1880}), .a ({signal_3025, signal_1816}), .c ({signal_3335, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_866 ( .s (signal_753), .b ({signal_2932, signal_1871}), .a ({signal_3336, signal_881}), .c ({signal_4058, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_867 ( .s (signal_744), .b ({signal_2957, signal_1879}), .a ({signal_3028, signal_1815}), .c ({signal_3336, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_870 ( .s (signal_753), .b ({signal_2935, signal_1870}), .a ({signal_3337, signal_884}), .c ({signal_4059, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_871 ( .s (signal_744), .b ({signal_2960, signal_1878}), .a ({signal_3031, signal_1814}), .c ({signal_3337, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_874 ( .s (signal_753), .b ({signal_2938, signal_1861}), .a ({signal_3338, signal_887}), .c ({signal_4060, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_875 ( .s (signal_744), .b ({signal_2963, signal_1869}), .a ({signal_3034, signal_1805}), .c ({signal_3338, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_878 ( .s (signal_753), .b ({signal_2941, signal_1860}), .a ({signal_3339, signal_890}), .c ({signal_4061, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_879 ( .s (signal_744), .b ({signal_2966, signal_1868}), .a ({signal_3037, signal_1804}), .c ({signal_3339, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_882 ( .s (signal_753), .b ({signal_2944, signal_1859}), .a ({signal_3340, signal_893}), .c ({signal_4062, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_883 ( .s (signal_744), .b ({signal_2969, signal_1867}), .a ({signal_3040, signal_1803}), .c ({signal_3340, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_886 ( .s (signal_753), .b ({signal_2947, signal_1858}), .a ({signal_3341, signal_896}), .c ({signal_4063, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_887 ( .s (signal_744), .b ({signal_2972, signal_1866}), .a ({signal_3043, signal_1802}), .c ({signal_3341, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_890 ( .s (signal_753), .b ({signal_2950, signal_1857}), .a ({signal_3342, signal_899}), .c ({signal_4064, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_891 ( .s (signal_744), .b ({signal_2975, signal_1865}), .a ({signal_3046, signal_1801}), .c ({signal_3342, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_894 ( .s (signal_753), .b ({signal_2953, signal_1856}), .a ({signal_3343, signal_902}), .c ({signal_4065, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_895 ( .s (signal_744), .b ({signal_2978, signal_1864}), .a ({signal_3049, signal_1800}), .c ({signal_3343, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_898 ( .s (signal_753), .b ({signal_2956, signal_1855}), .a ({signal_3344, signal_905}), .c ({signal_4066, signal_904}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_899 ( .s (signal_744), .b ({signal_2981, signal_1863}), .a ({signal_3052, signal_1799}), .c ({signal_3344, signal_905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_902 ( .s (signal_753), .b ({signal_2959, signal_1854}), .a ({signal_3345, signal_908}), .c ({signal_4067, signal_907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_903 ( .s (signal_744), .b ({signal_2984, signal_1862}), .a ({signal_3055, signal_1798}), .c ({signal_3345, signal_908}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_906 ( .s (signal_404), .b ({signal_2962, signal_1845}), .a ({signal_3346, signal_911}), .c ({signal_3675, signal_910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_907 ( .s (signal_745), .b ({signal_2987, signal_1853}), .a ({signal_3058, signal_1789}), .c ({signal_3346, signal_911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_910 ( .s (signal_404), .b ({signal_2965, signal_1844}), .a ({signal_3347, signal_914}), .c ({signal_3676, signal_913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_911 ( .s (signal_745), .b ({signal_2990, signal_1852}), .a ({signal_3061, signal_1788}), .c ({signal_3347, signal_914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_914 ( .s (signal_404), .b ({signal_2968, signal_1843}), .a ({signal_3348, signal_917}), .c ({signal_3677, signal_916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_915 ( .s (signal_745), .b ({signal_2993, signal_1851}), .a ({signal_3064, signal_1787}), .c ({signal_3348, signal_917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_918 ( .s (signal_404), .b ({signal_2971, signal_1842}), .a ({signal_3349, signal_920}), .c ({signal_3678, signal_919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_919 ( .s (signal_745), .b ({signal_2996, signal_1850}), .a ({signal_3067, signal_1786}), .c ({signal_3349, signal_920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_922 ( .s (signal_404), .b ({signal_2974, signal_1841}), .a ({signal_3350, signal_923}), .c ({signal_3679, signal_922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_923 ( .s (signal_745), .b ({signal_2999, signal_1849}), .a ({signal_3070, signal_1785}), .c ({signal_3350, signal_923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_926 ( .s (signal_404), .b ({signal_2977, signal_1840}), .a ({signal_3351, signal_926}), .c ({signal_3680, signal_925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_927 ( .s (signal_745), .b ({signal_3002, signal_1848}), .a ({signal_3073, signal_1784}), .c ({signal_3351, signal_926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_930 ( .s (signal_404), .b ({signal_2980, signal_1839}), .a ({signal_3352, signal_929}), .c ({signal_3681, signal_928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_931 ( .s (signal_745), .b ({signal_3005, signal_1847}), .a ({signal_3076, signal_1783}), .c ({signal_3352, signal_929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_934 ( .s (signal_404), .b ({signal_2983, signal_1838}), .a ({signal_3353, signal_932}), .c ({signal_3682, signal_931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_935 ( .s (signal_745), .b ({signal_3008, signal_1846}), .a ({signal_3079, signal_1782}), .c ({signal_3353, signal_932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_938 ( .s (signal_404), .b ({signal_2986, signal_1509}), .a ({signal_3354, signal_935}), .c ({signal_3683, signal_934}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_939 ( .s (signal_745), .b ({signal_3011, signal_1837}), .a ({signal_3082, signal_1773}), .c ({signal_3354, signal_935}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_942 ( .s (signal_404), .b ({signal_2989, signal_1508}), .a ({signal_3355, signal_938}), .c ({signal_3684, signal_937}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_943 ( .s (signal_745), .b ({signal_3014, signal_1836}), .a ({signal_3085, signal_1772}), .c ({signal_3355, signal_938}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_946 ( .s (signal_404), .b ({signal_2992, signal_1507}), .a ({signal_3356, signal_941}), .c ({signal_3685, signal_940}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_947 ( .s (signal_745), .b ({signal_3017, signal_1835}), .a ({signal_3088, signal_1771}), .c ({signal_3356, signal_941}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_950 ( .s (signal_404), .b ({signal_2995, signal_1506}), .a ({signal_3357, signal_944}), .c ({signal_3686, signal_943}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_951 ( .s (signal_745), .b ({signal_3020, signal_1834}), .a ({signal_3091, signal_1770}), .c ({signal_3357, signal_944}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_954 ( .s (signal_404), .b ({signal_2998, signal_1505}), .a ({signal_3358, signal_947}), .c ({signal_3687, signal_946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_955 ( .s (signal_745), .b ({signal_3023, signal_1833}), .a ({signal_3094, signal_1769}), .c ({signal_3358, signal_947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_958 ( .s (signal_404), .b ({signal_3001, signal_1504}), .a ({signal_3359, signal_950}), .c ({signal_3688, signal_949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_959 ( .s (signal_745), .b ({signal_3026, signal_1832}), .a ({signal_3097, signal_1768}), .c ({signal_3359, signal_950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_962 ( .s (signal_404), .b ({signal_3004, signal_1503}), .a ({signal_3360, signal_953}), .c ({signal_3689, signal_952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_963 ( .s (signal_745), .b ({signal_3029, signal_1831}), .a ({signal_3100, signal_1767}), .c ({signal_3360, signal_953}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_966 ( .s (signal_404), .b ({signal_3007, signal_1502}), .a ({signal_3361, signal_956}), .c ({signal_3690, signal_955}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_967 ( .s (signal_745), .b ({signal_3032, signal_1830}), .a ({signal_3103, signal_1766}), .c ({signal_3361, signal_956}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_970 ( .s (signal_754), .b ({signal_3010, signal_1821}), .a ({signal_3362, signal_959}), .c ({signal_4068, signal_958}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_971 ( .s (signal_746), .b ({signal_3035, signal_1829}), .a ({signal_3106, signal_1749}), .c ({signal_3362, signal_959}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_974 ( .s (signal_754), .b ({signal_3013, signal_1820}), .a ({signal_3363, signal_962}), .c ({signal_4069, signal_961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_975 ( .s (signal_746), .b ({signal_3038, signal_1828}), .a ({signal_3109, signal_1748}), .c ({signal_3363, signal_962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_978 ( .s (signal_754), .b ({signal_3016, signal_1819}), .a ({signal_3364, signal_965}), .c ({signal_4070, signal_964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_979 ( .s (signal_746), .b ({signal_3041, signal_1827}), .a ({signal_3112, signal_1747}), .c ({signal_3364, signal_965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_982 ( .s (signal_754), .b ({signal_3019, signal_1818}), .a ({signal_3365, signal_968}), .c ({signal_4071, signal_967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_983 ( .s (signal_746), .b ({signal_3044, signal_1826}), .a ({signal_3115, signal_1746}), .c ({signal_3365, signal_968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_986 ( .s (signal_754), .b ({signal_3022, signal_1817}), .a ({signal_3366, signal_971}), .c ({signal_4072, signal_970}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_987 ( .s (signal_746), .b ({signal_3047, signal_1825}), .a ({signal_3118, signal_1745}), .c ({signal_3366, signal_971}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_990 ( .s (signal_754), .b ({signal_3025, signal_1816}), .a ({signal_3367, signal_974}), .c ({signal_4073, signal_973}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_991 ( .s (signal_746), .b ({signal_3050, signal_1824}), .a ({signal_3121, signal_1744}), .c ({signal_3367, signal_974}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_994 ( .s (signal_754), .b ({signal_3028, signal_1815}), .a ({signal_3368, signal_977}), .c ({signal_4074, signal_976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_995 ( .s (signal_746), .b ({signal_3053, signal_1823}), .a ({signal_3124, signal_1743}), .c ({signal_3368, signal_977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_998 ( .s (signal_754), .b ({signal_3031, signal_1814}), .a ({signal_3369, signal_980}), .c ({signal_4075, signal_979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_999 ( .s (signal_746), .b ({signal_3056, signal_1822}), .a ({signal_3127, signal_1742}), .c ({signal_3369, signal_980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1002 ( .s (signal_754), .b ({signal_3034, signal_1805}), .a ({signal_3370, signal_983}), .c ({signal_4076, signal_982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1003 ( .s (signal_746), .b ({signal_3059, signal_1813}), .a ({signal_3130, signal_1733}), .c ({signal_3370, signal_983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1006 ( .s (signal_754), .b ({signal_3037, signal_1804}), .a ({signal_3371, signal_986}), .c ({signal_4077, signal_985}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1007 ( .s (signal_746), .b ({signal_3062, signal_1812}), .a ({signal_3133, signal_1732}), .c ({signal_3371, signal_986}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1010 ( .s (signal_754), .b ({signal_3040, signal_1803}), .a ({signal_3372, signal_989}), .c ({signal_4078, signal_988}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1011 ( .s (signal_746), .b ({signal_3065, signal_1811}), .a ({signal_3136, signal_1731}), .c ({signal_3372, signal_989}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1014 ( .s (signal_754), .b ({signal_3043, signal_1802}), .a ({signal_3373, signal_992}), .c ({signal_4079, signal_991}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1015 ( .s (signal_746), .b ({signal_3068, signal_1810}), .a ({signal_3139, signal_1730}), .c ({signal_3373, signal_992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1018 ( .s (signal_754), .b ({signal_3046, signal_1801}), .a ({signal_3374, signal_995}), .c ({signal_4080, signal_994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1019 ( .s (signal_746), .b ({signal_3071, signal_1809}), .a ({signal_3142, signal_1729}), .c ({signal_3374, signal_995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1022 ( .s (signal_754), .b ({signal_3049, signal_1800}), .a ({signal_3375, signal_998}), .c ({signal_4081, signal_997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1023 ( .s (signal_746), .b ({signal_3074, signal_1808}), .a ({signal_3145, signal_1728}), .c ({signal_3375, signal_998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1026 ( .s (signal_754), .b ({signal_3052, signal_1799}), .a ({signal_3376, signal_1001}), .c ({signal_4082, signal_1000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1027 ( .s (signal_746), .b ({signal_3077, signal_1807}), .a ({signal_3148, signal_1727}), .c ({signal_3376, signal_1001}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1030 ( .s (signal_754), .b ({signal_3055, signal_1798}), .a ({signal_3377, signal_1004}), .c ({signal_4083, signal_1003}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1031 ( .s (signal_746), .b ({signal_3080, signal_1806}), .a ({signal_3151, signal_1726}), .c ({signal_3377, signal_1004}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1034 ( .s (signal_755), .b ({signal_3058, signal_1789}), .a ({signal_3378, signal_1007}), .c ({signal_4084, signal_1006}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1035 ( .s (signal_747), .b ({signal_3083, signal_1797}), .a ({signal_3154, signal_1717}), .c ({signal_3378, signal_1007}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1038 ( .s (signal_755), .b ({signal_3061, signal_1788}), .a ({signal_3379, signal_1010}), .c ({signal_4085, signal_1009}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1039 ( .s (signal_747), .b ({signal_3086, signal_1796}), .a ({signal_3157, signal_1716}), .c ({signal_3379, signal_1010}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1042 ( .s (signal_755), .b ({signal_3064, signal_1787}), .a ({signal_3380, signal_1013}), .c ({signal_4086, signal_1012}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1043 ( .s (signal_747), .b ({signal_3089, signal_1795}), .a ({signal_3160, signal_1715}), .c ({signal_3380, signal_1013}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1046 ( .s (signal_755), .b ({signal_3067, signal_1786}), .a ({signal_3381, signal_1016}), .c ({signal_4087, signal_1015}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1047 ( .s (signal_747), .b ({signal_3092, signal_1794}), .a ({signal_3163, signal_1714}), .c ({signal_3381, signal_1016}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1050 ( .s (signal_755), .b ({signal_3070, signal_1785}), .a ({signal_3382, signal_1019}), .c ({signal_4088, signal_1018}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1051 ( .s (signal_747), .b ({signal_3095, signal_1793}), .a ({signal_3166, signal_1713}), .c ({signal_3382, signal_1019}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1054 ( .s (signal_755), .b ({signal_3073, signal_1784}), .a ({signal_3383, signal_1022}), .c ({signal_4089, signal_1021}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1055 ( .s (signal_747), .b ({signal_3098, signal_1792}), .a ({signal_3169, signal_1712}), .c ({signal_3383, signal_1022}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1058 ( .s (signal_755), .b ({signal_3076, signal_1783}), .a ({signal_3384, signal_1025}), .c ({signal_4090, signal_1024}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1059 ( .s (signal_747), .b ({signal_3101, signal_1791}), .a ({signal_3172, signal_1711}), .c ({signal_3384, signal_1025}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1062 ( .s (signal_755), .b ({signal_3079, signal_1782}), .a ({signal_3385, signal_1028}), .c ({signal_4091, signal_1027}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1063 ( .s (signal_747), .b ({signal_3104, signal_1790}), .a ({signal_3175, signal_1710}), .c ({signal_3385, signal_1028}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1066 ( .s (signal_755), .b ({signal_3082, signal_1773}), .a ({signal_3386, signal_1031}), .c ({signal_4092, signal_1030}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1067 ( .s (signal_747), .b ({signal_3107, signal_1781}), .a ({signal_3178, signal_1701}), .c ({signal_3386, signal_1031}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1070 ( .s (signal_755), .b ({signal_3085, signal_1772}), .a ({signal_3387, signal_1034}), .c ({signal_4093, signal_1033}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1071 ( .s (signal_747), .b ({signal_3110, signal_1780}), .a ({signal_3181, signal_1700}), .c ({signal_3387, signal_1034}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1074 ( .s (signal_755), .b ({signal_3088, signal_1771}), .a ({signal_3388, signal_1037}), .c ({signal_4094, signal_1036}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1075 ( .s (signal_747), .b ({signal_3113, signal_1779}), .a ({signal_3184, signal_1699}), .c ({signal_3388, signal_1037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1078 ( .s (signal_755), .b ({signal_3091, signal_1770}), .a ({signal_3389, signal_1040}), .c ({signal_4095, signal_1039}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1079 ( .s (signal_747), .b ({signal_3116, signal_1778}), .a ({signal_3187, signal_1698}), .c ({signal_3389, signal_1040}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1082 ( .s (signal_755), .b ({signal_3094, signal_1769}), .a ({signal_3390, signal_1043}), .c ({signal_4096, signal_1042}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1083 ( .s (signal_747), .b ({signal_3119, signal_1777}), .a ({signal_3190, signal_1697}), .c ({signal_3390, signal_1043}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1086 ( .s (signal_755), .b ({signal_3097, signal_1768}), .a ({signal_3391, signal_1046}), .c ({signal_4097, signal_1045}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1087 ( .s (signal_747), .b ({signal_3122, signal_1776}), .a ({signal_3193, signal_1696}), .c ({signal_3391, signal_1046}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1090 ( .s (signal_755), .b ({signal_3100, signal_1767}), .a ({signal_3392, signal_1049}), .c ({signal_4098, signal_1048}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1091 ( .s (signal_747), .b ({signal_3125, signal_1775}), .a ({signal_3196, signal_1695}), .c ({signal_3392, signal_1049}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1094 ( .s (signal_755), .b ({signal_3103, signal_1766}), .a ({signal_3393, signal_1052}), .c ({signal_4099, signal_1051}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1095 ( .s (signal_747), .b ({signal_3128, signal_1774}), .a ({signal_3199, signal_1694}), .c ({signal_3393, signal_1052}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1130 ( .s (signal_756), .b ({signal_3130, signal_1733}), .a ({signal_3394, signal_1079}), .c ({signal_4100, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1131 ( .s (signal_748), .b ({signal_3155, signal_1741}), .a ({signal_2443, signal_758}), .c ({signal_3394, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1134 ( .s (signal_756), .b ({signal_3133, signal_1732}), .a ({signal_3395, signal_1082}), .c ({signal_4101, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1135 ( .s (signal_748), .b ({signal_3158, signal_1740}), .a ({signal_2441, signal_759}), .c ({signal_3395, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1138 ( .s (signal_756), .b ({signal_3136, signal_1731}), .a ({signal_3396, signal_1085}), .c ({signal_4102, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1139 ( .s (signal_748), .b ({signal_3161, signal_1739}), .a ({signal_2439, signal_760}), .c ({signal_3396, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1142 ( .s (signal_756), .b ({signal_3139, signal_1730}), .a ({signal_3397, signal_1088}), .c ({signal_4103, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1143 ( .s (signal_748), .b ({signal_3164, signal_1738}), .a ({signal_2437, signal_761}), .c ({signal_3397, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1146 ( .s (signal_756), .b ({signal_3142, signal_1729}), .a ({signal_3398, signal_1091}), .c ({signal_4104, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1147 ( .s (signal_748), .b ({signal_3167, signal_1737}), .a ({signal_2435, signal_762}), .c ({signal_3398, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1150 ( .s (signal_756), .b ({signal_3145, signal_1728}), .a ({signal_3399, signal_1094}), .c ({signal_4105, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1151 ( .s (signal_748), .b ({signal_3170, signal_1736}), .a ({signal_2433, signal_763}), .c ({signal_3399, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1154 ( .s (signal_756), .b ({signal_3148, signal_1727}), .a ({signal_3400, signal_1097}), .c ({signal_4106, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1155 ( .s (signal_748), .b ({signal_3173, signal_1735}), .a ({signal_2431, signal_764}), .c ({signal_3400, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1158 ( .s (signal_756), .b ({signal_3151, signal_1726}), .a ({signal_3401, signal_1100}), .c ({signal_4107, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1159 ( .s (signal_748), .b ({signal_3176, signal_1734}), .a ({signal_2429, signal_765}), .c ({signal_3401, signal_1100}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1162 ( .s (signal_757), .b ({signal_3154, signal_1717}), .a ({signal_3402, signal_1103}), .c ({signal_4108, signal_1102}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1163 ( .s (signal_749), .b ({signal_3179, signal_1725}), .a ({signal_2866, signal_1909}), .c ({signal_3402, signal_1103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1166 ( .s (signal_757), .b ({signal_3157, signal_1716}), .a ({signal_3403, signal_1106}), .c ({signal_4109, signal_1105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1167 ( .s (signal_749), .b ({signal_3182, signal_1724}), .a ({signal_2869, signal_1908}), .c ({signal_3403, signal_1106}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1170 ( .s (signal_757), .b ({signal_3160, signal_1715}), .a ({signal_3404, signal_1109}), .c ({signal_4110, signal_1108}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1171 ( .s (signal_749), .b ({signal_3185, signal_1723}), .a ({signal_2872, signal_1907}), .c ({signal_3404, signal_1109}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1174 ( .s (signal_757), .b ({signal_3163, signal_1714}), .a ({signal_3405, signal_1112}), .c ({signal_4111, signal_1111}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1175 ( .s (signal_749), .b ({signal_3188, signal_1722}), .a ({signal_2875, signal_1906}), .c ({signal_3405, signal_1112}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1178 ( .s (signal_757), .b ({signal_3166, signal_1713}), .a ({signal_3406, signal_1115}), .c ({signal_4112, signal_1114}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1179 ( .s (signal_749), .b ({signal_3191, signal_1721}), .a ({signal_2878, signal_1905}), .c ({signal_3406, signal_1115}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1182 ( .s (signal_757), .b ({signal_3169, signal_1712}), .a ({signal_3407, signal_1118}), .c ({signal_4113, signal_1117}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1183 ( .s (signal_749), .b ({signal_3194, signal_1720}), .a ({signal_2881, signal_1904}), .c ({signal_3407, signal_1118}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1186 ( .s (signal_757), .b ({signal_3172, signal_1711}), .a ({signal_3408, signal_1121}), .c ({signal_4114, signal_1120}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1187 ( .s (signal_749), .b ({signal_3197, signal_1719}), .a ({signal_2884, signal_1903}), .c ({signal_3408, signal_1121}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1190 ( .s (signal_757), .b ({signal_3175, signal_1710}), .a ({signal_3409, signal_1124}), .c ({signal_4115, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1191 ( .s (signal_749), .b ({signal_3200, signal_1718}), .a ({signal_2887, signal_1902}), .c ({signal_3409, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1194 ( .s (signal_757), .b ({signal_3178, signal_1701}), .a ({signal_3410, signal_1127}), .c ({signal_4116, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1195 ( .s (signal_749), .b ({signal_3202, signal_1709}), .a ({signal_2890, signal_1893}), .c ({signal_3410, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1198 ( .s (signal_757), .b ({signal_3181, signal_1700}), .a ({signal_3411, signal_1130}), .c ({signal_4117, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1199 ( .s (signal_749), .b ({signal_3204, signal_1708}), .a ({signal_2893, signal_1892}), .c ({signal_3411, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1202 ( .s (signal_757), .b ({signal_3184, signal_1699}), .a ({signal_3412, signal_1133}), .c ({signal_4118, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1203 ( .s (signal_749), .b ({signal_3206, signal_1707}), .a ({signal_2896, signal_1891}), .c ({signal_3412, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1206 ( .s (signal_757), .b ({signal_3187, signal_1698}), .a ({signal_3413, signal_1136}), .c ({signal_4119, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1207 ( .s (signal_749), .b ({signal_3208, signal_1706}), .a ({signal_2899, signal_1890}), .c ({signal_3413, signal_1136}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1210 ( .s (signal_757), .b ({signal_3190, signal_1697}), .a ({signal_3414, signal_1139}), .c ({signal_4120, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1211 ( .s (signal_749), .b ({signal_3210, signal_1705}), .a ({signal_2902, signal_1889}), .c ({signal_3414, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1214 ( .s (signal_757), .b ({signal_3193, signal_1696}), .a ({signal_3415, signal_1142}), .c ({signal_4121, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1215 ( .s (signal_749), .b ({signal_3212, signal_1704}), .a ({signal_2905, signal_1888}), .c ({signal_3415, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1218 ( .s (signal_757), .b ({signal_3196, signal_1695}), .a ({signal_3416, signal_1145}), .c ({signal_4122, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1219 ( .s (signal_749), .b ({signal_3214, signal_1703}), .a ({signal_2908, signal_1887}), .c ({signal_3416, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1222 ( .s (signal_757), .b ({signal_3199, signal_1694}), .a ({signal_3417, signal_1148}), .c ({signal_4123, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1223 ( .s (signal_749), .b ({signal_3216, signal_1702}), .a ({signal_2911, signal_1886}), .c ({signal_3417, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1226 ( .s (signal_400), .b ({signal_2443, signal_758}), .a ({signal_2444, signal_1693}), .c ({signal_3691, signal_1685}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1227 ( .s (signal_400), .b ({signal_2441, signal_759}), .a ({signal_2442, signal_1692}), .c ({signal_3692, signal_1684}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1228 ( .s (signal_400), .b ({signal_2439, signal_760}), .a ({signal_2440, signal_1691}), .c ({signal_3693, signal_1683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1229 ( .s (signal_400), .b ({signal_2437, signal_761}), .a ({signal_2438, signal_1690}), .c ({signal_3694, signal_1682}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1230 ( .s (signal_400), .b ({signal_2435, signal_762}), .a ({signal_2436, signal_1689}), .c ({signal_3695, signal_1681}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1231 ( .s (signal_400), .b ({signal_2433, signal_763}), .a ({signal_2434, signal_1688}), .c ({signal_3696, signal_1680}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1232 ( .s (signal_400), .b ({signal_2431, signal_764}), .a ({signal_2432, signal_1687}), .c ({signal_3697, signal_1679}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1233 ( .s (signal_400), .b ({signal_2429, signal_765}), .a ({signal_2430, signal_1686}), .c ({signal_3698, signal_1678}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1234 ( .s (signal_733), .b ({key_s1[120], key_s0[120]}), .a ({signal_3691, signal_1685}), .c ({signal_3941, signal_1933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1235 ( .s (signal_733), .b ({key_s1[121], key_s0[121]}), .a ({signal_3692, signal_1684}), .c ({signal_3943, signal_1932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1236 ( .s (signal_733), .b ({key_s1[122], key_s0[122]}), .a ({signal_3693, signal_1683}), .c ({signal_3945, signal_1931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1237 ( .s (signal_733), .b ({key_s1[123], key_s0[123]}), .a ({signal_3694, signal_1682}), .c ({signal_3947, signal_1930}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1238 ( .s (signal_733), .b ({key_s1[124], key_s0[124]}), .a ({signal_3695, signal_1681}), .c ({signal_3949, signal_1929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1239 ( .s (signal_733), .b ({key_s1[125], key_s0[125]}), .a ({signal_3696, signal_1680}), .c ({signal_3951, signal_1928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1240 ( .s (signal_733), .b ({key_s1[126], key_s0[126]}), .a ({signal_3697, signal_1679}), .c ({signal_3953, signal_1927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1241 ( .s (signal_733), .b ({key_s1[127], key_s0[127]}), .a ({signal_3698, signal_1678}), .c ({signal_3955, signal_1926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1242 ( .s (signal_733), .b ({key_s1[112], key_s0[112]}), .a ({signal_2866, signal_1909}), .c ({signal_2867, signal_1925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1243 ( .s (signal_733), .b ({key_s1[113], key_s0[113]}), .a ({signal_2869, signal_1908}), .c ({signal_2870, signal_1924}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1244 ( .s (signal_733), .b ({key_s1[114], key_s0[114]}), .a ({signal_2872, signal_1907}), .c ({signal_2873, signal_1923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1245 ( .s (signal_733), .b ({key_s1[115], key_s0[115]}), .a ({signal_2875, signal_1906}), .c ({signal_2876, signal_1922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1246 ( .s (signal_733), .b ({key_s1[116], key_s0[116]}), .a ({signal_2878, signal_1905}), .c ({signal_2879, signal_1921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1247 ( .s (signal_733), .b ({key_s1[117], key_s0[117]}), .a ({signal_2881, signal_1904}), .c ({signal_2882, signal_1920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1248 ( .s (signal_733), .b ({key_s1[118], key_s0[118]}), .a ({signal_2884, signal_1903}), .c ({signal_2885, signal_1919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1249 ( .s (signal_733), .b ({key_s1[119], key_s0[119]}), .a ({signal_2887, signal_1902}), .c ({signal_2888, signal_1918}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1250 ( .s (signal_734), .b ({key_s1[104], key_s0[104]}), .a ({signal_2890, signal_1893}), .c ({signal_2891, signal_1917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1251 ( .s (signal_734), .b ({key_s1[105], key_s0[105]}), .a ({signal_2893, signal_1892}), .c ({signal_2894, signal_1916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1252 ( .s (signal_734), .b ({key_s1[106], key_s0[106]}), .a ({signal_2896, signal_1891}), .c ({signal_2897, signal_1915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1253 ( .s (signal_734), .b ({key_s1[107], key_s0[107]}), .a ({signal_2899, signal_1890}), .c ({signal_2900, signal_1914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1254 ( .s (signal_734), .b ({key_s1[108], key_s0[108]}), .a ({signal_2902, signal_1889}), .c ({signal_2903, signal_1913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1255 ( .s (signal_734), .b ({key_s1[109], key_s0[109]}), .a ({signal_2905, signal_1888}), .c ({signal_2906, signal_1912}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1256 ( .s (signal_734), .b ({key_s1[110], key_s0[110]}), .a ({signal_2908, signal_1887}), .c ({signal_2909, signal_1911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1257 ( .s (signal_734), .b ({key_s1[111], key_s0[111]}), .a ({signal_2911, signal_1886}), .c ({signal_2912, signal_1910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1258 ( .s (signal_734), .b ({key_s1[96], key_s0[96]}), .a ({signal_2914, signal_1877}), .c ({signal_2915, signal_1901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1259 ( .s (signal_734), .b ({key_s1[97], key_s0[97]}), .a ({signal_2917, signal_1876}), .c ({signal_2918, signal_1900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1260 ( .s (signal_734), .b ({key_s1[98], key_s0[98]}), .a ({signal_2920, signal_1875}), .c ({signal_2921, signal_1899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1261 ( .s (signal_734), .b ({key_s1[99], key_s0[99]}), .a ({signal_2923, signal_1874}), .c ({signal_2924, signal_1898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1262 ( .s (signal_734), .b ({key_s1[100], key_s0[100]}), .a ({signal_2926, signal_1873}), .c ({signal_2927, signal_1897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1263 ( .s (signal_734), .b ({key_s1[101], key_s0[101]}), .a ({signal_2929, signal_1872}), .c ({signal_2930, signal_1896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1264 ( .s (signal_734), .b ({key_s1[102], key_s0[102]}), .a ({signal_2932, signal_1871}), .c ({signal_2933, signal_1895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1265 ( .s (signal_734), .b ({key_s1[103], key_s0[103]}), .a ({signal_2935, signal_1870}), .c ({signal_2936, signal_1894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1266 ( .s (signal_735), .b ({key_s1[88], key_s0[88]}), .a ({signal_2938, signal_1861}), .c ({signal_2939, signal_1885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1267 ( .s (signal_735), .b ({key_s1[89], key_s0[89]}), .a ({signal_2941, signal_1860}), .c ({signal_2942, signal_1884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1268 ( .s (signal_735), .b ({key_s1[90], key_s0[90]}), .a ({signal_2944, signal_1859}), .c ({signal_2945, signal_1883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1269 ( .s (signal_735), .b ({key_s1[91], key_s0[91]}), .a ({signal_2947, signal_1858}), .c ({signal_2948, signal_1882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1270 ( .s (signal_735), .b ({key_s1[92], key_s0[92]}), .a ({signal_2950, signal_1857}), .c ({signal_2951, signal_1881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1271 ( .s (signal_735), .b ({key_s1[93], key_s0[93]}), .a ({signal_2953, signal_1856}), .c ({signal_2954, signal_1880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1272 ( .s (signal_735), .b ({key_s1[94], key_s0[94]}), .a ({signal_2956, signal_1855}), .c ({signal_2957, signal_1879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1273 ( .s (signal_735), .b ({key_s1[95], key_s0[95]}), .a ({signal_2959, signal_1854}), .c ({signal_2960, signal_1878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1274 ( .s (signal_735), .b ({key_s1[80], key_s0[80]}), .a ({signal_2962, signal_1845}), .c ({signal_2963, signal_1869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1275 ( .s (signal_735), .b ({key_s1[81], key_s0[81]}), .a ({signal_2965, signal_1844}), .c ({signal_2966, signal_1868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1276 ( .s (signal_735), .b ({key_s1[82], key_s0[82]}), .a ({signal_2968, signal_1843}), .c ({signal_2969, signal_1867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1277 ( .s (signal_735), .b ({key_s1[83], key_s0[83]}), .a ({signal_2971, signal_1842}), .c ({signal_2972, signal_1866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1278 ( .s (signal_735), .b ({key_s1[84], key_s0[84]}), .a ({signal_2974, signal_1841}), .c ({signal_2975, signal_1865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1279 ( .s (signal_735), .b ({key_s1[85], key_s0[85]}), .a ({signal_2977, signal_1840}), .c ({signal_2978, signal_1864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1280 ( .s (signal_735), .b ({key_s1[86], key_s0[86]}), .a ({signal_2980, signal_1839}), .c ({signal_2981, signal_1863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1281 ( .s (signal_735), .b ({key_s1[87], key_s0[87]}), .a ({signal_2983, signal_1838}), .c ({signal_2984, signal_1862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1282 ( .s (signal_736), .b ({key_s1[72], key_s0[72]}), .a ({signal_2986, signal_1509}), .c ({signal_2987, signal_1853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1283 ( .s (signal_736), .b ({key_s1[73], key_s0[73]}), .a ({signal_2989, signal_1508}), .c ({signal_2990, signal_1852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1284 ( .s (signal_736), .b ({key_s1[74], key_s0[74]}), .a ({signal_2992, signal_1507}), .c ({signal_2993, signal_1851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1285 ( .s (signal_736), .b ({key_s1[75], key_s0[75]}), .a ({signal_2995, signal_1506}), .c ({signal_2996, signal_1850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1286 ( .s (signal_736), .b ({key_s1[76], key_s0[76]}), .a ({signal_2998, signal_1505}), .c ({signal_2999, signal_1849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1287 ( .s (signal_736), .b ({key_s1[77], key_s0[77]}), .a ({signal_3001, signal_1504}), .c ({signal_3002, signal_1848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1288 ( .s (signal_736), .b ({key_s1[78], key_s0[78]}), .a ({signal_3004, signal_1503}), .c ({signal_3005, signal_1847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1289 ( .s (signal_736), .b ({key_s1[79], key_s0[79]}), .a ({signal_3007, signal_1502}), .c ({signal_3008, signal_1846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1290 ( .s (signal_736), .b ({key_s1[64], key_s0[64]}), .a ({signal_3010, signal_1821}), .c ({signal_3011, signal_1837}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1291 ( .s (signal_736), .b ({key_s1[65], key_s0[65]}), .a ({signal_3013, signal_1820}), .c ({signal_3014, signal_1836}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1292 ( .s (signal_736), .b ({key_s1[66], key_s0[66]}), .a ({signal_3016, signal_1819}), .c ({signal_3017, signal_1835}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1293 ( .s (signal_736), .b ({key_s1[67], key_s0[67]}), .a ({signal_3019, signal_1818}), .c ({signal_3020, signal_1834}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1294 ( .s (signal_736), .b ({key_s1[68], key_s0[68]}), .a ({signal_3022, signal_1817}), .c ({signal_3023, signal_1833}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1295 ( .s (signal_736), .b ({key_s1[69], key_s0[69]}), .a ({signal_3025, signal_1816}), .c ({signal_3026, signal_1832}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1296 ( .s (signal_736), .b ({key_s1[70], key_s0[70]}), .a ({signal_3028, signal_1815}), .c ({signal_3029, signal_1831}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1297 ( .s (signal_736), .b ({key_s1[71], key_s0[71]}), .a ({signal_3031, signal_1814}), .c ({signal_3032, signal_1830}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1298 ( .s (signal_737), .b ({key_s1[56], key_s0[56]}), .a ({signal_3034, signal_1805}), .c ({signal_3035, signal_1829}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1299 ( .s (signal_737), .b ({key_s1[57], key_s0[57]}), .a ({signal_3037, signal_1804}), .c ({signal_3038, signal_1828}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1300 ( .s (signal_737), .b ({key_s1[58], key_s0[58]}), .a ({signal_3040, signal_1803}), .c ({signal_3041, signal_1827}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1301 ( .s (signal_737), .b ({key_s1[59], key_s0[59]}), .a ({signal_3043, signal_1802}), .c ({signal_3044, signal_1826}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1302 ( .s (signal_737), .b ({key_s1[60], key_s0[60]}), .a ({signal_3046, signal_1801}), .c ({signal_3047, signal_1825}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1303 ( .s (signal_737), .b ({key_s1[61], key_s0[61]}), .a ({signal_3049, signal_1800}), .c ({signal_3050, signal_1824}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1304 ( .s (signal_737), .b ({key_s1[62], key_s0[62]}), .a ({signal_3052, signal_1799}), .c ({signal_3053, signal_1823}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1305 ( .s (signal_737), .b ({key_s1[63], key_s0[63]}), .a ({signal_3055, signal_1798}), .c ({signal_3056, signal_1822}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1306 ( .s (signal_737), .b ({key_s1[48], key_s0[48]}), .a ({signal_3058, signal_1789}), .c ({signal_3059, signal_1813}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1307 ( .s (signal_737), .b ({key_s1[49], key_s0[49]}), .a ({signal_3061, signal_1788}), .c ({signal_3062, signal_1812}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1308 ( .s (signal_737), .b ({key_s1[50], key_s0[50]}), .a ({signal_3064, signal_1787}), .c ({signal_3065, signal_1811}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1309 ( .s (signal_737), .b ({key_s1[51], key_s0[51]}), .a ({signal_3067, signal_1786}), .c ({signal_3068, signal_1810}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1310 ( .s (signal_737), .b ({key_s1[52], key_s0[52]}), .a ({signal_3070, signal_1785}), .c ({signal_3071, signal_1809}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1311 ( .s (signal_737), .b ({key_s1[53], key_s0[53]}), .a ({signal_3073, signal_1784}), .c ({signal_3074, signal_1808}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1312 ( .s (signal_737), .b ({key_s1[54], key_s0[54]}), .a ({signal_3076, signal_1783}), .c ({signal_3077, signal_1807}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1313 ( .s (signal_737), .b ({key_s1[55], key_s0[55]}), .a ({signal_3079, signal_1782}), .c ({signal_3080, signal_1806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1314 ( .s (signal_738), .b ({key_s1[40], key_s0[40]}), .a ({signal_3082, signal_1773}), .c ({signal_3083, signal_1797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1315 ( .s (signal_738), .b ({key_s1[41], key_s0[41]}), .a ({signal_3085, signal_1772}), .c ({signal_3086, signal_1796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1316 ( .s (signal_738), .b ({key_s1[42], key_s0[42]}), .a ({signal_3088, signal_1771}), .c ({signal_3089, signal_1795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1317 ( .s (signal_738), .b ({key_s1[43], key_s0[43]}), .a ({signal_3091, signal_1770}), .c ({signal_3092, signal_1794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1318 ( .s (signal_738), .b ({key_s1[44], key_s0[44]}), .a ({signal_3094, signal_1769}), .c ({signal_3095, signal_1793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1319 ( .s (signal_738), .b ({key_s1[45], key_s0[45]}), .a ({signal_3097, signal_1768}), .c ({signal_3098, signal_1792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1320 ( .s (signal_738), .b ({key_s1[46], key_s0[46]}), .a ({signal_3100, signal_1767}), .c ({signal_3101, signal_1791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1321 ( .s (signal_738), .b ({key_s1[47], key_s0[47]}), .a ({signal_3103, signal_1766}), .c ({signal_3104, signal_1790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1322 ( .s (signal_738), .b ({key_s1[32], key_s0[32]}), .a ({signal_3106, signal_1749}), .c ({signal_3107, signal_1781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1323 ( .s (signal_738), .b ({key_s1[33], key_s0[33]}), .a ({signal_3109, signal_1748}), .c ({signal_3110, signal_1780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1324 ( .s (signal_738), .b ({key_s1[34], key_s0[34]}), .a ({signal_3112, signal_1747}), .c ({signal_3113, signal_1779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1325 ( .s (signal_738), .b ({key_s1[35], key_s0[35]}), .a ({signal_3115, signal_1746}), .c ({signal_3116, signal_1778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1326 ( .s (signal_738), .b ({key_s1[36], key_s0[36]}), .a ({signal_3118, signal_1745}), .c ({signal_3119, signal_1777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1327 ( .s (signal_738), .b ({key_s1[37], key_s0[37]}), .a ({signal_3121, signal_1744}), .c ({signal_3122, signal_1776}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1328 ( .s (signal_738), .b ({key_s1[38], key_s0[38]}), .a ({signal_3124, signal_1743}), .c ({signal_3125, signal_1775}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1329 ( .s (signal_738), .b ({key_s1[39], key_s0[39]}), .a ({signal_3127, signal_1742}), .c ({signal_3128, signal_1774}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1330 ( .s (signal_739), .b ({key_s1[24], key_s0[24]}), .a ({signal_3130, signal_1733}), .c ({signal_3131, signal_1765}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1331 ( .s (signal_739), .b ({key_s1[25], key_s0[25]}), .a ({signal_3133, signal_1732}), .c ({signal_3134, signal_1764}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1332 ( .s (signal_739), .b ({key_s1[26], key_s0[26]}), .a ({signal_3136, signal_1731}), .c ({signal_3137, signal_1763}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1333 ( .s (signal_739), .b ({key_s1[27], key_s0[27]}), .a ({signal_3139, signal_1730}), .c ({signal_3140, signal_1762}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1334 ( .s (signal_739), .b ({key_s1[28], key_s0[28]}), .a ({signal_3142, signal_1729}), .c ({signal_3143, signal_1761}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1335 ( .s (signal_739), .b ({key_s1[29], key_s0[29]}), .a ({signal_3145, signal_1728}), .c ({signal_3146, signal_1760}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1336 ( .s (signal_739), .b ({key_s1[30], key_s0[30]}), .a ({signal_3148, signal_1727}), .c ({signal_3149, signal_1759}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1337 ( .s (signal_739), .b ({key_s1[31], key_s0[31]}), .a ({signal_3151, signal_1726}), .c ({signal_3152, signal_1758}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1338 ( .s (signal_739), .b ({key_s1[16], key_s0[16]}), .a ({signal_3154, signal_1717}), .c ({signal_3155, signal_1741}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1339 ( .s (signal_739), .b ({key_s1[17], key_s0[17]}), .a ({signal_3157, signal_1716}), .c ({signal_3158, signal_1740}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1340 ( .s (signal_739), .b ({key_s1[18], key_s0[18]}), .a ({signal_3160, signal_1715}), .c ({signal_3161, signal_1739}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1341 ( .s (signal_739), .b ({key_s1[19], key_s0[19]}), .a ({signal_3163, signal_1714}), .c ({signal_3164, signal_1738}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1342 ( .s (signal_739), .b ({key_s1[20], key_s0[20]}), .a ({signal_3166, signal_1713}), .c ({signal_3167, signal_1737}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1343 ( .s (signal_739), .b ({key_s1[21], key_s0[21]}), .a ({signal_3169, signal_1712}), .c ({signal_3170, signal_1736}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1344 ( .s (signal_739), .b ({key_s1[22], key_s0[22]}), .a ({signal_3172, signal_1711}), .c ({signal_3173, signal_1735}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1345 ( .s (signal_739), .b ({key_s1[23], key_s0[23]}), .a ({signal_3175, signal_1710}), .c ({signal_3176, signal_1734}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1346 ( .s (signal_740), .b ({key_s1[8], key_s0[8]}), .a ({signal_3178, signal_1701}), .c ({signal_3179, signal_1725}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1347 ( .s (signal_740), .b ({key_s1[9], key_s0[9]}), .a ({signal_3181, signal_1700}), .c ({signal_3182, signal_1724}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1348 ( .s (signal_740), .b ({key_s1[10], key_s0[10]}), .a ({signal_3184, signal_1699}), .c ({signal_3185, signal_1723}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1349 ( .s (signal_740), .b ({key_s1[11], key_s0[11]}), .a ({signal_3187, signal_1698}), .c ({signal_3188, signal_1722}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1350 ( .s (signal_740), .b ({key_s1[12], key_s0[12]}), .a ({signal_3190, signal_1697}), .c ({signal_3191, signal_1721}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1351 ( .s (signal_740), .b ({key_s1[13], key_s0[13]}), .a ({signal_3193, signal_1696}), .c ({signal_3194, signal_1720}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1352 ( .s (signal_740), .b ({key_s1[14], key_s0[14]}), .a ({signal_3196, signal_1695}), .c ({signal_3197, signal_1719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1353 ( .s (signal_740), .b ({key_s1[15], key_s0[15]}), .a ({signal_3199, signal_1694}), .c ({signal_3200, signal_1718}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1354 ( .s (signal_740), .b ({key_s1[0], key_s0[0]}), .a ({signal_2406, signal_1493}), .c ({signal_3202, signal_1709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1355 ( .s (signal_740), .b ({key_s1[1], key_s0[1]}), .a ({signal_2409, signal_1492}), .c ({signal_3204, signal_1708}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1356 ( .s (signal_740), .b ({key_s1[2], key_s0[2]}), .a ({signal_2412, signal_1491}), .c ({signal_3206, signal_1707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1357 ( .s (signal_740), .b ({key_s1[3], key_s0[3]}), .a ({signal_2415, signal_1490}), .c ({signal_3208, signal_1706}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1358 ( .s (signal_740), .b ({key_s1[4], key_s0[4]}), .a ({signal_2418, signal_1489}), .c ({signal_3210, signal_1705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1359 ( .s (signal_740), .b ({key_s1[5], key_s0[5]}), .a ({signal_2421, signal_1488}), .c ({signal_3212, signal_1704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1360 ( .s (signal_740), .b ({key_s1[6], key_s0[6]}), .a ({signal_2424, signal_1487}), .c ({signal_3214, signal_1703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1361 ( .s (signal_740), .b ({key_s1[7], key_s0[7]}), .a ({signal_2427, signal_1486}), .c ({signal_3216, signal_1702}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1362 ( .a ({signal_2545, signal_1150}), .b ({signal_2447, signal_1151}), .c ({signal_3217, signal_1454}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1363 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2447, signal_1151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1364 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2474, signal_1934}), .c ({signal_2545, signal_1150}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1365 ( .a ({signal_2546, signal_1152}), .b ({signal_2450, signal_1153}), .c ({signal_3218, signal_1455}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1366 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2450, signal_1153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1367 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2476, signal_1935}), .c ({signal_2546, signal_1152}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1368 ( .a ({signal_2547, signal_1154}), .b ({signal_2453, signal_1155}), .c ({signal_3219, signal_1456}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1369 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2453, signal_1155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1370 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2478, signal_1936}), .c ({signal_2547, signal_1154}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1371 ( .a ({signal_3220, signal_1156}), .b ({signal_2456, signal_1157}), .c ({signal_3261, signal_1457}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1372 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2456, signal_1157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1373 ( .a ({signal_2469, signal_1942}), .b ({signal_2550, signal_1937}), .c ({signal_3220, signal_1156}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1374 ( .a ({signal_3221, signal_1158}), .b ({signal_2459, signal_1159}), .c ({signal_3262, signal_1458}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1375 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2459, signal_1159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1376 ( .a ({signal_2470, signal_1943}), .b ({signal_2551, signal_1938}), .c ({signal_3221, signal_1158}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1377 ( .a ({signal_2548, signal_1160}), .b ({signal_2462, signal_1161}), .c ({signal_3222, signal_1459}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1378 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2462, signal_1161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1379 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2481, signal_1939}), .c ({signal_2548, signal_1160}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1380 ( .a ({signal_3223, signal_1162}), .b ({signal_2465, signal_1163}), .c ({signal_3263, signal_1460}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1381 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2465, signal_1163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1382 ( .a ({signal_2471, signal_1945}), .b ({signal_2552, signal_1940}), .c ({signal_3223, signal_1162}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1383 ( .a ({signal_2549, signal_1164}), .b ({signal_2468, signal_1165}), .c ({signal_3224, signal_1461}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1384 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2468, signal_1165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1385 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2483, signal_1941}), .c ({signal_2549, signal_1164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1386 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2469, signal_1942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1387 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2470, signal_1943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1388 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2471, signal_1945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1389 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2474, signal_1934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1390 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2476, signal_1935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1391 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2478, signal_1936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1392 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2485, signal_1946}), .c ({signal_2550, signal_1937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1393 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_2486, signal_1947}), .c ({signal_2551, signal_1938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1394 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2481, signal_1939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1395 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2487, signal_1949}), .c ({signal_2552, signal_1940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1396 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2483, signal_1941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1397 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2485, signal_1946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1398 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2486, signal_1947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1399 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2487, signal_1949}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1400 ( .a ({signal_2553, signal_1166}), .b ({signal_2488, signal_1167}), .c ({signal_3225, signal_1462}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1401 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2488, signal_1167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1402 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_2499, signal_1950}), .c ({signal_2553, signal_1166}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1403 ( .a ({signal_2554, signal_1168}), .b ({signal_2489, signal_1169}), .c ({signal_3226, signal_1463}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1404 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2489, signal_1169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1405 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_2500, signal_1951}), .c ({signal_2554, signal_1168}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1406 ( .a ({signal_2555, signal_1170}), .b ({signal_2490, signal_1171}), .c ({signal_3227, signal_1464}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1407 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2490, signal_1171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1408 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2501, signal_1952}), .c ({signal_2555, signal_1170}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1409 ( .a ({signal_3228, signal_1172}), .b ({signal_2491, signal_1173}), .c ({signal_3264, signal_1465}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1410 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2491, signal_1173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1411 ( .a ({signal_2496, signal_1184}), .b ({signal_2558, signal_1953}), .c ({signal_3228, signal_1172}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1412 ( .a ({signal_3229, signal_1174}), .b ({signal_2492, signal_1175}), .c ({signal_3265, signal_1466}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1413 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2492, signal_1175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1414 ( .a ({signal_2497, signal_1183}), .b ({signal_2559, signal_1954}), .c ({signal_3229, signal_1174}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1415 ( .a ({signal_2556, signal_1176}), .b ({signal_2493, signal_1177}), .c ({signal_3230, signal_1467}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1416 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2493, signal_1177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1417 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2502, signal_1955}), .c ({signal_2556, signal_1176}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1418 ( .a ({signal_3231, signal_1178}), .b ({signal_2494, signal_1179}), .c ({signal_3266, signal_1468}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1419 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2494, signal_1179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1420 ( .a ({signal_2498, signal_1182}), .b ({signal_2560, signal_1956}), .c ({signal_3231, signal_1178}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1421 ( .a ({signal_2557, signal_1180}), .b ({signal_2495, signal_1181}), .c ({signal_3232, signal_1469}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1422 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2495, signal_1181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1423 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_2503, signal_1957}), .c ({signal_2557, signal_1180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1424 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2496, signal_1184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1425 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2497, signal_1183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1426 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2498, signal_1182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1427 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2499, signal_1950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1428 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2500, signal_1951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1429 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2501, signal_1952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1430 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2504, signal_1958}), .c ({signal_2558, signal_1953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1431 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_2505, signal_1959}), .c ({signal_2559, signal_1954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1432 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_2502, signal_1955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1433 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2506, signal_1961}), .c ({signal_2560, signal_1956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1434 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2503, signal_1957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1435 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2504, signal_1958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1436 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2505, signal_1959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1437 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2506, signal_1961}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1438 ( .a ({signal_2561, signal_1185}), .b ({signal_2507, signal_1186}), .c ({signal_3233, signal_1470}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1439 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_2507, signal_1186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1440 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_2518, signal_1962}), .c ({signal_2561, signal_1185}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1441 ( .a ({signal_2562, signal_1187}), .b ({signal_2508, signal_1188}), .c ({signal_3234, signal_1471}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1442 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_2508, signal_1188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1443 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2519, signal_1963}), .c ({signal_2562, signal_1187}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1444 ( .a ({signal_2563, signal_1189}), .b ({signal_2509, signal_1190}), .c ({signal_3235, signal_1472}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1445 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_2509, signal_1190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1446 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2520, signal_1964}), .c ({signal_2563, signal_1189}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1447 ( .a ({signal_3236, signal_1191}), .b ({signal_2510, signal_1192}), .c ({signal_3267, signal_1473}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1448 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_2510, signal_1192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1449 ( .a ({signal_2515, signal_1203}), .b ({signal_2566, signal_1965}), .c ({signal_3236, signal_1191}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1450 ( .a ({signal_3237, signal_1193}), .b ({signal_2511, signal_1194}), .c ({signal_3268, signal_1474}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1451 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_2511, signal_1194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1452 ( .a ({signal_2516, signal_1202}), .b ({signal_2567, signal_1966}), .c ({signal_3237, signal_1193}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1453 ( .a ({signal_2564, signal_1195}), .b ({signal_2512, signal_1196}), .c ({signal_3238, signal_1475}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1454 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .c ({signal_2512, signal_1196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1455 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2521, signal_1967}), .c ({signal_2564, signal_1195}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1456 ( .a ({signal_3239, signal_1197}), .b ({signal_2513, signal_1198}), .c ({signal_3269, signal_1476}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1457 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2513, signal_1198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1458 ( .a ({signal_2517, signal_1201}), .b ({signal_2568, signal_1968}), .c ({signal_3239, signal_1197}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1459 ( .a ({signal_2565, signal_1199}), .b ({signal_2514, signal_1200}), .c ({signal_3240, signal_1477}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1460 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2514, signal_1200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1461 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_2522, signal_1969}), .c ({signal_2565, signal_1199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1462 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2515, signal_1203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1463 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2516, signal_1202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1464 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .c ({signal_2517, signal_1201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1465 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_2518, signal_1962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1466 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_2519, signal_1963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1467 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_2520, signal_1964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1468 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2523, signal_1970}), .c ({signal_2566, signal_1965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1469 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_2524, signal_1971}), .c ({signal_2567, signal_1966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1470 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_2521, signal_1967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1471 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2525, signal_1973}), .c ({signal_2568, signal_1968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1472 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_2522, signal_1969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1473 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2523, signal_1970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1474 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2524, signal_1971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1475 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2525, signal_1973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1476 ( .a ({signal_2569, signal_1204}), .b ({signal_2526, signal_1205}), .c ({signal_3241, signal_1478}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1477 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_2526, signal_1205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1478 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_2537, signal_1974}), .c ({signal_2569, signal_1204}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1479 ( .a ({signal_2570, signal_1206}), .b ({signal_2527, signal_1207}), .c ({signal_3242, signal_1479}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1480 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_2527, signal_1207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1481 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2538, signal_1975}), .c ({signal_2570, signal_1206}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1482 ( .a ({signal_2571, signal_1208}), .b ({signal_2528, signal_1209}), .c ({signal_3243, signal_1480}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1483 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_2528, signal_1209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1484 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2539, signal_1976}), .c ({signal_2571, signal_1208}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1485 ( .a ({signal_3244, signal_1210}), .b ({signal_2529, signal_1211}), .c ({signal_3270, signal_1481}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1486 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_2529, signal_1211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1487 ( .a ({signal_2534, signal_1222}), .b ({signal_2574, signal_1977}), .c ({signal_3244, signal_1210}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1488 ( .a ({signal_3245, signal_1212}), .b ({signal_2530, signal_1213}), .c ({signal_3271, signal_1482}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1489 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_2530, signal_1213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1490 ( .a ({signal_2535, signal_1221}), .b ({signal_2575, signal_1978}), .c ({signal_3245, signal_1212}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1491 ( .a ({signal_2572, signal_1214}), .b ({signal_2531, signal_1215}), .c ({signal_3246, signal_1483}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1492 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .c ({signal_2531, signal_1215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1493 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2540, signal_1979}), .c ({signal_2572, signal_1214}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1494 ( .a ({signal_3247, signal_1216}), .b ({signal_2532, signal_1217}), .c ({signal_3272, signal_1484}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1495 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_2532, signal_1217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1496 ( .a ({signal_2536, signal_1220}), .b ({signal_2576, signal_1980}), .c ({signal_3247, signal_1216}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1497 ( .a ({signal_2573, signal_1218}), .b ({signal_2533, signal_1219}), .c ({signal_3248, signal_1485}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_1498 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .c ({signal_2533, signal_1219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1499 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_2541, signal_1981}), .c ({signal_2573, signal_1218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1500 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_2534, signal_1222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1501 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .c ({signal_2535, signal_1221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1502 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .c ({signal_2536, signal_1220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1503 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_2537, signal_1974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1504 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_2538, signal_1975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1505 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_2539, signal_1976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1506 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2542, signal_1225}), .c ({signal_2574, signal_1977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1507 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2543, signal_1224}), .c ({signal_2575, signal_1978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1508 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_2540, signal_1979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1509 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2544, signal_1223}), .c ({signal_2576, signal_1980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1510 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_2541, signal_1981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1511 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_2542, signal_1225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1512 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .c ({signal_2543, signal_1224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_1513 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .c ({signal_2544, signal_1223}) ) ;
    NOR2_X1 cell_1514 ( .A1 (signal_1255), .A2 (signal_1226), .ZN (signal_1494) ) ;
    NOR2_X1 cell_1515 ( .A1 (signal_1257), .A2 (signal_1226), .ZN (signal_1495) ) ;
    AND2_X1 cell_1516 ( .A1 (signal_1273), .A2 (signal_397), .ZN (signal_1496) ) ;
    AND2_X1 cell_1517 ( .A1 (signal_1272), .A2 (signal_397), .ZN (signal_1497) ) ;
    NOR2_X1 cell_1518 ( .A1 (signal_1261), .A2 (signal_1226), .ZN (signal_1498) ) ;
    NOR2_X1 cell_1519 ( .A1 (signal_1263), .A2 (signal_1226), .ZN (signal_1499) ) ;
    NOR2_X1 cell_1520 ( .A1 (signal_1265), .A2 (signal_1226), .ZN (signal_1500) ) ;
    NOR2_X1 cell_1521 ( .A1 (signal_1267), .A2 (signal_1226), .ZN (signal_1501) ) ;
    INV_X1 cell_1522 ( .A (signal_397), .ZN (signal_1226) ) ;
    NAND2_X1 cell_1523 ( .A1 (signal_1227), .A2 (signal_1228), .ZN (signal_401) ) ;
    NOR2_X1 cell_1524 ( .A1 (signal_1229), .A2 (signal_1230), .ZN (signal_1228) ) ;
    NAND2_X1 cell_1525 ( .A1 (signal_1231), .A2 (signal_1232), .ZN (signal_1230) ) ;
    NOR2_X1 cell_1526 ( .A1 (signal_1269), .A2 (signal_1261), .ZN (signal_1232) ) ;
    NOR2_X1 cell_1527 ( .A1 (signal_1274), .A2 (signal_1267), .ZN (signal_1231) ) ;
    NAND2_X1 cell_1528 ( .A1 (signal_1270), .A2 (signal_1254), .ZN (signal_1229) ) ;
    NOR2_X1 cell_1529 ( .A1 (signal_1272), .A2 (signal_1273), .ZN (signal_1227) ) ;
    NAND2_X1 cell_1530 ( .A1 (signal_393), .A2 (signal_1233), .ZN (signal_1275) ) ;
    MUX2_X1 cell_1531 ( .S (signal_1253), .A (signal_1255), .B (signal_1267), .Z (signal_1233) ) ;
    NAND2_X1 cell_1532 ( .A1 (signal_1234), .A2 (signal_1235), .ZN (signal_1266) ) ;
    NAND2_X1 cell_1533 ( .A1 (signal_1236), .A2 (signal_1269), .ZN (signal_1235) ) ;
    NAND2_X1 cell_1534 ( .A1 (signal_1237), .A2 (signal_1238), .ZN (signal_1234) ) ;
    XOR2_X1 cell_1535 ( .A (signal_1268), .B (signal_1254), .Z (signal_1237) ) ;
    NAND2_X1 cell_1536 ( .A1 (signal_393), .A2 (signal_1239), .ZN (signal_1264) ) ;
    MUX2_X1 cell_1537 ( .S (signal_1253), .A (signal_1265), .B (signal_1263), .Z (signal_1239) ) ;
    NAND2_X1 cell_1538 ( .A1 (signal_393), .A2 (signal_1240), .ZN (signal_1262) ) ;
    MUX2_X1 cell_1539 ( .S (signal_1253), .A (signal_1241), .B (signal_1261), .Z (signal_1240) ) ;
    XNOR2_X1 cell_1540 ( .A (signal_1254), .B (signal_1270), .ZN (signal_1241) ) ;
    NAND2_X1 cell_1541 ( .A1 (signal_1242), .A2 (signal_1243), .ZN (signal_1260) ) ;
    NAND2_X1 cell_1542 ( .A1 (signal_1272), .A2 (signal_1236), .ZN (signal_1243) ) ;
    NAND2_X1 cell_1543 ( .A1 (signal_1244), .A2 (signal_1238), .ZN (signal_1242) ) ;
    XOR2_X1 cell_1544 ( .A (signal_1261), .B (signal_1255), .Z (signal_1244) ) ;
    NAND2_X1 cell_1545 ( .A1 (signal_1245), .A2 (signal_1246), .ZN (signal_1259) ) ;
    NAND2_X1 cell_1546 ( .A1 (signal_1272), .A2 (signal_1238), .ZN (signal_1246) ) ;
    NAND2_X1 cell_1547 ( .A1 (signal_1273), .A2 (signal_1236), .ZN (signal_1245) ) ;
    NAND2_X1 cell_1548 ( .A1 (signal_1247), .A2 (signal_1248), .ZN (signal_1258) ) ;
    NAND2_X1 cell_1549 ( .A1 (signal_1273), .A2 (signal_1238), .ZN (signal_1248) ) ;
    NOR2_X1 cell_1550 ( .A1 (signal_1253), .A2 (signal_1252), .ZN (signal_1238) ) ;
    NAND2_X1 cell_1551 ( .A1 (signal_1274), .A2 (signal_1236), .ZN (signal_1247) ) ;
    NOR2_X1 cell_1552 ( .A1 (signal_395), .A2 (signal_1252), .ZN (signal_1236) ) ;
    NAND2_X1 cell_1553 ( .A1 (signal_393), .A2 (signal_1249), .ZN (signal_1256) ) ;
    MUX2_X1 cell_1554 ( .S (signal_1253), .A (signal_1257), .B (signal_1255), .Z (signal_1249) ) ;
    NAND2_X1 cell_1555 ( .A1 (signal_1272), .A2 (signal_1270), .ZN (signal_1251) ) ;
    NAND2_X1 cell_1556 ( .A1 (signal_1269), .A2 (signal_1273), .ZN (signal_1250) ) ;
    INV_X1 cell_1557 ( .A (signal_393), .ZN (signal_1252) ) ;
    INV_X1 cell_1558 ( .A (signal_395), .ZN (signal_1253) ) ;
    NOR2_X1 cell_1559 ( .A1 (signal_1250), .A2 (signal_1251), .ZN (signal_399) ) ;
    INV_X1 cell_1560 ( .A (signal_1268), .ZN (signal_1267) ) ;
    INV_X1 cell_1562 ( .A (signal_1269), .ZN (signal_1265) ) ;
    INV_X1 cell_1564 ( .A (signal_1270), .ZN (signal_1263) ) ;
    INV_X1 cell_1566 ( .A (signal_1271), .ZN (signal_1261) ) ;
    INV_X1 cell_1572 ( .A (signal_1274), .ZN (signal_1257) ) ;
    INV_X1 cell_1574 ( .A (signal_1254), .ZN (signal_1255) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1576 ( .s (signal_394), .b ({signal_2407, signal_1413}), .a ({signal_2986, signal_1509}), .c ({signal_3249, signal_1517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1577 ( .s (signal_394), .b ({signal_2410, signal_1412}), .a ({signal_2989, signal_1508}), .c ({signal_3250, signal_1516}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1578 ( .s (signal_394), .b ({signal_2413, signal_1411}), .a ({signal_2992, signal_1507}), .c ({signal_3251, signal_1515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1579 ( .s (signal_394), .b ({signal_2416, signal_1410}), .a ({signal_2995, signal_1506}), .c ({signal_3252, signal_1514}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1580 ( .s (signal_394), .b ({signal_2419, signal_1409}), .a ({signal_2998, signal_1505}), .c ({signal_3253, signal_1513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1581 ( .s (signal_394), .b ({signal_2422, signal_1408}), .a ({signal_3001, signal_1504}), .c ({signal_3254, signal_1512}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1582 ( .s (signal_394), .b ({signal_2425, signal_1407}), .a ({signal_3004, signal_1503}), .c ({signal_3255, signal_1511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1583 ( .s (signal_394), .b ({signal_2428, signal_1406}), .a ({signal_3007, signal_1502}), .c ({signal_3256, signal_1510}) ) ;
    INV_X1 cell_1712 ( .A (signal_393), .ZN (signal_402) ) ;

    /* cells in depth 1 */
    buf_clk cell_2145 ( .C (clk), .D (signal_1511), .Q (signal_4691) ) ;
    buf_clk cell_2147 ( .C (clk), .D (signal_3255), .Q (signal_4693) ) ;
    buf_clk cell_2149 ( .C (clk), .D (signal_1512), .Q (signal_4695) ) ;
    buf_clk cell_2151 ( .C (clk), .D (signal_3254), .Q (signal_4697) ) ;
    buf_clk cell_2169 ( .C (clk), .D (signal_1513), .Q (signal_4715) ) ;
    buf_clk cell_2173 ( .C (clk), .D (signal_3253), .Q (signal_4719) ) ;
    buf_clk cell_2297 ( .C (clk), .D (signal_1514), .Q (signal_4843) ) ;
    buf_clk cell_2305 ( .C (clk), .D (signal_3252), .Q (signal_4851) ) ;
    buf_clk cell_2341 ( .C (clk), .D (signal_1515), .Q (signal_4887) ) ;
    buf_clk cell_2351 ( .C (clk), .D (signal_3251), .Q (signal_4897) ) ;
    buf_clk cell_2361 ( .C (clk), .D (signal_1516), .Q (signal_4907) ) ;
    buf_clk cell_2373 ( .C (clk), .D (signal_3250), .Q (signal_4919) ) ;
    buf_clk cell_2385 ( .C (clk), .D (signal_399), .Q (signal_4931) ) ;
    buf_clk cell_2401 ( .C (clk), .D (signal_1413), .Q (signal_4947) ) ;
    buf_clk cell_2417 ( .C (clk), .D (signal_2407), .Q (signal_4963) ) ;
    buf_clk cell_2433 ( .C (clk), .D (signal_1412), .Q (signal_4979) ) ;
    buf_clk cell_2449 ( .C (clk), .D (signal_2410), .Q (signal_4995) ) ;
    buf_clk cell_2465 ( .C (clk), .D (signal_1411), .Q (signal_5011) ) ;
    buf_clk cell_2481 ( .C (clk), .D (signal_2413), .Q (signal_5027) ) ;
    buf_clk cell_2497 ( .C (clk), .D (signal_1410), .Q (signal_5043) ) ;
    buf_clk cell_2513 ( .C (clk), .D (signal_2416), .Q (signal_5059) ) ;
    buf_clk cell_2529 ( .C (clk), .D (signal_1409), .Q (signal_5075) ) ;
    buf_clk cell_2545 ( .C (clk), .D (signal_2419), .Q (signal_5091) ) ;
    buf_clk cell_2561 ( .C (clk), .D (signal_1408), .Q (signal_5107) ) ;
    buf_clk cell_2577 ( .C (clk), .D (signal_2422), .Q (signal_5123) ) ;
    buf_clk cell_2593 ( .C (clk), .D (signal_1407), .Q (signal_5139) ) ;
    buf_clk cell_2609 ( .C (clk), .D (signal_2425), .Q (signal_5155) ) ;
    buf_clk cell_2625 ( .C (clk), .D (signal_1406), .Q (signal_5171) ) ;
    buf_clk cell_2641 ( .C (clk), .D (signal_2428), .Q (signal_5187) ) ;
    buf_clk cell_2657 ( .C (clk), .D (signal_464), .Q (signal_5203) ) ;
    buf_clk cell_2673 ( .C (clk), .D (ciphertext_s0[8]), .Q (signal_5219) ) ;
    buf_clk cell_2689 ( .C (clk), .D (ciphertext_s1[8]), .Q (signal_5235) ) ;
    buf_clk cell_2705 ( .C (clk), .D (ciphertext_s0[9]), .Q (signal_5251) ) ;
    buf_clk cell_2721 ( .C (clk), .D (ciphertext_s1[9]), .Q (signal_5267) ) ;
    buf_clk cell_2737 ( .C (clk), .D (ciphertext_s0[10]), .Q (signal_5283) ) ;
    buf_clk cell_2753 ( .C (clk), .D (ciphertext_s1[10]), .Q (signal_5299) ) ;
    buf_clk cell_2769 ( .C (clk), .D (ciphertext_s0[11]), .Q (signal_5315) ) ;
    buf_clk cell_2785 ( .C (clk), .D (ciphertext_s1[11]), .Q (signal_5331) ) ;
    buf_clk cell_2801 ( .C (clk), .D (ciphertext_s0[12]), .Q (signal_5347) ) ;
    buf_clk cell_2817 ( .C (clk), .D (ciphertext_s1[12]), .Q (signal_5363) ) ;
    buf_clk cell_2833 ( .C (clk), .D (ciphertext_s0[13]), .Q (signal_5379) ) ;
    buf_clk cell_2849 ( .C (clk), .D (ciphertext_s1[13]), .Q (signal_5395) ) ;
    buf_clk cell_2865 ( .C (clk), .D (ciphertext_s0[14]), .Q (signal_5411) ) ;
    buf_clk cell_2881 ( .C (clk), .D (ciphertext_s1[14]), .Q (signal_5427) ) ;
    buf_clk cell_2897 ( .C (clk), .D (ciphertext_s0[15]), .Q (signal_5443) ) ;
    buf_clk cell_2913 ( .C (clk), .D (ciphertext_s1[15]), .Q (signal_5459) ) ;
    buf_clk cell_2929 ( .C (clk), .D (signal_455), .Q (signal_5475) ) ;
    buf_clk cell_2945 ( .C (clk), .D (signal_1453), .Q (signal_5491) ) ;
    buf_clk cell_2961 ( .C (clk), .D (signal_3278), .Q (signal_5507) ) ;
    buf_clk cell_2977 ( .C (clk), .D (signal_1452), .Q (signal_5523) ) ;
    buf_clk cell_2993 ( .C (clk), .D (signal_3279), .Q (signal_5539) ) ;
    buf_clk cell_3009 ( .C (clk), .D (signal_1451), .Q (signal_5555) ) ;
    buf_clk cell_3025 ( .C (clk), .D (signal_3257), .Q (signal_5571) ) ;
    buf_clk cell_3041 ( .C (clk), .D (signal_1450), .Q (signal_5587) ) ;
    buf_clk cell_3057 ( .C (clk), .D (signal_3280), .Q (signal_5603) ) ;
    buf_clk cell_3073 ( .C (clk), .D (signal_1449), .Q (signal_5619) ) ;
    buf_clk cell_3089 ( .C (clk), .D (signal_3281), .Q (signal_5635) ) ;
    buf_clk cell_3105 ( .C (clk), .D (signal_1448), .Q (signal_5651) ) ;
    buf_clk cell_3121 ( .C (clk), .D (signal_3258), .Q (signal_5667) ) ;
    buf_clk cell_3137 ( .C (clk), .D (signal_1447), .Q (signal_5683) ) ;
    buf_clk cell_3153 ( .C (clk), .D (signal_3259), .Q (signal_5699) ) ;
    buf_clk cell_3169 ( .C (clk), .D (signal_1446), .Q (signal_5715) ) ;
    buf_clk cell_3185 ( .C (clk), .D (signal_3260), .Q (signal_5731) ) ;
    buf_clk cell_3201 ( .C (clk), .D (signal_452), .Q (signal_5747) ) ;
    buf_clk cell_3217 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_5763) ) ;
    buf_clk cell_3233 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_5779) ) ;
    buf_clk cell_3249 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_5795) ) ;
    buf_clk cell_3265 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_5811) ) ;
    buf_clk cell_3281 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_5827) ) ;
    buf_clk cell_3297 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_5843) ) ;
    buf_clk cell_3313 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_5859) ) ;
    buf_clk cell_3329 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_5875) ) ;
    buf_clk cell_3345 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_5891) ) ;
    buf_clk cell_3361 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_5907) ) ;
    buf_clk cell_3377 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_5923) ) ;
    buf_clk cell_3393 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_5939) ) ;
    buf_clk cell_3409 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_5955) ) ;
    buf_clk cell_3425 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_5971) ) ;
    buf_clk cell_3441 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_5987) ) ;
    buf_clk cell_3457 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_6003) ) ;
    buf_clk cell_3473 ( .C (clk), .D (signal_1486), .Q (signal_6019) ) ;
    buf_clk cell_3489 ( .C (clk), .D (signal_2427), .Q (signal_6035) ) ;
    buf_clk cell_3505 ( .C (clk), .D (signal_1494), .Q (signal_6051) ) ;
    buf_clk cell_3521 ( .C (clk), .D (signal_1487), .Q (signal_6067) ) ;
    buf_clk cell_3537 ( .C (clk), .D (signal_2424), .Q (signal_6083) ) ;
    buf_clk cell_3553 ( .C (clk), .D (signal_1495), .Q (signal_6099) ) ;
    buf_clk cell_3569 ( .C (clk), .D (signal_1488), .Q (signal_6115) ) ;
    buf_clk cell_3585 ( .C (clk), .D (signal_2421), .Q (signal_6131) ) ;
    buf_clk cell_3601 ( .C (clk), .D (signal_1496), .Q (signal_6147) ) ;
    buf_clk cell_3617 ( .C (clk), .D (signal_1489), .Q (signal_6163) ) ;
    buf_clk cell_3633 ( .C (clk), .D (signal_2418), .Q (signal_6179) ) ;
    buf_clk cell_3649 ( .C (clk), .D (signal_1497), .Q (signal_6195) ) ;
    buf_clk cell_3665 ( .C (clk), .D (signal_1490), .Q (signal_6211) ) ;
    buf_clk cell_3681 ( .C (clk), .D (signal_2415), .Q (signal_6227) ) ;
    buf_clk cell_3697 ( .C (clk), .D (signal_1498), .Q (signal_6243) ) ;
    buf_clk cell_3713 ( .C (clk), .D (signal_1491), .Q (signal_6259) ) ;
    buf_clk cell_3729 ( .C (clk), .D (signal_2412), .Q (signal_6275) ) ;
    buf_clk cell_3745 ( .C (clk), .D (signal_1499), .Q (signal_6291) ) ;
    buf_clk cell_3761 ( .C (clk), .D (signal_1492), .Q (signal_6307) ) ;
    buf_clk cell_3777 ( .C (clk), .D (signal_2409), .Q (signal_6323) ) ;
    buf_clk cell_3793 ( .C (clk), .D (signal_1500), .Q (signal_6339) ) ;
    buf_clk cell_3809 ( .C (clk), .D (signal_1493), .Q (signal_6355) ) ;
    buf_clk cell_3825 ( .C (clk), .D (signal_2406), .Q (signal_6371) ) ;
    buf_clk cell_3841 ( .C (clk), .D (signal_1501), .Q (signal_6387) ) ;
    buf_clk cell_3857 ( .C (clk), .D (signal_756), .Q (signal_6403) ) ;
    buf_clk cell_3873 ( .C (clk), .D (signal_1749), .Q (signal_6419) ) ;
    buf_clk cell_3889 ( .C (clk), .D (signal_3106), .Q (signal_6435) ) ;
    buf_clk cell_3905 ( .C (clk), .D (signal_748), .Q (signal_6451) ) ;
    buf_clk cell_3921 ( .C (clk), .D (signal_1765), .Q (signal_6467) ) ;
    buf_clk cell_3937 ( .C (clk), .D (signal_3131), .Q (signal_6483) ) ;
    buf_clk cell_3953 ( .C (clk), .D (signal_1748), .Q (signal_6499) ) ;
    buf_clk cell_3969 ( .C (clk), .D (signal_3109), .Q (signal_6515) ) ;
    buf_clk cell_3985 ( .C (clk), .D (signal_1764), .Q (signal_6531) ) ;
    buf_clk cell_4001 ( .C (clk), .D (signal_3134), .Q (signal_6547) ) ;
    buf_clk cell_4017 ( .C (clk), .D (signal_1747), .Q (signal_6563) ) ;
    buf_clk cell_4033 ( .C (clk), .D (signal_3112), .Q (signal_6579) ) ;
    buf_clk cell_4049 ( .C (clk), .D (signal_1763), .Q (signal_6595) ) ;
    buf_clk cell_4065 ( .C (clk), .D (signal_3137), .Q (signal_6611) ) ;
    buf_clk cell_4081 ( .C (clk), .D (signal_1746), .Q (signal_6627) ) ;
    buf_clk cell_4097 ( .C (clk), .D (signal_3115), .Q (signal_6643) ) ;
    buf_clk cell_4113 ( .C (clk), .D (signal_1762), .Q (signal_6659) ) ;
    buf_clk cell_4129 ( .C (clk), .D (signal_3140), .Q (signal_6675) ) ;
    buf_clk cell_4145 ( .C (clk), .D (signal_1745), .Q (signal_6691) ) ;
    buf_clk cell_4161 ( .C (clk), .D (signal_3118), .Q (signal_6707) ) ;
    buf_clk cell_4177 ( .C (clk), .D (signal_1761), .Q (signal_6723) ) ;
    buf_clk cell_4193 ( .C (clk), .D (signal_3143), .Q (signal_6739) ) ;
    buf_clk cell_4209 ( .C (clk), .D (signal_1744), .Q (signal_6755) ) ;
    buf_clk cell_4225 ( .C (clk), .D (signal_3121), .Q (signal_6771) ) ;
    buf_clk cell_4241 ( .C (clk), .D (signal_1760), .Q (signal_6787) ) ;
    buf_clk cell_4257 ( .C (clk), .D (signal_3146), .Q (signal_6803) ) ;
    buf_clk cell_4273 ( .C (clk), .D (signal_1743), .Q (signal_6819) ) ;
    buf_clk cell_4289 ( .C (clk), .D (signal_3124), .Q (signal_6835) ) ;
    buf_clk cell_4305 ( .C (clk), .D (signal_1759), .Q (signal_6851) ) ;
    buf_clk cell_4321 ( .C (clk), .D (signal_3149), .Q (signal_6867) ) ;
    buf_clk cell_4337 ( .C (clk), .D (signal_1742), .Q (signal_6883) ) ;
    buf_clk cell_4353 ( .C (clk), .D (signal_3127), .Q (signal_6899) ) ;
    buf_clk cell_4369 ( .C (clk), .D (signal_1758), .Q (signal_6915) ) ;
    buf_clk cell_4385 ( .C (clk), .D (signal_3152), .Q (signal_6931) ) ;
    buf_clk cell_4401 ( .C (clk), .D (signal_1517), .Q (signal_6947) ) ;
    buf_clk cell_4415 ( .C (clk), .D (signal_3249), .Q (signal_6961) ) ;
    buf_clk cell_4429 ( .C (clk), .D (signal_429), .Q (signal_6975) ) ;
    buf_clk cell_4445 ( .C (clk), .D (signal_431), .Q (signal_6991) ) ;
    buf_clk cell_4461 ( .C (clk), .D (signal_433), .Q (signal_7007) ) ;
    buf_clk cell_4477 ( .C (clk), .D (signal_435), .Q (signal_7023) ) ;
    buf_clk cell_4493 ( .C (clk), .D (signal_437), .Q (signal_7039) ) ;
    buf_clk cell_4509 ( .C (clk), .D (signal_439), .Q (signal_7055) ) ;
    buf_clk cell_4525 ( .C (clk), .D (signal_441), .Q (signal_7071) ) ;
    buf_clk cell_4541 ( .C (clk), .D (signal_419), .Q (signal_7087) ) ;
    buf_clk cell_4557 ( .C (clk), .D (signal_395), .Q (signal_7103) ) ;
    buf_clk cell_4573 ( .C (clk), .D (signal_465), .Q (signal_7119) ) ;
    buf_clk cell_4589 ( .C (clk), .D (signal_3820), .Q (signal_7135) ) ;
    buf_clk cell_4605 ( .C (clk), .D (signal_467), .Q (signal_7151) ) ;
    buf_clk cell_4621 ( .C (clk), .D (signal_3821), .Q (signal_7167) ) ;
    buf_clk cell_4637 ( .C (clk), .D (signal_469), .Q (signal_7183) ) ;
    buf_clk cell_4653 ( .C (clk), .D (signal_3822), .Q (signal_7199) ) ;
    buf_clk cell_4669 ( .C (clk), .D (signal_471), .Q (signal_7215) ) ;
    buf_clk cell_4685 ( .C (clk), .D (signal_3823), .Q (signal_7231) ) ;
    buf_clk cell_4701 ( .C (clk), .D (signal_473), .Q (signal_7247) ) ;
    buf_clk cell_4717 ( .C (clk), .D (signal_3824), .Q (signal_7263) ) ;
    buf_clk cell_4733 ( .C (clk), .D (signal_475), .Q (signal_7279) ) ;
    buf_clk cell_4749 ( .C (clk), .D (signal_3825), .Q (signal_7295) ) ;
    buf_clk cell_4765 ( .C (clk), .D (signal_477), .Q (signal_7311) ) ;
    buf_clk cell_4781 ( .C (clk), .D (signal_3826), .Q (signal_7327) ) ;
    buf_clk cell_4797 ( .C (clk), .D (signal_479), .Q (signal_7343) ) ;
    buf_clk cell_4813 ( .C (clk), .D (signal_3827), .Q (signal_7359) ) ;
    buf_clk cell_4829 ( .C (clk), .D (signal_481), .Q (signal_7375) ) ;
    buf_clk cell_4845 ( .C (clk), .D (signal_3828), .Q (signal_7391) ) ;
    buf_clk cell_4861 ( .C (clk), .D (signal_483), .Q (signal_7407) ) ;
    buf_clk cell_4877 ( .C (clk), .D (signal_3829), .Q (signal_7423) ) ;
    buf_clk cell_4893 ( .C (clk), .D (signal_485), .Q (signal_7439) ) ;
    buf_clk cell_4909 ( .C (clk), .D (signal_3830), .Q (signal_7455) ) ;
    buf_clk cell_4925 ( .C (clk), .D (signal_487), .Q (signal_7471) ) ;
    buf_clk cell_4941 ( .C (clk), .D (signal_3831), .Q (signal_7487) ) ;
    buf_clk cell_4957 ( .C (clk), .D (signal_489), .Q (signal_7503) ) ;
    buf_clk cell_4973 ( .C (clk), .D (signal_3832), .Q (signal_7519) ) ;
    buf_clk cell_4989 ( .C (clk), .D (signal_491), .Q (signal_7535) ) ;
    buf_clk cell_5005 ( .C (clk), .D (signal_3833), .Q (signal_7551) ) ;
    buf_clk cell_5021 ( .C (clk), .D (signal_493), .Q (signal_7567) ) ;
    buf_clk cell_5037 ( .C (clk), .D (signal_3834), .Q (signal_7583) ) ;
    buf_clk cell_5053 ( .C (clk), .D (signal_495), .Q (signal_7599) ) ;
    buf_clk cell_5069 ( .C (clk), .D (signal_3835), .Q (signal_7615) ) ;
    buf_clk cell_5085 ( .C (clk), .D (signal_497), .Q (signal_7631) ) ;
    buf_clk cell_5101 ( .C (clk), .D (signal_3836), .Q (signal_7647) ) ;
    buf_clk cell_5117 ( .C (clk), .D (signal_499), .Q (signal_7663) ) ;
    buf_clk cell_5133 ( .C (clk), .D (signal_3837), .Q (signal_7679) ) ;
    buf_clk cell_5149 ( .C (clk), .D (signal_501), .Q (signal_7695) ) ;
    buf_clk cell_5165 ( .C (clk), .D (signal_3838), .Q (signal_7711) ) ;
    buf_clk cell_5181 ( .C (clk), .D (signal_503), .Q (signal_7727) ) ;
    buf_clk cell_5197 ( .C (clk), .D (signal_3839), .Q (signal_7743) ) ;
    buf_clk cell_5213 ( .C (clk), .D (signal_505), .Q (signal_7759) ) ;
    buf_clk cell_5229 ( .C (clk), .D (signal_3840), .Q (signal_7775) ) ;
    buf_clk cell_5245 ( .C (clk), .D (signal_507), .Q (signal_7791) ) ;
    buf_clk cell_5261 ( .C (clk), .D (signal_3841), .Q (signal_7807) ) ;
    buf_clk cell_5277 ( .C (clk), .D (signal_509), .Q (signal_7823) ) ;
    buf_clk cell_5293 ( .C (clk), .D (signal_3842), .Q (signal_7839) ) ;
    buf_clk cell_5309 ( .C (clk), .D (signal_511), .Q (signal_7855) ) ;
    buf_clk cell_5325 ( .C (clk), .D (signal_3843), .Q (signal_7871) ) ;
    buf_clk cell_5341 ( .C (clk), .D (signal_513), .Q (signal_7887) ) ;
    buf_clk cell_5357 ( .C (clk), .D (signal_3844), .Q (signal_7903) ) ;
    buf_clk cell_5373 ( .C (clk), .D (signal_515), .Q (signal_7919) ) ;
    buf_clk cell_5389 ( .C (clk), .D (signal_3845), .Q (signal_7935) ) ;
    buf_clk cell_5405 ( .C (clk), .D (signal_517), .Q (signal_7951) ) ;
    buf_clk cell_5421 ( .C (clk), .D (signal_3846), .Q (signal_7967) ) ;
    buf_clk cell_5437 ( .C (clk), .D (signal_519), .Q (signal_7983) ) ;
    buf_clk cell_5453 ( .C (clk), .D (signal_3847), .Q (signal_7999) ) ;
    buf_clk cell_5469 ( .C (clk), .D (signal_521), .Q (signal_8015) ) ;
    buf_clk cell_5485 ( .C (clk), .D (signal_3848), .Q (signal_8031) ) ;
    buf_clk cell_5501 ( .C (clk), .D (signal_523), .Q (signal_8047) ) ;
    buf_clk cell_5517 ( .C (clk), .D (signal_3849), .Q (signal_8063) ) ;
    buf_clk cell_5533 ( .C (clk), .D (signal_525), .Q (signal_8079) ) ;
    buf_clk cell_5549 ( .C (clk), .D (signal_3850), .Q (signal_8095) ) ;
    buf_clk cell_5565 ( .C (clk), .D (signal_527), .Q (signal_8111) ) ;
    buf_clk cell_5581 ( .C (clk), .D (signal_3851), .Q (signal_8127) ) ;
    buf_clk cell_5597 ( .C (clk), .D (signal_529), .Q (signal_8143) ) ;
    buf_clk cell_5613 ( .C (clk), .D (signal_3852), .Q (signal_8159) ) ;
    buf_clk cell_5629 ( .C (clk), .D (signal_531), .Q (signal_8175) ) ;
    buf_clk cell_5645 ( .C (clk), .D (signal_3853), .Q (signal_8191) ) ;
    buf_clk cell_5661 ( .C (clk), .D (signal_533), .Q (signal_8207) ) ;
    buf_clk cell_5677 ( .C (clk), .D (signal_3854), .Q (signal_8223) ) ;
    buf_clk cell_5693 ( .C (clk), .D (signal_535), .Q (signal_8239) ) ;
    buf_clk cell_5709 ( .C (clk), .D (signal_3855), .Q (signal_8255) ) ;
    buf_clk cell_5725 ( .C (clk), .D (signal_537), .Q (signal_8271) ) ;
    buf_clk cell_5741 ( .C (clk), .D (signal_3856), .Q (signal_8287) ) ;
    buf_clk cell_5757 ( .C (clk), .D (signal_539), .Q (signal_8303) ) ;
    buf_clk cell_5773 ( .C (clk), .D (signal_3857), .Q (signal_8319) ) ;
    buf_clk cell_5789 ( .C (clk), .D (signal_541), .Q (signal_8335) ) ;
    buf_clk cell_5805 ( .C (clk), .D (signal_3858), .Q (signal_8351) ) ;
    buf_clk cell_5821 ( .C (clk), .D (signal_543), .Q (signal_8367) ) ;
    buf_clk cell_5837 ( .C (clk), .D (signal_3859), .Q (signal_8383) ) ;
    buf_clk cell_5853 ( .C (clk), .D (signal_545), .Q (signal_8399) ) ;
    buf_clk cell_5869 ( .C (clk), .D (signal_3860), .Q (signal_8415) ) ;
    buf_clk cell_5885 ( .C (clk), .D (signal_547), .Q (signal_8431) ) ;
    buf_clk cell_5901 ( .C (clk), .D (signal_3861), .Q (signal_8447) ) ;
    buf_clk cell_5917 ( .C (clk), .D (signal_549), .Q (signal_8463) ) ;
    buf_clk cell_5933 ( .C (clk), .D (signal_3862), .Q (signal_8479) ) ;
    buf_clk cell_5949 ( .C (clk), .D (signal_551), .Q (signal_8495) ) ;
    buf_clk cell_5965 ( .C (clk), .D (signal_3863), .Q (signal_8511) ) ;
    buf_clk cell_5981 ( .C (clk), .D (signal_553), .Q (signal_8527) ) ;
    buf_clk cell_5997 ( .C (clk), .D (signal_3864), .Q (signal_8543) ) ;
    buf_clk cell_6013 ( .C (clk), .D (signal_555), .Q (signal_8559) ) ;
    buf_clk cell_6029 ( .C (clk), .D (signal_3865), .Q (signal_8575) ) ;
    buf_clk cell_6045 ( .C (clk), .D (signal_557), .Q (signal_8591) ) ;
    buf_clk cell_6061 ( .C (clk), .D (signal_3866), .Q (signal_8607) ) ;
    buf_clk cell_6077 ( .C (clk), .D (signal_559), .Q (signal_8623) ) ;
    buf_clk cell_6093 ( .C (clk), .D (signal_3867), .Q (signal_8639) ) ;
    buf_clk cell_6109 ( .C (clk), .D (signal_561), .Q (signal_8655) ) ;
    buf_clk cell_6125 ( .C (clk), .D (signal_3868), .Q (signal_8671) ) ;
    buf_clk cell_6141 ( .C (clk), .D (signal_563), .Q (signal_8687) ) ;
    buf_clk cell_6157 ( .C (clk), .D (signal_3869), .Q (signal_8703) ) ;
    buf_clk cell_6173 ( .C (clk), .D (signal_565), .Q (signal_8719) ) ;
    buf_clk cell_6189 ( .C (clk), .D (signal_3870), .Q (signal_8735) ) ;
    buf_clk cell_6205 ( .C (clk), .D (signal_567), .Q (signal_8751) ) ;
    buf_clk cell_6221 ( .C (clk), .D (signal_3871), .Q (signal_8767) ) ;
    buf_clk cell_6237 ( .C (clk), .D (signal_569), .Q (signal_8783) ) ;
    buf_clk cell_6253 ( .C (clk), .D (signal_3872), .Q (signal_8799) ) ;
    buf_clk cell_6269 ( .C (clk), .D (signal_571), .Q (signal_8815) ) ;
    buf_clk cell_6285 ( .C (clk), .D (signal_3873), .Q (signal_8831) ) ;
    buf_clk cell_6301 ( .C (clk), .D (signal_573), .Q (signal_8847) ) ;
    buf_clk cell_6317 ( .C (clk), .D (signal_3874), .Q (signal_8863) ) ;
    buf_clk cell_6333 ( .C (clk), .D (signal_575), .Q (signal_8879) ) ;
    buf_clk cell_6349 ( .C (clk), .D (signal_3875), .Q (signal_8895) ) ;
    buf_clk cell_6365 ( .C (clk), .D (signal_577), .Q (signal_8911) ) ;
    buf_clk cell_6381 ( .C (clk), .D (signal_3876), .Q (signal_8927) ) ;
    buf_clk cell_6397 ( .C (clk), .D (signal_579), .Q (signal_8943) ) ;
    buf_clk cell_6413 ( .C (clk), .D (signal_3877), .Q (signal_8959) ) ;
    buf_clk cell_6429 ( .C (clk), .D (signal_581), .Q (signal_8975) ) ;
    buf_clk cell_6445 ( .C (clk), .D (signal_3878), .Q (signal_8991) ) ;
    buf_clk cell_6461 ( .C (clk), .D (signal_583), .Q (signal_9007) ) ;
    buf_clk cell_6477 ( .C (clk), .D (signal_3879), .Q (signal_9023) ) ;
    buf_clk cell_6493 ( .C (clk), .D (signal_585), .Q (signal_9039) ) ;
    buf_clk cell_6509 ( .C (clk), .D (signal_3880), .Q (signal_9055) ) ;
    buf_clk cell_6525 ( .C (clk), .D (signal_587), .Q (signal_9071) ) ;
    buf_clk cell_6541 ( .C (clk), .D (signal_3881), .Q (signal_9087) ) ;
    buf_clk cell_6557 ( .C (clk), .D (signal_589), .Q (signal_9103) ) ;
    buf_clk cell_6573 ( .C (clk), .D (signal_3882), .Q (signal_9119) ) ;
    buf_clk cell_6589 ( .C (clk), .D (signal_591), .Q (signal_9135) ) ;
    buf_clk cell_6605 ( .C (clk), .D (signal_3883), .Q (signal_9151) ) ;
    buf_clk cell_6621 ( .C (clk), .D (signal_593), .Q (signal_9167) ) ;
    buf_clk cell_6637 ( .C (clk), .D (signal_3884), .Q (signal_9183) ) ;
    buf_clk cell_6653 ( .C (clk), .D (signal_595), .Q (signal_9199) ) ;
    buf_clk cell_6669 ( .C (clk), .D (signal_3885), .Q (signal_9215) ) ;
    buf_clk cell_6685 ( .C (clk), .D (signal_597), .Q (signal_9231) ) ;
    buf_clk cell_6701 ( .C (clk), .D (signal_3886), .Q (signal_9247) ) ;
    buf_clk cell_6717 ( .C (clk), .D (signal_599), .Q (signal_9263) ) ;
    buf_clk cell_6733 ( .C (clk), .D (signal_3887), .Q (signal_9279) ) ;
    buf_clk cell_6749 ( .C (clk), .D (signal_601), .Q (signal_9295) ) ;
    buf_clk cell_6765 ( .C (clk), .D (signal_3888), .Q (signal_9311) ) ;
    buf_clk cell_6781 ( .C (clk), .D (signal_603), .Q (signal_9327) ) ;
    buf_clk cell_6797 ( .C (clk), .D (signal_3889), .Q (signal_9343) ) ;
    buf_clk cell_6813 ( .C (clk), .D (signal_605), .Q (signal_9359) ) ;
    buf_clk cell_6829 ( .C (clk), .D (signal_3890), .Q (signal_9375) ) ;
    buf_clk cell_6845 ( .C (clk), .D (signal_607), .Q (signal_9391) ) ;
    buf_clk cell_6861 ( .C (clk), .D (signal_3891), .Q (signal_9407) ) ;
    buf_clk cell_6877 ( .C (clk), .D (signal_609), .Q (signal_9423) ) ;
    buf_clk cell_6893 ( .C (clk), .D (signal_3892), .Q (signal_9439) ) ;
    buf_clk cell_6909 ( .C (clk), .D (signal_611), .Q (signal_9455) ) ;
    buf_clk cell_6925 ( .C (clk), .D (signal_3893), .Q (signal_9471) ) ;
    buf_clk cell_6941 ( .C (clk), .D (signal_613), .Q (signal_9487) ) ;
    buf_clk cell_6957 ( .C (clk), .D (signal_3894), .Q (signal_9503) ) ;
    buf_clk cell_6973 ( .C (clk), .D (signal_615), .Q (signal_9519) ) ;
    buf_clk cell_6989 ( .C (clk), .D (signal_3895), .Q (signal_9535) ) ;
    buf_clk cell_7005 ( .C (clk), .D (signal_617), .Q (signal_9551) ) ;
    buf_clk cell_7021 ( .C (clk), .D (signal_3896), .Q (signal_9567) ) ;
    buf_clk cell_7037 ( .C (clk), .D (signal_619), .Q (signal_9583) ) ;
    buf_clk cell_7053 ( .C (clk), .D (signal_3897), .Q (signal_9599) ) ;
    buf_clk cell_7069 ( .C (clk), .D (signal_621), .Q (signal_9615) ) ;
    buf_clk cell_7085 ( .C (clk), .D (signal_3898), .Q (signal_9631) ) ;
    buf_clk cell_7101 ( .C (clk), .D (signal_623), .Q (signal_9647) ) ;
    buf_clk cell_7117 ( .C (clk), .D (signal_3899), .Q (signal_9663) ) ;
    buf_clk cell_7133 ( .C (clk), .D (signal_625), .Q (signal_9679) ) ;
    buf_clk cell_7149 ( .C (clk), .D (signal_3900), .Q (signal_9695) ) ;
    buf_clk cell_7165 ( .C (clk), .D (signal_627), .Q (signal_9711) ) ;
    buf_clk cell_7181 ( .C (clk), .D (signal_3901), .Q (signal_9727) ) ;
    buf_clk cell_7197 ( .C (clk), .D (signal_629), .Q (signal_9743) ) ;
    buf_clk cell_7213 ( .C (clk), .D (signal_3902), .Q (signal_9759) ) ;
    buf_clk cell_7229 ( .C (clk), .D (signal_631), .Q (signal_9775) ) ;
    buf_clk cell_7245 ( .C (clk), .D (signal_3903), .Q (signal_9791) ) ;
    buf_clk cell_7261 ( .C (clk), .D (signal_633), .Q (signal_9807) ) ;
    buf_clk cell_7277 ( .C (clk), .D (signal_3904), .Q (signal_9823) ) ;
    buf_clk cell_7293 ( .C (clk), .D (signal_635), .Q (signal_9839) ) ;
    buf_clk cell_7309 ( .C (clk), .D (signal_3905), .Q (signal_9855) ) ;
    buf_clk cell_7325 ( .C (clk), .D (signal_637), .Q (signal_9871) ) ;
    buf_clk cell_7341 ( .C (clk), .D (signal_3906), .Q (signal_9887) ) ;
    buf_clk cell_7357 ( .C (clk), .D (signal_639), .Q (signal_9903) ) ;
    buf_clk cell_7373 ( .C (clk), .D (signal_3907), .Q (signal_9919) ) ;
    buf_clk cell_7389 ( .C (clk), .D (signal_641), .Q (signal_9935) ) ;
    buf_clk cell_7405 ( .C (clk), .D (signal_3908), .Q (signal_9951) ) ;
    buf_clk cell_7421 ( .C (clk), .D (signal_643), .Q (signal_9967) ) ;
    buf_clk cell_7437 ( .C (clk), .D (signal_3909), .Q (signal_9983) ) ;
    buf_clk cell_7453 ( .C (clk), .D (signal_645), .Q (signal_9999) ) ;
    buf_clk cell_7469 ( .C (clk), .D (signal_3910), .Q (signal_10015) ) ;
    buf_clk cell_7485 ( .C (clk), .D (signal_647), .Q (signal_10031) ) ;
    buf_clk cell_7501 ( .C (clk), .D (signal_3911), .Q (signal_10047) ) ;
    buf_clk cell_7517 ( .C (clk), .D (signal_649), .Q (signal_10063) ) ;
    buf_clk cell_7533 ( .C (clk), .D (signal_3912), .Q (signal_10079) ) ;
    buf_clk cell_7549 ( .C (clk), .D (signal_651), .Q (signal_10095) ) ;
    buf_clk cell_7565 ( .C (clk), .D (signal_3913), .Q (signal_10111) ) ;
    buf_clk cell_7581 ( .C (clk), .D (signal_653), .Q (signal_10127) ) ;
    buf_clk cell_7597 ( .C (clk), .D (signal_3914), .Q (signal_10143) ) ;
    buf_clk cell_7613 ( .C (clk), .D (signal_655), .Q (signal_10159) ) ;
    buf_clk cell_7629 ( .C (clk), .D (signal_3915), .Q (signal_10175) ) ;
    buf_clk cell_7645 ( .C (clk), .D (signal_657), .Q (signal_10191) ) ;
    buf_clk cell_7661 ( .C (clk), .D (signal_3916), .Q (signal_10207) ) ;
    buf_clk cell_7677 ( .C (clk), .D (signal_659), .Q (signal_10223) ) ;
    buf_clk cell_7693 ( .C (clk), .D (signal_3917), .Q (signal_10239) ) ;
    buf_clk cell_7709 ( .C (clk), .D (signal_661), .Q (signal_10255) ) ;
    buf_clk cell_7725 ( .C (clk), .D (signal_3918), .Q (signal_10271) ) ;
    buf_clk cell_7741 ( .C (clk), .D (signal_663), .Q (signal_10287) ) ;
    buf_clk cell_7757 ( .C (clk), .D (signal_3919), .Q (signal_10303) ) ;
    buf_clk cell_7773 ( .C (clk), .D (signal_665), .Q (signal_10319) ) ;
    buf_clk cell_7789 ( .C (clk), .D (signal_3920), .Q (signal_10335) ) ;
    buf_clk cell_7805 ( .C (clk), .D (signal_667), .Q (signal_10351) ) ;
    buf_clk cell_7821 ( .C (clk), .D (signal_3921), .Q (signal_10367) ) ;
    buf_clk cell_7837 ( .C (clk), .D (signal_669), .Q (signal_10383) ) ;
    buf_clk cell_7853 ( .C (clk), .D (signal_3922), .Q (signal_10399) ) ;
    buf_clk cell_7869 ( .C (clk), .D (signal_671), .Q (signal_10415) ) ;
    buf_clk cell_7885 ( .C (clk), .D (signal_3923), .Q (signal_10431) ) ;
    buf_clk cell_7901 ( .C (clk), .D (signal_673), .Q (signal_10447) ) ;
    buf_clk cell_7917 ( .C (clk), .D (signal_3924), .Q (signal_10463) ) ;
    buf_clk cell_7933 ( .C (clk), .D (signal_675), .Q (signal_10479) ) ;
    buf_clk cell_7949 ( .C (clk), .D (signal_3925), .Q (signal_10495) ) ;
    buf_clk cell_7965 ( .C (clk), .D (signal_677), .Q (signal_10511) ) ;
    buf_clk cell_7981 ( .C (clk), .D (signal_3926), .Q (signal_10527) ) ;
    buf_clk cell_7997 ( .C (clk), .D (signal_679), .Q (signal_10543) ) ;
    buf_clk cell_8013 ( .C (clk), .D (signal_3927), .Q (signal_10559) ) ;
    buf_clk cell_8029 ( .C (clk), .D (signal_681), .Q (signal_10575) ) ;
    buf_clk cell_8045 ( .C (clk), .D (signal_3928), .Q (signal_10591) ) ;
    buf_clk cell_8061 ( .C (clk), .D (signal_683), .Q (signal_10607) ) ;
    buf_clk cell_8077 ( .C (clk), .D (signal_3929), .Q (signal_10623) ) ;
    buf_clk cell_8093 ( .C (clk), .D (signal_685), .Q (signal_10639) ) ;
    buf_clk cell_8109 ( .C (clk), .D (signal_3930), .Q (signal_10655) ) ;
    buf_clk cell_8125 ( .C (clk), .D (signal_687), .Q (signal_10671) ) ;
    buf_clk cell_8141 ( .C (clk), .D (signal_3931), .Q (signal_10687) ) ;
    buf_clk cell_8157 ( .C (clk), .D (signal_689), .Q (signal_10703) ) ;
    buf_clk cell_8173 ( .C (clk), .D (signal_3932), .Q (signal_10719) ) ;
    buf_clk cell_8189 ( .C (clk), .D (signal_691), .Q (signal_10735) ) ;
    buf_clk cell_8205 ( .C (clk), .D (signal_3933), .Q (signal_10751) ) ;
    buf_clk cell_8221 ( .C (clk), .D (signal_693), .Q (signal_10767) ) ;
    buf_clk cell_8237 ( .C (clk), .D (signal_3934), .Q (signal_10783) ) ;
    buf_clk cell_8253 ( .C (clk), .D (signal_695), .Q (signal_10799) ) ;
    buf_clk cell_8269 ( .C (clk), .D (signal_3935), .Q (signal_10815) ) ;
    buf_clk cell_8285 ( .C (clk), .D (signal_697), .Q (signal_10831) ) ;
    buf_clk cell_8301 ( .C (clk), .D (signal_3936), .Q (signal_10847) ) ;
    buf_clk cell_8317 ( .C (clk), .D (signal_699), .Q (signal_10863) ) ;
    buf_clk cell_8333 ( .C (clk), .D (signal_3937), .Q (signal_10879) ) ;
    buf_clk cell_8349 ( .C (clk), .D (signal_701), .Q (signal_10895) ) ;
    buf_clk cell_8365 ( .C (clk), .D (signal_3938), .Q (signal_10911) ) ;
    buf_clk cell_8381 ( .C (clk), .D (signal_703), .Q (signal_10927) ) ;
    buf_clk cell_8397 ( .C (clk), .D (signal_3939), .Q (signal_10943) ) ;
    buf_clk cell_8413 ( .C (clk), .D (signal_766), .Q (signal_10959) ) ;
    buf_clk cell_8429 ( .C (clk), .D (signal_4156), .Q (signal_10975) ) ;
    buf_clk cell_8445 ( .C (clk), .D (signal_769), .Q (signal_10991) ) ;
    buf_clk cell_8461 ( .C (clk), .D (signal_4157), .Q (signal_11007) ) ;
    buf_clk cell_8477 ( .C (clk), .D (signal_772), .Q (signal_11023) ) ;
    buf_clk cell_8493 ( .C (clk), .D (signal_4158), .Q (signal_11039) ) ;
    buf_clk cell_8509 ( .C (clk), .D (signal_775), .Q (signal_11055) ) ;
    buf_clk cell_8525 ( .C (clk), .D (signal_4159), .Q (signal_11071) ) ;
    buf_clk cell_8541 ( .C (clk), .D (signal_778), .Q (signal_11087) ) ;
    buf_clk cell_8557 ( .C (clk), .D (signal_4160), .Q (signal_11103) ) ;
    buf_clk cell_8573 ( .C (clk), .D (signal_781), .Q (signal_11119) ) ;
    buf_clk cell_8589 ( .C (clk), .D (signal_4161), .Q (signal_11135) ) ;
    buf_clk cell_8605 ( .C (clk), .D (signal_784), .Q (signal_11151) ) ;
    buf_clk cell_8621 ( .C (clk), .D (signal_4162), .Q (signal_11167) ) ;
    buf_clk cell_8637 ( .C (clk), .D (signal_787), .Q (signal_11183) ) ;
    buf_clk cell_8653 ( .C (clk), .D (signal_4163), .Q (signal_11199) ) ;
    buf_clk cell_8669 ( .C (clk), .D (signal_790), .Q (signal_11215) ) ;
    buf_clk cell_8685 ( .C (clk), .D (signal_4028), .Q (signal_11231) ) ;
    buf_clk cell_8701 ( .C (clk), .D (signal_793), .Q (signal_11247) ) ;
    buf_clk cell_8717 ( .C (clk), .D (signal_4029), .Q (signal_11263) ) ;
    buf_clk cell_8733 ( .C (clk), .D (signal_796), .Q (signal_11279) ) ;
    buf_clk cell_8749 ( .C (clk), .D (signal_4030), .Q (signal_11295) ) ;
    buf_clk cell_8765 ( .C (clk), .D (signal_799), .Q (signal_11311) ) ;
    buf_clk cell_8781 ( .C (clk), .D (signal_4031), .Q (signal_11327) ) ;
    buf_clk cell_8797 ( .C (clk), .D (signal_802), .Q (signal_11343) ) ;
    buf_clk cell_8813 ( .C (clk), .D (signal_4032), .Q (signal_11359) ) ;
    buf_clk cell_8829 ( .C (clk), .D (signal_805), .Q (signal_11375) ) ;
    buf_clk cell_8845 ( .C (clk), .D (signal_4033), .Q (signal_11391) ) ;
    buf_clk cell_8861 ( .C (clk), .D (signal_808), .Q (signal_11407) ) ;
    buf_clk cell_8877 ( .C (clk), .D (signal_4034), .Q (signal_11423) ) ;
    buf_clk cell_8893 ( .C (clk), .D (signal_811), .Q (signal_11439) ) ;
    buf_clk cell_8909 ( .C (clk), .D (signal_4035), .Q (signal_11455) ) ;
    buf_clk cell_8925 ( .C (clk), .D (signal_814), .Q (signal_11471) ) ;
    buf_clk cell_8941 ( .C (clk), .D (signal_4036), .Q (signal_11487) ) ;
    buf_clk cell_8957 ( .C (clk), .D (signal_817), .Q (signal_11503) ) ;
    buf_clk cell_8973 ( .C (clk), .D (signal_4037), .Q (signal_11519) ) ;
    buf_clk cell_8989 ( .C (clk), .D (signal_820), .Q (signal_11535) ) ;
    buf_clk cell_9005 ( .C (clk), .D (signal_4038), .Q (signal_11551) ) ;
    buf_clk cell_9021 ( .C (clk), .D (signal_823), .Q (signal_11567) ) ;
    buf_clk cell_9037 ( .C (clk), .D (signal_4039), .Q (signal_11583) ) ;
    buf_clk cell_9053 ( .C (clk), .D (signal_826), .Q (signal_11599) ) ;
    buf_clk cell_9069 ( .C (clk), .D (signal_4040), .Q (signal_11615) ) ;
    buf_clk cell_9085 ( .C (clk), .D (signal_829), .Q (signal_11631) ) ;
    buf_clk cell_9101 ( .C (clk), .D (signal_4041), .Q (signal_11647) ) ;
    buf_clk cell_9117 ( .C (clk), .D (signal_832), .Q (signal_11663) ) ;
    buf_clk cell_9133 ( .C (clk), .D (signal_4042), .Q (signal_11679) ) ;
    buf_clk cell_9149 ( .C (clk), .D (signal_835), .Q (signal_11695) ) ;
    buf_clk cell_9165 ( .C (clk), .D (signal_4043), .Q (signal_11711) ) ;
    buf_clk cell_9181 ( .C (clk), .D (signal_838), .Q (signal_11727) ) ;
    buf_clk cell_9197 ( .C (clk), .D (signal_4044), .Q (signal_11743) ) ;
    buf_clk cell_9213 ( .C (clk), .D (signal_841), .Q (signal_11759) ) ;
    buf_clk cell_9229 ( .C (clk), .D (signal_4045), .Q (signal_11775) ) ;
    buf_clk cell_9245 ( .C (clk), .D (signal_844), .Q (signal_11791) ) ;
    buf_clk cell_9261 ( .C (clk), .D (signal_4046), .Q (signal_11807) ) ;
    buf_clk cell_9277 ( .C (clk), .D (signal_847), .Q (signal_11823) ) ;
    buf_clk cell_9293 ( .C (clk), .D (signal_4047), .Q (signal_11839) ) ;
    buf_clk cell_9309 ( .C (clk), .D (signal_850), .Q (signal_11855) ) ;
    buf_clk cell_9325 ( .C (clk), .D (signal_4048), .Q (signal_11871) ) ;
    buf_clk cell_9341 ( .C (clk), .D (signal_853), .Q (signal_11887) ) ;
    buf_clk cell_9357 ( .C (clk), .D (signal_4049), .Q (signal_11903) ) ;
    buf_clk cell_9373 ( .C (clk), .D (signal_856), .Q (signal_11919) ) ;
    buf_clk cell_9389 ( .C (clk), .D (signal_4050), .Q (signal_11935) ) ;
    buf_clk cell_9405 ( .C (clk), .D (signal_859), .Q (signal_11951) ) ;
    buf_clk cell_9421 ( .C (clk), .D (signal_4051), .Q (signal_11967) ) ;
    buf_clk cell_9437 ( .C (clk), .D (signal_862), .Q (signal_11983) ) ;
    buf_clk cell_9453 ( .C (clk), .D (signal_4052), .Q (signal_11999) ) ;
    buf_clk cell_9469 ( .C (clk), .D (signal_865), .Q (signal_12015) ) ;
    buf_clk cell_9485 ( .C (clk), .D (signal_4053), .Q (signal_12031) ) ;
    buf_clk cell_9501 ( .C (clk), .D (signal_868), .Q (signal_12047) ) ;
    buf_clk cell_9517 ( .C (clk), .D (signal_4054), .Q (signal_12063) ) ;
    buf_clk cell_9533 ( .C (clk), .D (signal_871), .Q (signal_12079) ) ;
    buf_clk cell_9549 ( .C (clk), .D (signal_4055), .Q (signal_12095) ) ;
    buf_clk cell_9565 ( .C (clk), .D (signal_874), .Q (signal_12111) ) ;
    buf_clk cell_9581 ( .C (clk), .D (signal_4056), .Q (signal_12127) ) ;
    buf_clk cell_9597 ( .C (clk), .D (signal_877), .Q (signal_12143) ) ;
    buf_clk cell_9613 ( .C (clk), .D (signal_4057), .Q (signal_12159) ) ;
    buf_clk cell_9629 ( .C (clk), .D (signal_880), .Q (signal_12175) ) ;
    buf_clk cell_9645 ( .C (clk), .D (signal_4058), .Q (signal_12191) ) ;
    buf_clk cell_9661 ( .C (clk), .D (signal_883), .Q (signal_12207) ) ;
    buf_clk cell_9677 ( .C (clk), .D (signal_4059), .Q (signal_12223) ) ;
    buf_clk cell_9693 ( .C (clk), .D (signal_886), .Q (signal_12239) ) ;
    buf_clk cell_9709 ( .C (clk), .D (signal_4060), .Q (signal_12255) ) ;
    buf_clk cell_9725 ( .C (clk), .D (signal_889), .Q (signal_12271) ) ;
    buf_clk cell_9741 ( .C (clk), .D (signal_4061), .Q (signal_12287) ) ;
    buf_clk cell_9757 ( .C (clk), .D (signal_892), .Q (signal_12303) ) ;
    buf_clk cell_9773 ( .C (clk), .D (signal_4062), .Q (signal_12319) ) ;
    buf_clk cell_9789 ( .C (clk), .D (signal_895), .Q (signal_12335) ) ;
    buf_clk cell_9805 ( .C (clk), .D (signal_4063), .Q (signal_12351) ) ;
    buf_clk cell_9821 ( .C (clk), .D (signal_898), .Q (signal_12367) ) ;
    buf_clk cell_9837 ( .C (clk), .D (signal_4064), .Q (signal_12383) ) ;
    buf_clk cell_9853 ( .C (clk), .D (signal_901), .Q (signal_12399) ) ;
    buf_clk cell_9869 ( .C (clk), .D (signal_4065), .Q (signal_12415) ) ;
    buf_clk cell_9885 ( .C (clk), .D (signal_904), .Q (signal_12431) ) ;
    buf_clk cell_9901 ( .C (clk), .D (signal_4066), .Q (signal_12447) ) ;
    buf_clk cell_9917 ( .C (clk), .D (signal_907), .Q (signal_12463) ) ;
    buf_clk cell_9933 ( .C (clk), .D (signal_4067), .Q (signal_12479) ) ;
    buf_clk cell_9949 ( .C (clk), .D (signal_910), .Q (signal_12495) ) ;
    buf_clk cell_9965 ( .C (clk), .D (signal_3675), .Q (signal_12511) ) ;
    buf_clk cell_9981 ( .C (clk), .D (signal_913), .Q (signal_12527) ) ;
    buf_clk cell_9997 ( .C (clk), .D (signal_3676), .Q (signal_12543) ) ;
    buf_clk cell_10013 ( .C (clk), .D (signal_916), .Q (signal_12559) ) ;
    buf_clk cell_10029 ( .C (clk), .D (signal_3677), .Q (signal_12575) ) ;
    buf_clk cell_10045 ( .C (clk), .D (signal_919), .Q (signal_12591) ) ;
    buf_clk cell_10061 ( .C (clk), .D (signal_3678), .Q (signal_12607) ) ;
    buf_clk cell_10077 ( .C (clk), .D (signal_922), .Q (signal_12623) ) ;
    buf_clk cell_10093 ( .C (clk), .D (signal_3679), .Q (signal_12639) ) ;
    buf_clk cell_10109 ( .C (clk), .D (signal_925), .Q (signal_12655) ) ;
    buf_clk cell_10125 ( .C (clk), .D (signal_3680), .Q (signal_12671) ) ;
    buf_clk cell_10141 ( .C (clk), .D (signal_928), .Q (signal_12687) ) ;
    buf_clk cell_10157 ( .C (clk), .D (signal_3681), .Q (signal_12703) ) ;
    buf_clk cell_10173 ( .C (clk), .D (signal_931), .Q (signal_12719) ) ;
    buf_clk cell_10189 ( .C (clk), .D (signal_3682), .Q (signal_12735) ) ;
    buf_clk cell_10205 ( .C (clk), .D (signal_934), .Q (signal_12751) ) ;
    buf_clk cell_10221 ( .C (clk), .D (signal_3683), .Q (signal_12767) ) ;
    buf_clk cell_10237 ( .C (clk), .D (signal_937), .Q (signal_12783) ) ;
    buf_clk cell_10253 ( .C (clk), .D (signal_3684), .Q (signal_12799) ) ;
    buf_clk cell_10269 ( .C (clk), .D (signal_940), .Q (signal_12815) ) ;
    buf_clk cell_10285 ( .C (clk), .D (signal_3685), .Q (signal_12831) ) ;
    buf_clk cell_10301 ( .C (clk), .D (signal_943), .Q (signal_12847) ) ;
    buf_clk cell_10317 ( .C (clk), .D (signal_3686), .Q (signal_12863) ) ;
    buf_clk cell_10333 ( .C (clk), .D (signal_946), .Q (signal_12879) ) ;
    buf_clk cell_10349 ( .C (clk), .D (signal_3687), .Q (signal_12895) ) ;
    buf_clk cell_10365 ( .C (clk), .D (signal_949), .Q (signal_12911) ) ;
    buf_clk cell_10381 ( .C (clk), .D (signal_3688), .Q (signal_12927) ) ;
    buf_clk cell_10397 ( .C (clk), .D (signal_952), .Q (signal_12943) ) ;
    buf_clk cell_10413 ( .C (clk), .D (signal_3689), .Q (signal_12959) ) ;
    buf_clk cell_10429 ( .C (clk), .D (signal_955), .Q (signal_12975) ) ;
    buf_clk cell_10445 ( .C (clk), .D (signal_3690), .Q (signal_12991) ) ;
    buf_clk cell_10461 ( .C (clk), .D (signal_958), .Q (signal_13007) ) ;
    buf_clk cell_10477 ( .C (clk), .D (signal_4068), .Q (signal_13023) ) ;
    buf_clk cell_10493 ( .C (clk), .D (signal_961), .Q (signal_13039) ) ;
    buf_clk cell_10509 ( .C (clk), .D (signal_4069), .Q (signal_13055) ) ;
    buf_clk cell_10525 ( .C (clk), .D (signal_964), .Q (signal_13071) ) ;
    buf_clk cell_10541 ( .C (clk), .D (signal_4070), .Q (signal_13087) ) ;
    buf_clk cell_10557 ( .C (clk), .D (signal_967), .Q (signal_13103) ) ;
    buf_clk cell_10573 ( .C (clk), .D (signal_4071), .Q (signal_13119) ) ;
    buf_clk cell_10589 ( .C (clk), .D (signal_970), .Q (signal_13135) ) ;
    buf_clk cell_10605 ( .C (clk), .D (signal_4072), .Q (signal_13151) ) ;
    buf_clk cell_10621 ( .C (clk), .D (signal_973), .Q (signal_13167) ) ;
    buf_clk cell_10637 ( .C (clk), .D (signal_4073), .Q (signal_13183) ) ;
    buf_clk cell_10653 ( .C (clk), .D (signal_976), .Q (signal_13199) ) ;
    buf_clk cell_10669 ( .C (clk), .D (signal_4074), .Q (signal_13215) ) ;
    buf_clk cell_10685 ( .C (clk), .D (signal_979), .Q (signal_13231) ) ;
    buf_clk cell_10701 ( .C (clk), .D (signal_4075), .Q (signal_13247) ) ;
    buf_clk cell_10717 ( .C (clk), .D (signal_982), .Q (signal_13263) ) ;
    buf_clk cell_10733 ( .C (clk), .D (signal_4076), .Q (signal_13279) ) ;
    buf_clk cell_10749 ( .C (clk), .D (signal_985), .Q (signal_13295) ) ;
    buf_clk cell_10765 ( .C (clk), .D (signal_4077), .Q (signal_13311) ) ;
    buf_clk cell_10781 ( .C (clk), .D (signal_988), .Q (signal_13327) ) ;
    buf_clk cell_10797 ( .C (clk), .D (signal_4078), .Q (signal_13343) ) ;
    buf_clk cell_10813 ( .C (clk), .D (signal_991), .Q (signal_13359) ) ;
    buf_clk cell_10829 ( .C (clk), .D (signal_4079), .Q (signal_13375) ) ;
    buf_clk cell_10845 ( .C (clk), .D (signal_994), .Q (signal_13391) ) ;
    buf_clk cell_10861 ( .C (clk), .D (signal_4080), .Q (signal_13407) ) ;
    buf_clk cell_10877 ( .C (clk), .D (signal_997), .Q (signal_13423) ) ;
    buf_clk cell_10893 ( .C (clk), .D (signal_4081), .Q (signal_13439) ) ;
    buf_clk cell_10909 ( .C (clk), .D (signal_1000), .Q (signal_13455) ) ;
    buf_clk cell_10925 ( .C (clk), .D (signal_4082), .Q (signal_13471) ) ;
    buf_clk cell_10941 ( .C (clk), .D (signal_1003), .Q (signal_13487) ) ;
    buf_clk cell_10957 ( .C (clk), .D (signal_4083), .Q (signal_13503) ) ;
    buf_clk cell_10973 ( .C (clk), .D (signal_1006), .Q (signal_13519) ) ;
    buf_clk cell_10989 ( .C (clk), .D (signal_4084), .Q (signal_13535) ) ;
    buf_clk cell_11005 ( .C (clk), .D (signal_1009), .Q (signal_13551) ) ;
    buf_clk cell_11021 ( .C (clk), .D (signal_4085), .Q (signal_13567) ) ;
    buf_clk cell_11037 ( .C (clk), .D (signal_1012), .Q (signal_13583) ) ;
    buf_clk cell_11053 ( .C (clk), .D (signal_4086), .Q (signal_13599) ) ;
    buf_clk cell_11069 ( .C (clk), .D (signal_1015), .Q (signal_13615) ) ;
    buf_clk cell_11085 ( .C (clk), .D (signal_4087), .Q (signal_13631) ) ;
    buf_clk cell_11101 ( .C (clk), .D (signal_1018), .Q (signal_13647) ) ;
    buf_clk cell_11117 ( .C (clk), .D (signal_4088), .Q (signal_13663) ) ;
    buf_clk cell_11133 ( .C (clk), .D (signal_1021), .Q (signal_13679) ) ;
    buf_clk cell_11149 ( .C (clk), .D (signal_4089), .Q (signal_13695) ) ;
    buf_clk cell_11165 ( .C (clk), .D (signal_1024), .Q (signal_13711) ) ;
    buf_clk cell_11181 ( .C (clk), .D (signal_4090), .Q (signal_13727) ) ;
    buf_clk cell_11197 ( .C (clk), .D (signal_1027), .Q (signal_13743) ) ;
    buf_clk cell_11213 ( .C (clk), .D (signal_4091), .Q (signal_13759) ) ;
    buf_clk cell_11229 ( .C (clk), .D (signal_1030), .Q (signal_13775) ) ;
    buf_clk cell_11245 ( .C (clk), .D (signal_4092), .Q (signal_13791) ) ;
    buf_clk cell_11261 ( .C (clk), .D (signal_1033), .Q (signal_13807) ) ;
    buf_clk cell_11277 ( .C (clk), .D (signal_4093), .Q (signal_13823) ) ;
    buf_clk cell_11293 ( .C (clk), .D (signal_1036), .Q (signal_13839) ) ;
    buf_clk cell_11309 ( .C (clk), .D (signal_4094), .Q (signal_13855) ) ;
    buf_clk cell_11325 ( .C (clk), .D (signal_1039), .Q (signal_13871) ) ;
    buf_clk cell_11341 ( .C (clk), .D (signal_4095), .Q (signal_13887) ) ;
    buf_clk cell_11357 ( .C (clk), .D (signal_1042), .Q (signal_13903) ) ;
    buf_clk cell_11373 ( .C (clk), .D (signal_4096), .Q (signal_13919) ) ;
    buf_clk cell_11389 ( .C (clk), .D (signal_1045), .Q (signal_13935) ) ;
    buf_clk cell_11405 ( .C (clk), .D (signal_4097), .Q (signal_13951) ) ;
    buf_clk cell_11421 ( .C (clk), .D (signal_1048), .Q (signal_13967) ) ;
    buf_clk cell_11437 ( .C (clk), .D (signal_4098), .Q (signal_13983) ) ;
    buf_clk cell_11453 ( .C (clk), .D (signal_1051), .Q (signal_13999) ) ;
    buf_clk cell_11469 ( .C (clk), .D (signal_4099), .Q (signal_14015) ) ;
    buf_clk cell_11485 ( .C (clk), .D (signal_1078), .Q (signal_14031) ) ;
    buf_clk cell_11501 ( .C (clk), .D (signal_4100), .Q (signal_14047) ) ;
    buf_clk cell_11517 ( .C (clk), .D (signal_1081), .Q (signal_14063) ) ;
    buf_clk cell_11533 ( .C (clk), .D (signal_4101), .Q (signal_14079) ) ;
    buf_clk cell_11549 ( .C (clk), .D (signal_1084), .Q (signal_14095) ) ;
    buf_clk cell_11565 ( .C (clk), .D (signal_4102), .Q (signal_14111) ) ;
    buf_clk cell_11581 ( .C (clk), .D (signal_1087), .Q (signal_14127) ) ;
    buf_clk cell_11597 ( .C (clk), .D (signal_4103), .Q (signal_14143) ) ;
    buf_clk cell_11613 ( .C (clk), .D (signal_1090), .Q (signal_14159) ) ;
    buf_clk cell_11629 ( .C (clk), .D (signal_4104), .Q (signal_14175) ) ;
    buf_clk cell_11645 ( .C (clk), .D (signal_1093), .Q (signal_14191) ) ;
    buf_clk cell_11661 ( .C (clk), .D (signal_4105), .Q (signal_14207) ) ;
    buf_clk cell_11677 ( .C (clk), .D (signal_1096), .Q (signal_14223) ) ;
    buf_clk cell_11693 ( .C (clk), .D (signal_4106), .Q (signal_14239) ) ;
    buf_clk cell_11709 ( .C (clk), .D (signal_1099), .Q (signal_14255) ) ;
    buf_clk cell_11725 ( .C (clk), .D (signal_4107), .Q (signal_14271) ) ;
    buf_clk cell_11741 ( .C (clk), .D (signal_1102), .Q (signal_14287) ) ;
    buf_clk cell_11757 ( .C (clk), .D (signal_4108), .Q (signal_14303) ) ;
    buf_clk cell_11773 ( .C (clk), .D (signal_1105), .Q (signal_14319) ) ;
    buf_clk cell_11789 ( .C (clk), .D (signal_4109), .Q (signal_14335) ) ;
    buf_clk cell_11805 ( .C (clk), .D (signal_1108), .Q (signal_14351) ) ;
    buf_clk cell_11821 ( .C (clk), .D (signal_4110), .Q (signal_14367) ) ;
    buf_clk cell_11837 ( .C (clk), .D (signal_1111), .Q (signal_14383) ) ;
    buf_clk cell_11853 ( .C (clk), .D (signal_4111), .Q (signal_14399) ) ;
    buf_clk cell_11869 ( .C (clk), .D (signal_1114), .Q (signal_14415) ) ;
    buf_clk cell_11885 ( .C (clk), .D (signal_4112), .Q (signal_14431) ) ;
    buf_clk cell_11901 ( .C (clk), .D (signal_1117), .Q (signal_14447) ) ;
    buf_clk cell_11917 ( .C (clk), .D (signal_4113), .Q (signal_14463) ) ;
    buf_clk cell_11933 ( .C (clk), .D (signal_1120), .Q (signal_14479) ) ;
    buf_clk cell_11949 ( .C (clk), .D (signal_4114), .Q (signal_14495) ) ;
    buf_clk cell_11965 ( .C (clk), .D (signal_1123), .Q (signal_14511) ) ;
    buf_clk cell_11981 ( .C (clk), .D (signal_4115), .Q (signal_14527) ) ;
    buf_clk cell_11997 ( .C (clk), .D (signal_1126), .Q (signal_14543) ) ;
    buf_clk cell_12013 ( .C (clk), .D (signal_4116), .Q (signal_14559) ) ;
    buf_clk cell_12029 ( .C (clk), .D (signal_1129), .Q (signal_14575) ) ;
    buf_clk cell_12045 ( .C (clk), .D (signal_4117), .Q (signal_14591) ) ;
    buf_clk cell_12061 ( .C (clk), .D (signal_1132), .Q (signal_14607) ) ;
    buf_clk cell_12077 ( .C (clk), .D (signal_4118), .Q (signal_14623) ) ;
    buf_clk cell_12093 ( .C (clk), .D (signal_1135), .Q (signal_14639) ) ;
    buf_clk cell_12109 ( .C (clk), .D (signal_4119), .Q (signal_14655) ) ;
    buf_clk cell_12125 ( .C (clk), .D (signal_1138), .Q (signal_14671) ) ;
    buf_clk cell_12141 ( .C (clk), .D (signal_4120), .Q (signal_14687) ) ;
    buf_clk cell_12157 ( .C (clk), .D (signal_1141), .Q (signal_14703) ) ;
    buf_clk cell_12173 ( .C (clk), .D (signal_4121), .Q (signal_14719) ) ;
    buf_clk cell_12189 ( .C (clk), .D (signal_1144), .Q (signal_14735) ) ;
    buf_clk cell_12205 ( .C (clk), .D (signal_4122), .Q (signal_14751) ) ;
    buf_clk cell_12221 ( .C (clk), .D (signal_1147), .Q (signal_14767) ) ;
    buf_clk cell_12237 ( .C (clk), .D (signal_4123), .Q (signal_14783) ) ;
    buf_clk cell_12253 ( .C (clk), .D (signal_1275), .Q (signal_14799) ) ;
    buf_clk cell_12269 ( .C (clk), .D (signal_1266), .Q (signal_14815) ) ;
    buf_clk cell_12285 ( .C (clk), .D (signal_1264), .Q (signal_14831) ) ;
    buf_clk cell_12301 ( .C (clk), .D (signal_1262), .Q (signal_14847) ) ;
    buf_clk cell_12317 ( .C (clk), .D (signal_1260), .Q (signal_14863) ) ;
    buf_clk cell_12333 ( .C (clk), .D (signal_1259), .Q (signal_14879) ) ;
    buf_clk cell_12349 ( .C (clk), .D (signal_1258), .Q (signal_14895) ) ;
    buf_clk cell_12365 ( .C (clk), .D (signal_1256), .Q (signal_14911) ) ;
    buf_clk cell_12381 ( .C (clk), .D (signal_403), .Q (signal_14927) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1714 ( .s ({signal_3256, signal_1510}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[0]), .c ({signal_3273, signal_1982}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1715 ( .s ({signal_3256, signal_1510}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[1]), .c ({signal_3274, signal_1983}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1716 ( .s ({signal_3255, signal_1511}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_3275, signal_1984}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1717 ( .s ({signal_3255, signal_1511}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[3]), .c ({signal_3276, signal_1985}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1718 ( .s ({signal_3254, signal_1512}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[4]), .c ({signal_3277, signal_1986}) ) ;
    buf_clk cell_2146 ( .C (clk), .D (signal_4691), .Q (signal_4692) ) ;
    buf_clk cell_2148 ( .C (clk), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_2150 ( .C (clk), .D (signal_4695), .Q (signal_4696) ) ;
    buf_clk cell_2152 ( .C (clk), .D (signal_4697), .Q (signal_4698) ) ;
    buf_clk cell_2170 ( .C (clk), .D (signal_4715), .Q (signal_4716) ) ;
    buf_clk cell_2174 ( .C (clk), .D (signal_4719), .Q (signal_4720) ) ;
    buf_clk cell_2298 ( .C (clk), .D (signal_4843), .Q (signal_4844) ) ;
    buf_clk cell_2306 ( .C (clk), .D (signal_4851), .Q (signal_4852) ) ;
    buf_clk cell_2342 ( .C (clk), .D (signal_4887), .Q (signal_4888) ) ;
    buf_clk cell_2352 ( .C (clk), .D (signal_4897), .Q (signal_4898) ) ;
    buf_clk cell_2362 ( .C (clk), .D (signal_4907), .Q (signal_4908) ) ;
    buf_clk cell_2374 ( .C (clk), .D (signal_4919), .Q (signal_4920) ) ;
    buf_clk cell_2386 ( .C (clk), .D (signal_4931), .Q (signal_4932) ) ;
    buf_clk cell_2402 ( .C (clk), .D (signal_4947), .Q (signal_4948) ) ;
    buf_clk cell_2418 ( .C (clk), .D (signal_4963), .Q (signal_4964) ) ;
    buf_clk cell_2434 ( .C (clk), .D (signal_4979), .Q (signal_4980) ) ;
    buf_clk cell_2450 ( .C (clk), .D (signal_4995), .Q (signal_4996) ) ;
    buf_clk cell_2466 ( .C (clk), .D (signal_5011), .Q (signal_5012) ) ;
    buf_clk cell_2482 ( .C (clk), .D (signal_5027), .Q (signal_5028) ) ;
    buf_clk cell_2498 ( .C (clk), .D (signal_5043), .Q (signal_5044) ) ;
    buf_clk cell_2514 ( .C (clk), .D (signal_5059), .Q (signal_5060) ) ;
    buf_clk cell_2530 ( .C (clk), .D (signal_5075), .Q (signal_5076) ) ;
    buf_clk cell_2546 ( .C (clk), .D (signal_5091), .Q (signal_5092) ) ;
    buf_clk cell_2562 ( .C (clk), .D (signal_5107), .Q (signal_5108) ) ;
    buf_clk cell_2578 ( .C (clk), .D (signal_5123), .Q (signal_5124) ) ;
    buf_clk cell_2594 ( .C (clk), .D (signal_5139), .Q (signal_5140) ) ;
    buf_clk cell_2610 ( .C (clk), .D (signal_5155), .Q (signal_5156) ) ;
    buf_clk cell_2626 ( .C (clk), .D (signal_5171), .Q (signal_5172) ) ;
    buf_clk cell_2642 ( .C (clk), .D (signal_5187), .Q (signal_5188) ) ;
    buf_clk cell_2658 ( .C (clk), .D (signal_5203), .Q (signal_5204) ) ;
    buf_clk cell_2674 ( .C (clk), .D (signal_5219), .Q (signal_5220) ) ;
    buf_clk cell_2690 ( .C (clk), .D (signal_5235), .Q (signal_5236) ) ;
    buf_clk cell_2706 ( .C (clk), .D (signal_5251), .Q (signal_5252) ) ;
    buf_clk cell_2722 ( .C (clk), .D (signal_5267), .Q (signal_5268) ) ;
    buf_clk cell_2738 ( .C (clk), .D (signal_5283), .Q (signal_5284) ) ;
    buf_clk cell_2754 ( .C (clk), .D (signal_5299), .Q (signal_5300) ) ;
    buf_clk cell_2770 ( .C (clk), .D (signal_5315), .Q (signal_5316) ) ;
    buf_clk cell_2786 ( .C (clk), .D (signal_5331), .Q (signal_5332) ) ;
    buf_clk cell_2802 ( .C (clk), .D (signal_5347), .Q (signal_5348) ) ;
    buf_clk cell_2818 ( .C (clk), .D (signal_5363), .Q (signal_5364) ) ;
    buf_clk cell_2834 ( .C (clk), .D (signal_5379), .Q (signal_5380) ) ;
    buf_clk cell_2850 ( .C (clk), .D (signal_5395), .Q (signal_5396) ) ;
    buf_clk cell_2866 ( .C (clk), .D (signal_5411), .Q (signal_5412) ) ;
    buf_clk cell_2882 ( .C (clk), .D (signal_5427), .Q (signal_5428) ) ;
    buf_clk cell_2898 ( .C (clk), .D (signal_5443), .Q (signal_5444) ) ;
    buf_clk cell_2914 ( .C (clk), .D (signal_5459), .Q (signal_5460) ) ;
    buf_clk cell_2930 ( .C (clk), .D (signal_5475), .Q (signal_5476) ) ;
    buf_clk cell_2946 ( .C (clk), .D (signal_5491), .Q (signal_5492) ) ;
    buf_clk cell_2962 ( .C (clk), .D (signal_5507), .Q (signal_5508) ) ;
    buf_clk cell_2978 ( .C (clk), .D (signal_5523), .Q (signal_5524) ) ;
    buf_clk cell_2994 ( .C (clk), .D (signal_5539), .Q (signal_5540) ) ;
    buf_clk cell_3010 ( .C (clk), .D (signal_5555), .Q (signal_5556) ) ;
    buf_clk cell_3026 ( .C (clk), .D (signal_5571), .Q (signal_5572) ) ;
    buf_clk cell_3042 ( .C (clk), .D (signal_5587), .Q (signal_5588) ) ;
    buf_clk cell_3058 ( .C (clk), .D (signal_5603), .Q (signal_5604) ) ;
    buf_clk cell_3074 ( .C (clk), .D (signal_5619), .Q (signal_5620) ) ;
    buf_clk cell_3090 ( .C (clk), .D (signal_5635), .Q (signal_5636) ) ;
    buf_clk cell_3106 ( .C (clk), .D (signal_5651), .Q (signal_5652) ) ;
    buf_clk cell_3122 ( .C (clk), .D (signal_5667), .Q (signal_5668) ) ;
    buf_clk cell_3138 ( .C (clk), .D (signal_5683), .Q (signal_5684) ) ;
    buf_clk cell_3154 ( .C (clk), .D (signal_5699), .Q (signal_5700) ) ;
    buf_clk cell_3170 ( .C (clk), .D (signal_5715), .Q (signal_5716) ) ;
    buf_clk cell_3186 ( .C (clk), .D (signal_5731), .Q (signal_5732) ) ;
    buf_clk cell_3202 ( .C (clk), .D (signal_5747), .Q (signal_5748) ) ;
    buf_clk cell_3218 ( .C (clk), .D (signal_5763), .Q (signal_5764) ) ;
    buf_clk cell_3234 ( .C (clk), .D (signal_5779), .Q (signal_5780) ) ;
    buf_clk cell_3250 ( .C (clk), .D (signal_5795), .Q (signal_5796) ) ;
    buf_clk cell_3266 ( .C (clk), .D (signal_5811), .Q (signal_5812) ) ;
    buf_clk cell_3282 ( .C (clk), .D (signal_5827), .Q (signal_5828) ) ;
    buf_clk cell_3298 ( .C (clk), .D (signal_5843), .Q (signal_5844) ) ;
    buf_clk cell_3314 ( .C (clk), .D (signal_5859), .Q (signal_5860) ) ;
    buf_clk cell_3330 ( .C (clk), .D (signal_5875), .Q (signal_5876) ) ;
    buf_clk cell_3346 ( .C (clk), .D (signal_5891), .Q (signal_5892) ) ;
    buf_clk cell_3362 ( .C (clk), .D (signal_5907), .Q (signal_5908) ) ;
    buf_clk cell_3378 ( .C (clk), .D (signal_5923), .Q (signal_5924) ) ;
    buf_clk cell_3394 ( .C (clk), .D (signal_5939), .Q (signal_5940) ) ;
    buf_clk cell_3410 ( .C (clk), .D (signal_5955), .Q (signal_5956) ) ;
    buf_clk cell_3426 ( .C (clk), .D (signal_5971), .Q (signal_5972) ) ;
    buf_clk cell_3442 ( .C (clk), .D (signal_5987), .Q (signal_5988) ) ;
    buf_clk cell_3458 ( .C (clk), .D (signal_6003), .Q (signal_6004) ) ;
    buf_clk cell_3474 ( .C (clk), .D (signal_6019), .Q (signal_6020) ) ;
    buf_clk cell_3490 ( .C (clk), .D (signal_6035), .Q (signal_6036) ) ;
    buf_clk cell_3506 ( .C (clk), .D (signal_6051), .Q (signal_6052) ) ;
    buf_clk cell_3522 ( .C (clk), .D (signal_6067), .Q (signal_6068) ) ;
    buf_clk cell_3538 ( .C (clk), .D (signal_6083), .Q (signal_6084) ) ;
    buf_clk cell_3554 ( .C (clk), .D (signal_6099), .Q (signal_6100) ) ;
    buf_clk cell_3570 ( .C (clk), .D (signal_6115), .Q (signal_6116) ) ;
    buf_clk cell_3586 ( .C (clk), .D (signal_6131), .Q (signal_6132) ) ;
    buf_clk cell_3602 ( .C (clk), .D (signal_6147), .Q (signal_6148) ) ;
    buf_clk cell_3618 ( .C (clk), .D (signal_6163), .Q (signal_6164) ) ;
    buf_clk cell_3634 ( .C (clk), .D (signal_6179), .Q (signal_6180) ) ;
    buf_clk cell_3650 ( .C (clk), .D (signal_6195), .Q (signal_6196) ) ;
    buf_clk cell_3666 ( .C (clk), .D (signal_6211), .Q (signal_6212) ) ;
    buf_clk cell_3682 ( .C (clk), .D (signal_6227), .Q (signal_6228) ) ;
    buf_clk cell_3698 ( .C (clk), .D (signal_6243), .Q (signal_6244) ) ;
    buf_clk cell_3714 ( .C (clk), .D (signal_6259), .Q (signal_6260) ) ;
    buf_clk cell_3730 ( .C (clk), .D (signal_6275), .Q (signal_6276) ) ;
    buf_clk cell_3746 ( .C (clk), .D (signal_6291), .Q (signal_6292) ) ;
    buf_clk cell_3762 ( .C (clk), .D (signal_6307), .Q (signal_6308) ) ;
    buf_clk cell_3778 ( .C (clk), .D (signal_6323), .Q (signal_6324) ) ;
    buf_clk cell_3794 ( .C (clk), .D (signal_6339), .Q (signal_6340) ) ;
    buf_clk cell_3810 ( .C (clk), .D (signal_6355), .Q (signal_6356) ) ;
    buf_clk cell_3826 ( .C (clk), .D (signal_6371), .Q (signal_6372) ) ;
    buf_clk cell_3842 ( .C (clk), .D (signal_6387), .Q (signal_6388) ) ;
    buf_clk cell_3858 ( .C (clk), .D (signal_6403), .Q (signal_6404) ) ;
    buf_clk cell_3874 ( .C (clk), .D (signal_6419), .Q (signal_6420) ) ;
    buf_clk cell_3890 ( .C (clk), .D (signal_6435), .Q (signal_6436) ) ;
    buf_clk cell_3906 ( .C (clk), .D (signal_6451), .Q (signal_6452) ) ;
    buf_clk cell_3922 ( .C (clk), .D (signal_6467), .Q (signal_6468) ) ;
    buf_clk cell_3938 ( .C (clk), .D (signal_6483), .Q (signal_6484) ) ;
    buf_clk cell_3954 ( .C (clk), .D (signal_6499), .Q (signal_6500) ) ;
    buf_clk cell_3970 ( .C (clk), .D (signal_6515), .Q (signal_6516) ) ;
    buf_clk cell_3986 ( .C (clk), .D (signal_6531), .Q (signal_6532) ) ;
    buf_clk cell_4002 ( .C (clk), .D (signal_6547), .Q (signal_6548) ) ;
    buf_clk cell_4018 ( .C (clk), .D (signal_6563), .Q (signal_6564) ) ;
    buf_clk cell_4034 ( .C (clk), .D (signal_6579), .Q (signal_6580) ) ;
    buf_clk cell_4050 ( .C (clk), .D (signal_6595), .Q (signal_6596) ) ;
    buf_clk cell_4066 ( .C (clk), .D (signal_6611), .Q (signal_6612) ) ;
    buf_clk cell_4082 ( .C (clk), .D (signal_6627), .Q (signal_6628) ) ;
    buf_clk cell_4098 ( .C (clk), .D (signal_6643), .Q (signal_6644) ) ;
    buf_clk cell_4114 ( .C (clk), .D (signal_6659), .Q (signal_6660) ) ;
    buf_clk cell_4130 ( .C (clk), .D (signal_6675), .Q (signal_6676) ) ;
    buf_clk cell_4146 ( .C (clk), .D (signal_6691), .Q (signal_6692) ) ;
    buf_clk cell_4162 ( .C (clk), .D (signal_6707), .Q (signal_6708) ) ;
    buf_clk cell_4178 ( .C (clk), .D (signal_6723), .Q (signal_6724) ) ;
    buf_clk cell_4194 ( .C (clk), .D (signal_6739), .Q (signal_6740) ) ;
    buf_clk cell_4210 ( .C (clk), .D (signal_6755), .Q (signal_6756) ) ;
    buf_clk cell_4226 ( .C (clk), .D (signal_6771), .Q (signal_6772) ) ;
    buf_clk cell_4242 ( .C (clk), .D (signal_6787), .Q (signal_6788) ) ;
    buf_clk cell_4258 ( .C (clk), .D (signal_6803), .Q (signal_6804) ) ;
    buf_clk cell_4274 ( .C (clk), .D (signal_6819), .Q (signal_6820) ) ;
    buf_clk cell_4290 ( .C (clk), .D (signal_6835), .Q (signal_6836) ) ;
    buf_clk cell_4306 ( .C (clk), .D (signal_6851), .Q (signal_6852) ) ;
    buf_clk cell_4322 ( .C (clk), .D (signal_6867), .Q (signal_6868) ) ;
    buf_clk cell_4338 ( .C (clk), .D (signal_6883), .Q (signal_6884) ) ;
    buf_clk cell_4354 ( .C (clk), .D (signal_6899), .Q (signal_6900) ) ;
    buf_clk cell_4370 ( .C (clk), .D (signal_6915), .Q (signal_6916) ) ;
    buf_clk cell_4386 ( .C (clk), .D (signal_6931), .Q (signal_6932) ) ;
    buf_clk cell_4402 ( .C (clk), .D (signal_6947), .Q (signal_6948) ) ;
    buf_clk cell_4416 ( .C (clk), .D (signal_6961), .Q (signal_6962) ) ;
    buf_clk cell_4430 ( .C (clk), .D (signal_6975), .Q (signal_6976) ) ;
    buf_clk cell_4446 ( .C (clk), .D (signal_6991), .Q (signal_6992) ) ;
    buf_clk cell_4462 ( .C (clk), .D (signal_7007), .Q (signal_7008) ) ;
    buf_clk cell_4478 ( .C (clk), .D (signal_7023), .Q (signal_7024) ) ;
    buf_clk cell_4494 ( .C (clk), .D (signal_7039), .Q (signal_7040) ) ;
    buf_clk cell_4510 ( .C (clk), .D (signal_7055), .Q (signal_7056) ) ;
    buf_clk cell_4526 ( .C (clk), .D (signal_7071), .Q (signal_7072) ) ;
    buf_clk cell_4542 ( .C (clk), .D (signal_7087), .Q (signal_7088) ) ;
    buf_clk cell_4558 ( .C (clk), .D (signal_7103), .Q (signal_7104) ) ;
    buf_clk cell_4574 ( .C (clk), .D (signal_7119), .Q (signal_7120) ) ;
    buf_clk cell_4590 ( .C (clk), .D (signal_7135), .Q (signal_7136) ) ;
    buf_clk cell_4606 ( .C (clk), .D (signal_7151), .Q (signal_7152) ) ;
    buf_clk cell_4622 ( .C (clk), .D (signal_7167), .Q (signal_7168) ) ;
    buf_clk cell_4638 ( .C (clk), .D (signal_7183), .Q (signal_7184) ) ;
    buf_clk cell_4654 ( .C (clk), .D (signal_7199), .Q (signal_7200) ) ;
    buf_clk cell_4670 ( .C (clk), .D (signal_7215), .Q (signal_7216) ) ;
    buf_clk cell_4686 ( .C (clk), .D (signal_7231), .Q (signal_7232) ) ;
    buf_clk cell_4702 ( .C (clk), .D (signal_7247), .Q (signal_7248) ) ;
    buf_clk cell_4718 ( .C (clk), .D (signal_7263), .Q (signal_7264) ) ;
    buf_clk cell_4734 ( .C (clk), .D (signal_7279), .Q (signal_7280) ) ;
    buf_clk cell_4750 ( .C (clk), .D (signal_7295), .Q (signal_7296) ) ;
    buf_clk cell_4766 ( .C (clk), .D (signal_7311), .Q (signal_7312) ) ;
    buf_clk cell_4782 ( .C (clk), .D (signal_7327), .Q (signal_7328) ) ;
    buf_clk cell_4798 ( .C (clk), .D (signal_7343), .Q (signal_7344) ) ;
    buf_clk cell_4814 ( .C (clk), .D (signal_7359), .Q (signal_7360) ) ;
    buf_clk cell_4830 ( .C (clk), .D (signal_7375), .Q (signal_7376) ) ;
    buf_clk cell_4846 ( .C (clk), .D (signal_7391), .Q (signal_7392) ) ;
    buf_clk cell_4862 ( .C (clk), .D (signal_7407), .Q (signal_7408) ) ;
    buf_clk cell_4878 ( .C (clk), .D (signal_7423), .Q (signal_7424) ) ;
    buf_clk cell_4894 ( .C (clk), .D (signal_7439), .Q (signal_7440) ) ;
    buf_clk cell_4910 ( .C (clk), .D (signal_7455), .Q (signal_7456) ) ;
    buf_clk cell_4926 ( .C (clk), .D (signal_7471), .Q (signal_7472) ) ;
    buf_clk cell_4942 ( .C (clk), .D (signal_7487), .Q (signal_7488) ) ;
    buf_clk cell_4958 ( .C (clk), .D (signal_7503), .Q (signal_7504) ) ;
    buf_clk cell_4974 ( .C (clk), .D (signal_7519), .Q (signal_7520) ) ;
    buf_clk cell_4990 ( .C (clk), .D (signal_7535), .Q (signal_7536) ) ;
    buf_clk cell_5006 ( .C (clk), .D (signal_7551), .Q (signal_7552) ) ;
    buf_clk cell_5022 ( .C (clk), .D (signal_7567), .Q (signal_7568) ) ;
    buf_clk cell_5038 ( .C (clk), .D (signal_7583), .Q (signal_7584) ) ;
    buf_clk cell_5054 ( .C (clk), .D (signal_7599), .Q (signal_7600) ) ;
    buf_clk cell_5070 ( .C (clk), .D (signal_7615), .Q (signal_7616) ) ;
    buf_clk cell_5086 ( .C (clk), .D (signal_7631), .Q (signal_7632) ) ;
    buf_clk cell_5102 ( .C (clk), .D (signal_7647), .Q (signal_7648) ) ;
    buf_clk cell_5118 ( .C (clk), .D (signal_7663), .Q (signal_7664) ) ;
    buf_clk cell_5134 ( .C (clk), .D (signal_7679), .Q (signal_7680) ) ;
    buf_clk cell_5150 ( .C (clk), .D (signal_7695), .Q (signal_7696) ) ;
    buf_clk cell_5166 ( .C (clk), .D (signal_7711), .Q (signal_7712) ) ;
    buf_clk cell_5182 ( .C (clk), .D (signal_7727), .Q (signal_7728) ) ;
    buf_clk cell_5198 ( .C (clk), .D (signal_7743), .Q (signal_7744) ) ;
    buf_clk cell_5214 ( .C (clk), .D (signal_7759), .Q (signal_7760) ) ;
    buf_clk cell_5230 ( .C (clk), .D (signal_7775), .Q (signal_7776) ) ;
    buf_clk cell_5246 ( .C (clk), .D (signal_7791), .Q (signal_7792) ) ;
    buf_clk cell_5262 ( .C (clk), .D (signal_7807), .Q (signal_7808) ) ;
    buf_clk cell_5278 ( .C (clk), .D (signal_7823), .Q (signal_7824) ) ;
    buf_clk cell_5294 ( .C (clk), .D (signal_7839), .Q (signal_7840) ) ;
    buf_clk cell_5310 ( .C (clk), .D (signal_7855), .Q (signal_7856) ) ;
    buf_clk cell_5326 ( .C (clk), .D (signal_7871), .Q (signal_7872) ) ;
    buf_clk cell_5342 ( .C (clk), .D (signal_7887), .Q (signal_7888) ) ;
    buf_clk cell_5358 ( .C (clk), .D (signal_7903), .Q (signal_7904) ) ;
    buf_clk cell_5374 ( .C (clk), .D (signal_7919), .Q (signal_7920) ) ;
    buf_clk cell_5390 ( .C (clk), .D (signal_7935), .Q (signal_7936) ) ;
    buf_clk cell_5406 ( .C (clk), .D (signal_7951), .Q (signal_7952) ) ;
    buf_clk cell_5422 ( .C (clk), .D (signal_7967), .Q (signal_7968) ) ;
    buf_clk cell_5438 ( .C (clk), .D (signal_7983), .Q (signal_7984) ) ;
    buf_clk cell_5454 ( .C (clk), .D (signal_7999), .Q (signal_8000) ) ;
    buf_clk cell_5470 ( .C (clk), .D (signal_8015), .Q (signal_8016) ) ;
    buf_clk cell_5486 ( .C (clk), .D (signal_8031), .Q (signal_8032) ) ;
    buf_clk cell_5502 ( .C (clk), .D (signal_8047), .Q (signal_8048) ) ;
    buf_clk cell_5518 ( .C (clk), .D (signal_8063), .Q (signal_8064) ) ;
    buf_clk cell_5534 ( .C (clk), .D (signal_8079), .Q (signal_8080) ) ;
    buf_clk cell_5550 ( .C (clk), .D (signal_8095), .Q (signal_8096) ) ;
    buf_clk cell_5566 ( .C (clk), .D (signal_8111), .Q (signal_8112) ) ;
    buf_clk cell_5582 ( .C (clk), .D (signal_8127), .Q (signal_8128) ) ;
    buf_clk cell_5598 ( .C (clk), .D (signal_8143), .Q (signal_8144) ) ;
    buf_clk cell_5614 ( .C (clk), .D (signal_8159), .Q (signal_8160) ) ;
    buf_clk cell_5630 ( .C (clk), .D (signal_8175), .Q (signal_8176) ) ;
    buf_clk cell_5646 ( .C (clk), .D (signal_8191), .Q (signal_8192) ) ;
    buf_clk cell_5662 ( .C (clk), .D (signal_8207), .Q (signal_8208) ) ;
    buf_clk cell_5678 ( .C (clk), .D (signal_8223), .Q (signal_8224) ) ;
    buf_clk cell_5694 ( .C (clk), .D (signal_8239), .Q (signal_8240) ) ;
    buf_clk cell_5710 ( .C (clk), .D (signal_8255), .Q (signal_8256) ) ;
    buf_clk cell_5726 ( .C (clk), .D (signal_8271), .Q (signal_8272) ) ;
    buf_clk cell_5742 ( .C (clk), .D (signal_8287), .Q (signal_8288) ) ;
    buf_clk cell_5758 ( .C (clk), .D (signal_8303), .Q (signal_8304) ) ;
    buf_clk cell_5774 ( .C (clk), .D (signal_8319), .Q (signal_8320) ) ;
    buf_clk cell_5790 ( .C (clk), .D (signal_8335), .Q (signal_8336) ) ;
    buf_clk cell_5806 ( .C (clk), .D (signal_8351), .Q (signal_8352) ) ;
    buf_clk cell_5822 ( .C (clk), .D (signal_8367), .Q (signal_8368) ) ;
    buf_clk cell_5838 ( .C (clk), .D (signal_8383), .Q (signal_8384) ) ;
    buf_clk cell_5854 ( .C (clk), .D (signal_8399), .Q (signal_8400) ) ;
    buf_clk cell_5870 ( .C (clk), .D (signal_8415), .Q (signal_8416) ) ;
    buf_clk cell_5886 ( .C (clk), .D (signal_8431), .Q (signal_8432) ) ;
    buf_clk cell_5902 ( .C (clk), .D (signal_8447), .Q (signal_8448) ) ;
    buf_clk cell_5918 ( .C (clk), .D (signal_8463), .Q (signal_8464) ) ;
    buf_clk cell_5934 ( .C (clk), .D (signal_8479), .Q (signal_8480) ) ;
    buf_clk cell_5950 ( .C (clk), .D (signal_8495), .Q (signal_8496) ) ;
    buf_clk cell_5966 ( .C (clk), .D (signal_8511), .Q (signal_8512) ) ;
    buf_clk cell_5982 ( .C (clk), .D (signal_8527), .Q (signal_8528) ) ;
    buf_clk cell_5998 ( .C (clk), .D (signal_8543), .Q (signal_8544) ) ;
    buf_clk cell_6014 ( .C (clk), .D (signal_8559), .Q (signal_8560) ) ;
    buf_clk cell_6030 ( .C (clk), .D (signal_8575), .Q (signal_8576) ) ;
    buf_clk cell_6046 ( .C (clk), .D (signal_8591), .Q (signal_8592) ) ;
    buf_clk cell_6062 ( .C (clk), .D (signal_8607), .Q (signal_8608) ) ;
    buf_clk cell_6078 ( .C (clk), .D (signal_8623), .Q (signal_8624) ) ;
    buf_clk cell_6094 ( .C (clk), .D (signal_8639), .Q (signal_8640) ) ;
    buf_clk cell_6110 ( .C (clk), .D (signal_8655), .Q (signal_8656) ) ;
    buf_clk cell_6126 ( .C (clk), .D (signal_8671), .Q (signal_8672) ) ;
    buf_clk cell_6142 ( .C (clk), .D (signal_8687), .Q (signal_8688) ) ;
    buf_clk cell_6158 ( .C (clk), .D (signal_8703), .Q (signal_8704) ) ;
    buf_clk cell_6174 ( .C (clk), .D (signal_8719), .Q (signal_8720) ) ;
    buf_clk cell_6190 ( .C (clk), .D (signal_8735), .Q (signal_8736) ) ;
    buf_clk cell_6206 ( .C (clk), .D (signal_8751), .Q (signal_8752) ) ;
    buf_clk cell_6222 ( .C (clk), .D (signal_8767), .Q (signal_8768) ) ;
    buf_clk cell_6238 ( .C (clk), .D (signal_8783), .Q (signal_8784) ) ;
    buf_clk cell_6254 ( .C (clk), .D (signal_8799), .Q (signal_8800) ) ;
    buf_clk cell_6270 ( .C (clk), .D (signal_8815), .Q (signal_8816) ) ;
    buf_clk cell_6286 ( .C (clk), .D (signal_8831), .Q (signal_8832) ) ;
    buf_clk cell_6302 ( .C (clk), .D (signal_8847), .Q (signal_8848) ) ;
    buf_clk cell_6318 ( .C (clk), .D (signal_8863), .Q (signal_8864) ) ;
    buf_clk cell_6334 ( .C (clk), .D (signal_8879), .Q (signal_8880) ) ;
    buf_clk cell_6350 ( .C (clk), .D (signal_8895), .Q (signal_8896) ) ;
    buf_clk cell_6366 ( .C (clk), .D (signal_8911), .Q (signal_8912) ) ;
    buf_clk cell_6382 ( .C (clk), .D (signal_8927), .Q (signal_8928) ) ;
    buf_clk cell_6398 ( .C (clk), .D (signal_8943), .Q (signal_8944) ) ;
    buf_clk cell_6414 ( .C (clk), .D (signal_8959), .Q (signal_8960) ) ;
    buf_clk cell_6430 ( .C (clk), .D (signal_8975), .Q (signal_8976) ) ;
    buf_clk cell_6446 ( .C (clk), .D (signal_8991), .Q (signal_8992) ) ;
    buf_clk cell_6462 ( .C (clk), .D (signal_9007), .Q (signal_9008) ) ;
    buf_clk cell_6478 ( .C (clk), .D (signal_9023), .Q (signal_9024) ) ;
    buf_clk cell_6494 ( .C (clk), .D (signal_9039), .Q (signal_9040) ) ;
    buf_clk cell_6510 ( .C (clk), .D (signal_9055), .Q (signal_9056) ) ;
    buf_clk cell_6526 ( .C (clk), .D (signal_9071), .Q (signal_9072) ) ;
    buf_clk cell_6542 ( .C (clk), .D (signal_9087), .Q (signal_9088) ) ;
    buf_clk cell_6558 ( .C (clk), .D (signal_9103), .Q (signal_9104) ) ;
    buf_clk cell_6574 ( .C (clk), .D (signal_9119), .Q (signal_9120) ) ;
    buf_clk cell_6590 ( .C (clk), .D (signal_9135), .Q (signal_9136) ) ;
    buf_clk cell_6606 ( .C (clk), .D (signal_9151), .Q (signal_9152) ) ;
    buf_clk cell_6622 ( .C (clk), .D (signal_9167), .Q (signal_9168) ) ;
    buf_clk cell_6638 ( .C (clk), .D (signal_9183), .Q (signal_9184) ) ;
    buf_clk cell_6654 ( .C (clk), .D (signal_9199), .Q (signal_9200) ) ;
    buf_clk cell_6670 ( .C (clk), .D (signal_9215), .Q (signal_9216) ) ;
    buf_clk cell_6686 ( .C (clk), .D (signal_9231), .Q (signal_9232) ) ;
    buf_clk cell_6702 ( .C (clk), .D (signal_9247), .Q (signal_9248) ) ;
    buf_clk cell_6718 ( .C (clk), .D (signal_9263), .Q (signal_9264) ) ;
    buf_clk cell_6734 ( .C (clk), .D (signal_9279), .Q (signal_9280) ) ;
    buf_clk cell_6750 ( .C (clk), .D (signal_9295), .Q (signal_9296) ) ;
    buf_clk cell_6766 ( .C (clk), .D (signal_9311), .Q (signal_9312) ) ;
    buf_clk cell_6782 ( .C (clk), .D (signal_9327), .Q (signal_9328) ) ;
    buf_clk cell_6798 ( .C (clk), .D (signal_9343), .Q (signal_9344) ) ;
    buf_clk cell_6814 ( .C (clk), .D (signal_9359), .Q (signal_9360) ) ;
    buf_clk cell_6830 ( .C (clk), .D (signal_9375), .Q (signal_9376) ) ;
    buf_clk cell_6846 ( .C (clk), .D (signal_9391), .Q (signal_9392) ) ;
    buf_clk cell_6862 ( .C (clk), .D (signal_9407), .Q (signal_9408) ) ;
    buf_clk cell_6878 ( .C (clk), .D (signal_9423), .Q (signal_9424) ) ;
    buf_clk cell_6894 ( .C (clk), .D (signal_9439), .Q (signal_9440) ) ;
    buf_clk cell_6910 ( .C (clk), .D (signal_9455), .Q (signal_9456) ) ;
    buf_clk cell_6926 ( .C (clk), .D (signal_9471), .Q (signal_9472) ) ;
    buf_clk cell_6942 ( .C (clk), .D (signal_9487), .Q (signal_9488) ) ;
    buf_clk cell_6958 ( .C (clk), .D (signal_9503), .Q (signal_9504) ) ;
    buf_clk cell_6974 ( .C (clk), .D (signal_9519), .Q (signal_9520) ) ;
    buf_clk cell_6990 ( .C (clk), .D (signal_9535), .Q (signal_9536) ) ;
    buf_clk cell_7006 ( .C (clk), .D (signal_9551), .Q (signal_9552) ) ;
    buf_clk cell_7022 ( .C (clk), .D (signal_9567), .Q (signal_9568) ) ;
    buf_clk cell_7038 ( .C (clk), .D (signal_9583), .Q (signal_9584) ) ;
    buf_clk cell_7054 ( .C (clk), .D (signal_9599), .Q (signal_9600) ) ;
    buf_clk cell_7070 ( .C (clk), .D (signal_9615), .Q (signal_9616) ) ;
    buf_clk cell_7086 ( .C (clk), .D (signal_9631), .Q (signal_9632) ) ;
    buf_clk cell_7102 ( .C (clk), .D (signal_9647), .Q (signal_9648) ) ;
    buf_clk cell_7118 ( .C (clk), .D (signal_9663), .Q (signal_9664) ) ;
    buf_clk cell_7134 ( .C (clk), .D (signal_9679), .Q (signal_9680) ) ;
    buf_clk cell_7150 ( .C (clk), .D (signal_9695), .Q (signal_9696) ) ;
    buf_clk cell_7166 ( .C (clk), .D (signal_9711), .Q (signal_9712) ) ;
    buf_clk cell_7182 ( .C (clk), .D (signal_9727), .Q (signal_9728) ) ;
    buf_clk cell_7198 ( .C (clk), .D (signal_9743), .Q (signal_9744) ) ;
    buf_clk cell_7214 ( .C (clk), .D (signal_9759), .Q (signal_9760) ) ;
    buf_clk cell_7230 ( .C (clk), .D (signal_9775), .Q (signal_9776) ) ;
    buf_clk cell_7246 ( .C (clk), .D (signal_9791), .Q (signal_9792) ) ;
    buf_clk cell_7262 ( .C (clk), .D (signal_9807), .Q (signal_9808) ) ;
    buf_clk cell_7278 ( .C (clk), .D (signal_9823), .Q (signal_9824) ) ;
    buf_clk cell_7294 ( .C (clk), .D (signal_9839), .Q (signal_9840) ) ;
    buf_clk cell_7310 ( .C (clk), .D (signal_9855), .Q (signal_9856) ) ;
    buf_clk cell_7326 ( .C (clk), .D (signal_9871), .Q (signal_9872) ) ;
    buf_clk cell_7342 ( .C (clk), .D (signal_9887), .Q (signal_9888) ) ;
    buf_clk cell_7358 ( .C (clk), .D (signal_9903), .Q (signal_9904) ) ;
    buf_clk cell_7374 ( .C (clk), .D (signal_9919), .Q (signal_9920) ) ;
    buf_clk cell_7390 ( .C (clk), .D (signal_9935), .Q (signal_9936) ) ;
    buf_clk cell_7406 ( .C (clk), .D (signal_9951), .Q (signal_9952) ) ;
    buf_clk cell_7422 ( .C (clk), .D (signal_9967), .Q (signal_9968) ) ;
    buf_clk cell_7438 ( .C (clk), .D (signal_9983), .Q (signal_9984) ) ;
    buf_clk cell_7454 ( .C (clk), .D (signal_9999), .Q (signal_10000) ) ;
    buf_clk cell_7470 ( .C (clk), .D (signal_10015), .Q (signal_10016) ) ;
    buf_clk cell_7486 ( .C (clk), .D (signal_10031), .Q (signal_10032) ) ;
    buf_clk cell_7502 ( .C (clk), .D (signal_10047), .Q (signal_10048) ) ;
    buf_clk cell_7518 ( .C (clk), .D (signal_10063), .Q (signal_10064) ) ;
    buf_clk cell_7534 ( .C (clk), .D (signal_10079), .Q (signal_10080) ) ;
    buf_clk cell_7550 ( .C (clk), .D (signal_10095), .Q (signal_10096) ) ;
    buf_clk cell_7566 ( .C (clk), .D (signal_10111), .Q (signal_10112) ) ;
    buf_clk cell_7582 ( .C (clk), .D (signal_10127), .Q (signal_10128) ) ;
    buf_clk cell_7598 ( .C (clk), .D (signal_10143), .Q (signal_10144) ) ;
    buf_clk cell_7614 ( .C (clk), .D (signal_10159), .Q (signal_10160) ) ;
    buf_clk cell_7630 ( .C (clk), .D (signal_10175), .Q (signal_10176) ) ;
    buf_clk cell_7646 ( .C (clk), .D (signal_10191), .Q (signal_10192) ) ;
    buf_clk cell_7662 ( .C (clk), .D (signal_10207), .Q (signal_10208) ) ;
    buf_clk cell_7678 ( .C (clk), .D (signal_10223), .Q (signal_10224) ) ;
    buf_clk cell_7694 ( .C (clk), .D (signal_10239), .Q (signal_10240) ) ;
    buf_clk cell_7710 ( .C (clk), .D (signal_10255), .Q (signal_10256) ) ;
    buf_clk cell_7726 ( .C (clk), .D (signal_10271), .Q (signal_10272) ) ;
    buf_clk cell_7742 ( .C (clk), .D (signal_10287), .Q (signal_10288) ) ;
    buf_clk cell_7758 ( .C (clk), .D (signal_10303), .Q (signal_10304) ) ;
    buf_clk cell_7774 ( .C (clk), .D (signal_10319), .Q (signal_10320) ) ;
    buf_clk cell_7790 ( .C (clk), .D (signal_10335), .Q (signal_10336) ) ;
    buf_clk cell_7806 ( .C (clk), .D (signal_10351), .Q (signal_10352) ) ;
    buf_clk cell_7822 ( .C (clk), .D (signal_10367), .Q (signal_10368) ) ;
    buf_clk cell_7838 ( .C (clk), .D (signal_10383), .Q (signal_10384) ) ;
    buf_clk cell_7854 ( .C (clk), .D (signal_10399), .Q (signal_10400) ) ;
    buf_clk cell_7870 ( .C (clk), .D (signal_10415), .Q (signal_10416) ) ;
    buf_clk cell_7886 ( .C (clk), .D (signal_10431), .Q (signal_10432) ) ;
    buf_clk cell_7902 ( .C (clk), .D (signal_10447), .Q (signal_10448) ) ;
    buf_clk cell_7918 ( .C (clk), .D (signal_10463), .Q (signal_10464) ) ;
    buf_clk cell_7934 ( .C (clk), .D (signal_10479), .Q (signal_10480) ) ;
    buf_clk cell_7950 ( .C (clk), .D (signal_10495), .Q (signal_10496) ) ;
    buf_clk cell_7966 ( .C (clk), .D (signal_10511), .Q (signal_10512) ) ;
    buf_clk cell_7982 ( .C (clk), .D (signal_10527), .Q (signal_10528) ) ;
    buf_clk cell_7998 ( .C (clk), .D (signal_10543), .Q (signal_10544) ) ;
    buf_clk cell_8014 ( .C (clk), .D (signal_10559), .Q (signal_10560) ) ;
    buf_clk cell_8030 ( .C (clk), .D (signal_10575), .Q (signal_10576) ) ;
    buf_clk cell_8046 ( .C (clk), .D (signal_10591), .Q (signal_10592) ) ;
    buf_clk cell_8062 ( .C (clk), .D (signal_10607), .Q (signal_10608) ) ;
    buf_clk cell_8078 ( .C (clk), .D (signal_10623), .Q (signal_10624) ) ;
    buf_clk cell_8094 ( .C (clk), .D (signal_10639), .Q (signal_10640) ) ;
    buf_clk cell_8110 ( .C (clk), .D (signal_10655), .Q (signal_10656) ) ;
    buf_clk cell_8126 ( .C (clk), .D (signal_10671), .Q (signal_10672) ) ;
    buf_clk cell_8142 ( .C (clk), .D (signal_10687), .Q (signal_10688) ) ;
    buf_clk cell_8158 ( .C (clk), .D (signal_10703), .Q (signal_10704) ) ;
    buf_clk cell_8174 ( .C (clk), .D (signal_10719), .Q (signal_10720) ) ;
    buf_clk cell_8190 ( .C (clk), .D (signal_10735), .Q (signal_10736) ) ;
    buf_clk cell_8206 ( .C (clk), .D (signal_10751), .Q (signal_10752) ) ;
    buf_clk cell_8222 ( .C (clk), .D (signal_10767), .Q (signal_10768) ) ;
    buf_clk cell_8238 ( .C (clk), .D (signal_10783), .Q (signal_10784) ) ;
    buf_clk cell_8254 ( .C (clk), .D (signal_10799), .Q (signal_10800) ) ;
    buf_clk cell_8270 ( .C (clk), .D (signal_10815), .Q (signal_10816) ) ;
    buf_clk cell_8286 ( .C (clk), .D (signal_10831), .Q (signal_10832) ) ;
    buf_clk cell_8302 ( .C (clk), .D (signal_10847), .Q (signal_10848) ) ;
    buf_clk cell_8318 ( .C (clk), .D (signal_10863), .Q (signal_10864) ) ;
    buf_clk cell_8334 ( .C (clk), .D (signal_10879), .Q (signal_10880) ) ;
    buf_clk cell_8350 ( .C (clk), .D (signal_10895), .Q (signal_10896) ) ;
    buf_clk cell_8366 ( .C (clk), .D (signal_10911), .Q (signal_10912) ) ;
    buf_clk cell_8382 ( .C (clk), .D (signal_10927), .Q (signal_10928) ) ;
    buf_clk cell_8398 ( .C (clk), .D (signal_10943), .Q (signal_10944) ) ;
    buf_clk cell_8414 ( .C (clk), .D (signal_10959), .Q (signal_10960) ) ;
    buf_clk cell_8430 ( .C (clk), .D (signal_10975), .Q (signal_10976) ) ;
    buf_clk cell_8446 ( .C (clk), .D (signal_10991), .Q (signal_10992) ) ;
    buf_clk cell_8462 ( .C (clk), .D (signal_11007), .Q (signal_11008) ) ;
    buf_clk cell_8478 ( .C (clk), .D (signal_11023), .Q (signal_11024) ) ;
    buf_clk cell_8494 ( .C (clk), .D (signal_11039), .Q (signal_11040) ) ;
    buf_clk cell_8510 ( .C (clk), .D (signal_11055), .Q (signal_11056) ) ;
    buf_clk cell_8526 ( .C (clk), .D (signal_11071), .Q (signal_11072) ) ;
    buf_clk cell_8542 ( .C (clk), .D (signal_11087), .Q (signal_11088) ) ;
    buf_clk cell_8558 ( .C (clk), .D (signal_11103), .Q (signal_11104) ) ;
    buf_clk cell_8574 ( .C (clk), .D (signal_11119), .Q (signal_11120) ) ;
    buf_clk cell_8590 ( .C (clk), .D (signal_11135), .Q (signal_11136) ) ;
    buf_clk cell_8606 ( .C (clk), .D (signal_11151), .Q (signal_11152) ) ;
    buf_clk cell_8622 ( .C (clk), .D (signal_11167), .Q (signal_11168) ) ;
    buf_clk cell_8638 ( .C (clk), .D (signal_11183), .Q (signal_11184) ) ;
    buf_clk cell_8654 ( .C (clk), .D (signal_11199), .Q (signal_11200) ) ;
    buf_clk cell_8670 ( .C (clk), .D (signal_11215), .Q (signal_11216) ) ;
    buf_clk cell_8686 ( .C (clk), .D (signal_11231), .Q (signal_11232) ) ;
    buf_clk cell_8702 ( .C (clk), .D (signal_11247), .Q (signal_11248) ) ;
    buf_clk cell_8718 ( .C (clk), .D (signal_11263), .Q (signal_11264) ) ;
    buf_clk cell_8734 ( .C (clk), .D (signal_11279), .Q (signal_11280) ) ;
    buf_clk cell_8750 ( .C (clk), .D (signal_11295), .Q (signal_11296) ) ;
    buf_clk cell_8766 ( .C (clk), .D (signal_11311), .Q (signal_11312) ) ;
    buf_clk cell_8782 ( .C (clk), .D (signal_11327), .Q (signal_11328) ) ;
    buf_clk cell_8798 ( .C (clk), .D (signal_11343), .Q (signal_11344) ) ;
    buf_clk cell_8814 ( .C (clk), .D (signal_11359), .Q (signal_11360) ) ;
    buf_clk cell_8830 ( .C (clk), .D (signal_11375), .Q (signal_11376) ) ;
    buf_clk cell_8846 ( .C (clk), .D (signal_11391), .Q (signal_11392) ) ;
    buf_clk cell_8862 ( .C (clk), .D (signal_11407), .Q (signal_11408) ) ;
    buf_clk cell_8878 ( .C (clk), .D (signal_11423), .Q (signal_11424) ) ;
    buf_clk cell_8894 ( .C (clk), .D (signal_11439), .Q (signal_11440) ) ;
    buf_clk cell_8910 ( .C (clk), .D (signal_11455), .Q (signal_11456) ) ;
    buf_clk cell_8926 ( .C (clk), .D (signal_11471), .Q (signal_11472) ) ;
    buf_clk cell_8942 ( .C (clk), .D (signal_11487), .Q (signal_11488) ) ;
    buf_clk cell_8958 ( .C (clk), .D (signal_11503), .Q (signal_11504) ) ;
    buf_clk cell_8974 ( .C (clk), .D (signal_11519), .Q (signal_11520) ) ;
    buf_clk cell_8990 ( .C (clk), .D (signal_11535), .Q (signal_11536) ) ;
    buf_clk cell_9006 ( .C (clk), .D (signal_11551), .Q (signal_11552) ) ;
    buf_clk cell_9022 ( .C (clk), .D (signal_11567), .Q (signal_11568) ) ;
    buf_clk cell_9038 ( .C (clk), .D (signal_11583), .Q (signal_11584) ) ;
    buf_clk cell_9054 ( .C (clk), .D (signal_11599), .Q (signal_11600) ) ;
    buf_clk cell_9070 ( .C (clk), .D (signal_11615), .Q (signal_11616) ) ;
    buf_clk cell_9086 ( .C (clk), .D (signal_11631), .Q (signal_11632) ) ;
    buf_clk cell_9102 ( .C (clk), .D (signal_11647), .Q (signal_11648) ) ;
    buf_clk cell_9118 ( .C (clk), .D (signal_11663), .Q (signal_11664) ) ;
    buf_clk cell_9134 ( .C (clk), .D (signal_11679), .Q (signal_11680) ) ;
    buf_clk cell_9150 ( .C (clk), .D (signal_11695), .Q (signal_11696) ) ;
    buf_clk cell_9166 ( .C (clk), .D (signal_11711), .Q (signal_11712) ) ;
    buf_clk cell_9182 ( .C (clk), .D (signal_11727), .Q (signal_11728) ) ;
    buf_clk cell_9198 ( .C (clk), .D (signal_11743), .Q (signal_11744) ) ;
    buf_clk cell_9214 ( .C (clk), .D (signal_11759), .Q (signal_11760) ) ;
    buf_clk cell_9230 ( .C (clk), .D (signal_11775), .Q (signal_11776) ) ;
    buf_clk cell_9246 ( .C (clk), .D (signal_11791), .Q (signal_11792) ) ;
    buf_clk cell_9262 ( .C (clk), .D (signal_11807), .Q (signal_11808) ) ;
    buf_clk cell_9278 ( .C (clk), .D (signal_11823), .Q (signal_11824) ) ;
    buf_clk cell_9294 ( .C (clk), .D (signal_11839), .Q (signal_11840) ) ;
    buf_clk cell_9310 ( .C (clk), .D (signal_11855), .Q (signal_11856) ) ;
    buf_clk cell_9326 ( .C (clk), .D (signal_11871), .Q (signal_11872) ) ;
    buf_clk cell_9342 ( .C (clk), .D (signal_11887), .Q (signal_11888) ) ;
    buf_clk cell_9358 ( .C (clk), .D (signal_11903), .Q (signal_11904) ) ;
    buf_clk cell_9374 ( .C (clk), .D (signal_11919), .Q (signal_11920) ) ;
    buf_clk cell_9390 ( .C (clk), .D (signal_11935), .Q (signal_11936) ) ;
    buf_clk cell_9406 ( .C (clk), .D (signal_11951), .Q (signal_11952) ) ;
    buf_clk cell_9422 ( .C (clk), .D (signal_11967), .Q (signal_11968) ) ;
    buf_clk cell_9438 ( .C (clk), .D (signal_11983), .Q (signal_11984) ) ;
    buf_clk cell_9454 ( .C (clk), .D (signal_11999), .Q (signal_12000) ) ;
    buf_clk cell_9470 ( .C (clk), .D (signal_12015), .Q (signal_12016) ) ;
    buf_clk cell_9486 ( .C (clk), .D (signal_12031), .Q (signal_12032) ) ;
    buf_clk cell_9502 ( .C (clk), .D (signal_12047), .Q (signal_12048) ) ;
    buf_clk cell_9518 ( .C (clk), .D (signal_12063), .Q (signal_12064) ) ;
    buf_clk cell_9534 ( .C (clk), .D (signal_12079), .Q (signal_12080) ) ;
    buf_clk cell_9550 ( .C (clk), .D (signal_12095), .Q (signal_12096) ) ;
    buf_clk cell_9566 ( .C (clk), .D (signal_12111), .Q (signal_12112) ) ;
    buf_clk cell_9582 ( .C (clk), .D (signal_12127), .Q (signal_12128) ) ;
    buf_clk cell_9598 ( .C (clk), .D (signal_12143), .Q (signal_12144) ) ;
    buf_clk cell_9614 ( .C (clk), .D (signal_12159), .Q (signal_12160) ) ;
    buf_clk cell_9630 ( .C (clk), .D (signal_12175), .Q (signal_12176) ) ;
    buf_clk cell_9646 ( .C (clk), .D (signal_12191), .Q (signal_12192) ) ;
    buf_clk cell_9662 ( .C (clk), .D (signal_12207), .Q (signal_12208) ) ;
    buf_clk cell_9678 ( .C (clk), .D (signal_12223), .Q (signal_12224) ) ;
    buf_clk cell_9694 ( .C (clk), .D (signal_12239), .Q (signal_12240) ) ;
    buf_clk cell_9710 ( .C (clk), .D (signal_12255), .Q (signal_12256) ) ;
    buf_clk cell_9726 ( .C (clk), .D (signal_12271), .Q (signal_12272) ) ;
    buf_clk cell_9742 ( .C (clk), .D (signal_12287), .Q (signal_12288) ) ;
    buf_clk cell_9758 ( .C (clk), .D (signal_12303), .Q (signal_12304) ) ;
    buf_clk cell_9774 ( .C (clk), .D (signal_12319), .Q (signal_12320) ) ;
    buf_clk cell_9790 ( .C (clk), .D (signal_12335), .Q (signal_12336) ) ;
    buf_clk cell_9806 ( .C (clk), .D (signal_12351), .Q (signal_12352) ) ;
    buf_clk cell_9822 ( .C (clk), .D (signal_12367), .Q (signal_12368) ) ;
    buf_clk cell_9838 ( .C (clk), .D (signal_12383), .Q (signal_12384) ) ;
    buf_clk cell_9854 ( .C (clk), .D (signal_12399), .Q (signal_12400) ) ;
    buf_clk cell_9870 ( .C (clk), .D (signal_12415), .Q (signal_12416) ) ;
    buf_clk cell_9886 ( .C (clk), .D (signal_12431), .Q (signal_12432) ) ;
    buf_clk cell_9902 ( .C (clk), .D (signal_12447), .Q (signal_12448) ) ;
    buf_clk cell_9918 ( .C (clk), .D (signal_12463), .Q (signal_12464) ) ;
    buf_clk cell_9934 ( .C (clk), .D (signal_12479), .Q (signal_12480) ) ;
    buf_clk cell_9950 ( .C (clk), .D (signal_12495), .Q (signal_12496) ) ;
    buf_clk cell_9966 ( .C (clk), .D (signal_12511), .Q (signal_12512) ) ;
    buf_clk cell_9982 ( .C (clk), .D (signal_12527), .Q (signal_12528) ) ;
    buf_clk cell_9998 ( .C (clk), .D (signal_12543), .Q (signal_12544) ) ;
    buf_clk cell_10014 ( .C (clk), .D (signal_12559), .Q (signal_12560) ) ;
    buf_clk cell_10030 ( .C (clk), .D (signal_12575), .Q (signal_12576) ) ;
    buf_clk cell_10046 ( .C (clk), .D (signal_12591), .Q (signal_12592) ) ;
    buf_clk cell_10062 ( .C (clk), .D (signal_12607), .Q (signal_12608) ) ;
    buf_clk cell_10078 ( .C (clk), .D (signal_12623), .Q (signal_12624) ) ;
    buf_clk cell_10094 ( .C (clk), .D (signal_12639), .Q (signal_12640) ) ;
    buf_clk cell_10110 ( .C (clk), .D (signal_12655), .Q (signal_12656) ) ;
    buf_clk cell_10126 ( .C (clk), .D (signal_12671), .Q (signal_12672) ) ;
    buf_clk cell_10142 ( .C (clk), .D (signal_12687), .Q (signal_12688) ) ;
    buf_clk cell_10158 ( .C (clk), .D (signal_12703), .Q (signal_12704) ) ;
    buf_clk cell_10174 ( .C (clk), .D (signal_12719), .Q (signal_12720) ) ;
    buf_clk cell_10190 ( .C (clk), .D (signal_12735), .Q (signal_12736) ) ;
    buf_clk cell_10206 ( .C (clk), .D (signal_12751), .Q (signal_12752) ) ;
    buf_clk cell_10222 ( .C (clk), .D (signal_12767), .Q (signal_12768) ) ;
    buf_clk cell_10238 ( .C (clk), .D (signal_12783), .Q (signal_12784) ) ;
    buf_clk cell_10254 ( .C (clk), .D (signal_12799), .Q (signal_12800) ) ;
    buf_clk cell_10270 ( .C (clk), .D (signal_12815), .Q (signal_12816) ) ;
    buf_clk cell_10286 ( .C (clk), .D (signal_12831), .Q (signal_12832) ) ;
    buf_clk cell_10302 ( .C (clk), .D (signal_12847), .Q (signal_12848) ) ;
    buf_clk cell_10318 ( .C (clk), .D (signal_12863), .Q (signal_12864) ) ;
    buf_clk cell_10334 ( .C (clk), .D (signal_12879), .Q (signal_12880) ) ;
    buf_clk cell_10350 ( .C (clk), .D (signal_12895), .Q (signal_12896) ) ;
    buf_clk cell_10366 ( .C (clk), .D (signal_12911), .Q (signal_12912) ) ;
    buf_clk cell_10382 ( .C (clk), .D (signal_12927), .Q (signal_12928) ) ;
    buf_clk cell_10398 ( .C (clk), .D (signal_12943), .Q (signal_12944) ) ;
    buf_clk cell_10414 ( .C (clk), .D (signal_12959), .Q (signal_12960) ) ;
    buf_clk cell_10430 ( .C (clk), .D (signal_12975), .Q (signal_12976) ) ;
    buf_clk cell_10446 ( .C (clk), .D (signal_12991), .Q (signal_12992) ) ;
    buf_clk cell_10462 ( .C (clk), .D (signal_13007), .Q (signal_13008) ) ;
    buf_clk cell_10478 ( .C (clk), .D (signal_13023), .Q (signal_13024) ) ;
    buf_clk cell_10494 ( .C (clk), .D (signal_13039), .Q (signal_13040) ) ;
    buf_clk cell_10510 ( .C (clk), .D (signal_13055), .Q (signal_13056) ) ;
    buf_clk cell_10526 ( .C (clk), .D (signal_13071), .Q (signal_13072) ) ;
    buf_clk cell_10542 ( .C (clk), .D (signal_13087), .Q (signal_13088) ) ;
    buf_clk cell_10558 ( .C (clk), .D (signal_13103), .Q (signal_13104) ) ;
    buf_clk cell_10574 ( .C (clk), .D (signal_13119), .Q (signal_13120) ) ;
    buf_clk cell_10590 ( .C (clk), .D (signal_13135), .Q (signal_13136) ) ;
    buf_clk cell_10606 ( .C (clk), .D (signal_13151), .Q (signal_13152) ) ;
    buf_clk cell_10622 ( .C (clk), .D (signal_13167), .Q (signal_13168) ) ;
    buf_clk cell_10638 ( .C (clk), .D (signal_13183), .Q (signal_13184) ) ;
    buf_clk cell_10654 ( .C (clk), .D (signal_13199), .Q (signal_13200) ) ;
    buf_clk cell_10670 ( .C (clk), .D (signal_13215), .Q (signal_13216) ) ;
    buf_clk cell_10686 ( .C (clk), .D (signal_13231), .Q (signal_13232) ) ;
    buf_clk cell_10702 ( .C (clk), .D (signal_13247), .Q (signal_13248) ) ;
    buf_clk cell_10718 ( .C (clk), .D (signal_13263), .Q (signal_13264) ) ;
    buf_clk cell_10734 ( .C (clk), .D (signal_13279), .Q (signal_13280) ) ;
    buf_clk cell_10750 ( .C (clk), .D (signal_13295), .Q (signal_13296) ) ;
    buf_clk cell_10766 ( .C (clk), .D (signal_13311), .Q (signal_13312) ) ;
    buf_clk cell_10782 ( .C (clk), .D (signal_13327), .Q (signal_13328) ) ;
    buf_clk cell_10798 ( .C (clk), .D (signal_13343), .Q (signal_13344) ) ;
    buf_clk cell_10814 ( .C (clk), .D (signal_13359), .Q (signal_13360) ) ;
    buf_clk cell_10830 ( .C (clk), .D (signal_13375), .Q (signal_13376) ) ;
    buf_clk cell_10846 ( .C (clk), .D (signal_13391), .Q (signal_13392) ) ;
    buf_clk cell_10862 ( .C (clk), .D (signal_13407), .Q (signal_13408) ) ;
    buf_clk cell_10878 ( .C (clk), .D (signal_13423), .Q (signal_13424) ) ;
    buf_clk cell_10894 ( .C (clk), .D (signal_13439), .Q (signal_13440) ) ;
    buf_clk cell_10910 ( .C (clk), .D (signal_13455), .Q (signal_13456) ) ;
    buf_clk cell_10926 ( .C (clk), .D (signal_13471), .Q (signal_13472) ) ;
    buf_clk cell_10942 ( .C (clk), .D (signal_13487), .Q (signal_13488) ) ;
    buf_clk cell_10958 ( .C (clk), .D (signal_13503), .Q (signal_13504) ) ;
    buf_clk cell_10974 ( .C (clk), .D (signal_13519), .Q (signal_13520) ) ;
    buf_clk cell_10990 ( .C (clk), .D (signal_13535), .Q (signal_13536) ) ;
    buf_clk cell_11006 ( .C (clk), .D (signal_13551), .Q (signal_13552) ) ;
    buf_clk cell_11022 ( .C (clk), .D (signal_13567), .Q (signal_13568) ) ;
    buf_clk cell_11038 ( .C (clk), .D (signal_13583), .Q (signal_13584) ) ;
    buf_clk cell_11054 ( .C (clk), .D (signal_13599), .Q (signal_13600) ) ;
    buf_clk cell_11070 ( .C (clk), .D (signal_13615), .Q (signal_13616) ) ;
    buf_clk cell_11086 ( .C (clk), .D (signal_13631), .Q (signal_13632) ) ;
    buf_clk cell_11102 ( .C (clk), .D (signal_13647), .Q (signal_13648) ) ;
    buf_clk cell_11118 ( .C (clk), .D (signal_13663), .Q (signal_13664) ) ;
    buf_clk cell_11134 ( .C (clk), .D (signal_13679), .Q (signal_13680) ) ;
    buf_clk cell_11150 ( .C (clk), .D (signal_13695), .Q (signal_13696) ) ;
    buf_clk cell_11166 ( .C (clk), .D (signal_13711), .Q (signal_13712) ) ;
    buf_clk cell_11182 ( .C (clk), .D (signal_13727), .Q (signal_13728) ) ;
    buf_clk cell_11198 ( .C (clk), .D (signal_13743), .Q (signal_13744) ) ;
    buf_clk cell_11214 ( .C (clk), .D (signal_13759), .Q (signal_13760) ) ;
    buf_clk cell_11230 ( .C (clk), .D (signal_13775), .Q (signal_13776) ) ;
    buf_clk cell_11246 ( .C (clk), .D (signal_13791), .Q (signal_13792) ) ;
    buf_clk cell_11262 ( .C (clk), .D (signal_13807), .Q (signal_13808) ) ;
    buf_clk cell_11278 ( .C (clk), .D (signal_13823), .Q (signal_13824) ) ;
    buf_clk cell_11294 ( .C (clk), .D (signal_13839), .Q (signal_13840) ) ;
    buf_clk cell_11310 ( .C (clk), .D (signal_13855), .Q (signal_13856) ) ;
    buf_clk cell_11326 ( .C (clk), .D (signal_13871), .Q (signal_13872) ) ;
    buf_clk cell_11342 ( .C (clk), .D (signal_13887), .Q (signal_13888) ) ;
    buf_clk cell_11358 ( .C (clk), .D (signal_13903), .Q (signal_13904) ) ;
    buf_clk cell_11374 ( .C (clk), .D (signal_13919), .Q (signal_13920) ) ;
    buf_clk cell_11390 ( .C (clk), .D (signal_13935), .Q (signal_13936) ) ;
    buf_clk cell_11406 ( .C (clk), .D (signal_13951), .Q (signal_13952) ) ;
    buf_clk cell_11422 ( .C (clk), .D (signal_13967), .Q (signal_13968) ) ;
    buf_clk cell_11438 ( .C (clk), .D (signal_13983), .Q (signal_13984) ) ;
    buf_clk cell_11454 ( .C (clk), .D (signal_13999), .Q (signal_14000) ) ;
    buf_clk cell_11470 ( .C (clk), .D (signal_14015), .Q (signal_14016) ) ;
    buf_clk cell_11486 ( .C (clk), .D (signal_14031), .Q (signal_14032) ) ;
    buf_clk cell_11502 ( .C (clk), .D (signal_14047), .Q (signal_14048) ) ;
    buf_clk cell_11518 ( .C (clk), .D (signal_14063), .Q (signal_14064) ) ;
    buf_clk cell_11534 ( .C (clk), .D (signal_14079), .Q (signal_14080) ) ;
    buf_clk cell_11550 ( .C (clk), .D (signal_14095), .Q (signal_14096) ) ;
    buf_clk cell_11566 ( .C (clk), .D (signal_14111), .Q (signal_14112) ) ;
    buf_clk cell_11582 ( .C (clk), .D (signal_14127), .Q (signal_14128) ) ;
    buf_clk cell_11598 ( .C (clk), .D (signal_14143), .Q (signal_14144) ) ;
    buf_clk cell_11614 ( .C (clk), .D (signal_14159), .Q (signal_14160) ) ;
    buf_clk cell_11630 ( .C (clk), .D (signal_14175), .Q (signal_14176) ) ;
    buf_clk cell_11646 ( .C (clk), .D (signal_14191), .Q (signal_14192) ) ;
    buf_clk cell_11662 ( .C (clk), .D (signal_14207), .Q (signal_14208) ) ;
    buf_clk cell_11678 ( .C (clk), .D (signal_14223), .Q (signal_14224) ) ;
    buf_clk cell_11694 ( .C (clk), .D (signal_14239), .Q (signal_14240) ) ;
    buf_clk cell_11710 ( .C (clk), .D (signal_14255), .Q (signal_14256) ) ;
    buf_clk cell_11726 ( .C (clk), .D (signal_14271), .Q (signal_14272) ) ;
    buf_clk cell_11742 ( .C (clk), .D (signal_14287), .Q (signal_14288) ) ;
    buf_clk cell_11758 ( .C (clk), .D (signal_14303), .Q (signal_14304) ) ;
    buf_clk cell_11774 ( .C (clk), .D (signal_14319), .Q (signal_14320) ) ;
    buf_clk cell_11790 ( .C (clk), .D (signal_14335), .Q (signal_14336) ) ;
    buf_clk cell_11806 ( .C (clk), .D (signal_14351), .Q (signal_14352) ) ;
    buf_clk cell_11822 ( .C (clk), .D (signal_14367), .Q (signal_14368) ) ;
    buf_clk cell_11838 ( .C (clk), .D (signal_14383), .Q (signal_14384) ) ;
    buf_clk cell_11854 ( .C (clk), .D (signal_14399), .Q (signal_14400) ) ;
    buf_clk cell_11870 ( .C (clk), .D (signal_14415), .Q (signal_14416) ) ;
    buf_clk cell_11886 ( .C (clk), .D (signal_14431), .Q (signal_14432) ) ;
    buf_clk cell_11902 ( .C (clk), .D (signal_14447), .Q (signal_14448) ) ;
    buf_clk cell_11918 ( .C (clk), .D (signal_14463), .Q (signal_14464) ) ;
    buf_clk cell_11934 ( .C (clk), .D (signal_14479), .Q (signal_14480) ) ;
    buf_clk cell_11950 ( .C (clk), .D (signal_14495), .Q (signal_14496) ) ;
    buf_clk cell_11966 ( .C (clk), .D (signal_14511), .Q (signal_14512) ) ;
    buf_clk cell_11982 ( .C (clk), .D (signal_14527), .Q (signal_14528) ) ;
    buf_clk cell_11998 ( .C (clk), .D (signal_14543), .Q (signal_14544) ) ;
    buf_clk cell_12014 ( .C (clk), .D (signal_14559), .Q (signal_14560) ) ;
    buf_clk cell_12030 ( .C (clk), .D (signal_14575), .Q (signal_14576) ) ;
    buf_clk cell_12046 ( .C (clk), .D (signal_14591), .Q (signal_14592) ) ;
    buf_clk cell_12062 ( .C (clk), .D (signal_14607), .Q (signal_14608) ) ;
    buf_clk cell_12078 ( .C (clk), .D (signal_14623), .Q (signal_14624) ) ;
    buf_clk cell_12094 ( .C (clk), .D (signal_14639), .Q (signal_14640) ) ;
    buf_clk cell_12110 ( .C (clk), .D (signal_14655), .Q (signal_14656) ) ;
    buf_clk cell_12126 ( .C (clk), .D (signal_14671), .Q (signal_14672) ) ;
    buf_clk cell_12142 ( .C (clk), .D (signal_14687), .Q (signal_14688) ) ;
    buf_clk cell_12158 ( .C (clk), .D (signal_14703), .Q (signal_14704) ) ;
    buf_clk cell_12174 ( .C (clk), .D (signal_14719), .Q (signal_14720) ) ;
    buf_clk cell_12190 ( .C (clk), .D (signal_14735), .Q (signal_14736) ) ;
    buf_clk cell_12206 ( .C (clk), .D (signal_14751), .Q (signal_14752) ) ;
    buf_clk cell_12222 ( .C (clk), .D (signal_14767), .Q (signal_14768) ) ;
    buf_clk cell_12238 ( .C (clk), .D (signal_14783), .Q (signal_14784) ) ;
    buf_clk cell_12254 ( .C (clk), .D (signal_14799), .Q (signal_14800) ) ;
    buf_clk cell_12270 ( .C (clk), .D (signal_14815), .Q (signal_14816) ) ;
    buf_clk cell_12286 ( .C (clk), .D (signal_14831), .Q (signal_14832) ) ;
    buf_clk cell_12302 ( .C (clk), .D (signal_14847), .Q (signal_14848) ) ;
    buf_clk cell_12318 ( .C (clk), .D (signal_14863), .Q (signal_14864) ) ;
    buf_clk cell_12334 ( .C (clk), .D (signal_14879), .Q (signal_14880) ) ;
    buf_clk cell_12350 ( .C (clk), .D (signal_14895), .Q (signal_14896) ) ;
    buf_clk cell_12366 ( .C (clk), .D (signal_14911), .Q (signal_14912) ) ;
    buf_clk cell_12382 ( .C (clk), .D (signal_14927), .Q (signal_14928) ) ;

    /* cells in depth 3 */
    buf_clk cell_2153 ( .C (clk), .D (signal_4696), .Q (signal_4699) ) ;
    buf_clk cell_2155 ( .C (clk), .D (signal_4698), .Q (signal_4701) ) ;
    buf_clk cell_2157 ( .C (clk), .D (signal_1984), .Q (signal_4703) ) ;
    buf_clk cell_2159 ( .C (clk), .D (signal_3275), .Q (signal_4705) ) ;
    buf_clk cell_2161 ( .C (clk), .D (signal_1985), .Q (signal_4707) ) ;
    buf_clk cell_2163 ( .C (clk), .D (signal_3276), .Q (signal_4709) ) ;
    buf_clk cell_2165 ( .C (clk), .D (signal_1982), .Q (signal_4711) ) ;
    buf_clk cell_2167 ( .C (clk), .D (signal_3273), .Q (signal_4713) ) ;
    buf_clk cell_2171 ( .C (clk), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_2175 ( .C (clk), .D (signal_4720), .Q (signal_4721) ) ;
    buf_clk cell_2177 ( .C (clk), .D (signal_1983), .Q (signal_4723) ) ;
    buf_clk cell_2179 ( .C (clk), .D (signal_3274), .Q (signal_4725) ) ;
    buf_clk cell_2181 ( .C (clk), .D (signal_1986), .Q (signal_4727) ) ;
    buf_clk cell_2183 ( .C (clk), .D (signal_3277), .Q (signal_4729) ) ;
    buf_clk cell_2299 ( .C (clk), .D (signal_4844), .Q (signal_4845) ) ;
    buf_clk cell_2307 ( .C (clk), .D (signal_4852), .Q (signal_4853) ) ;
    buf_clk cell_2343 ( .C (clk), .D (signal_4888), .Q (signal_4889) ) ;
    buf_clk cell_2353 ( .C (clk), .D (signal_4898), .Q (signal_4899) ) ;
    buf_clk cell_2363 ( .C (clk), .D (signal_4908), .Q (signal_4909) ) ;
    buf_clk cell_2375 ( .C (clk), .D (signal_4920), .Q (signal_4921) ) ;
    buf_clk cell_2387 ( .C (clk), .D (signal_4932), .Q (signal_4933) ) ;
    buf_clk cell_2403 ( .C (clk), .D (signal_4948), .Q (signal_4949) ) ;
    buf_clk cell_2419 ( .C (clk), .D (signal_4964), .Q (signal_4965) ) ;
    buf_clk cell_2435 ( .C (clk), .D (signal_4980), .Q (signal_4981) ) ;
    buf_clk cell_2451 ( .C (clk), .D (signal_4996), .Q (signal_4997) ) ;
    buf_clk cell_2467 ( .C (clk), .D (signal_5012), .Q (signal_5013) ) ;
    buf_clk cell_2483 ( .C (clk), .D (signal_5028), .Q (signal_5029) ) ;
    buf_clk cell_2499 ( .C (clk), .D (signal_5044), .Q (signal_5045) ) ;
    buf_clk cell_2515 ( .C (clk), .D (signal_5060), .Q (signal_5061) ) ;
    buf_clk cell_2531 ( .C (clk), .D (signal_5076), .Q (signal_5077) ) ;
    buf_clk cell_2547 ( .C (clk), .D (signal_5092), .Q (signal_5093) ) ;
    buf_clk cell_2563 ( .C (clk), .D (signal_5108), .Q (signal_5109) ) ;
    buf_clk cell_2579 ( .C (clk), .D (signal_5124), .Q (signal_5125) ) ;
    buf_clk cell_2595 ( .C (clk), .D (signal_5140), .Q (signal_5141) ) ;
    buf_clk cell_2611 ( .C (clk), .D (signal_5156), .Q (signal_5157) ) ;
    buf_clk cell_2627 ( .C (clk), .D (signal_5172), .Q (signal_5173) ) ;
    buf_clk cell_2643 ( .C (clk), .D (signal_5188), .Q (signal_5189) ) ;
    buf_clk cell_2659 ( .C (clk), .D (signal_5204), .Q (signal_5205) ) ;
    buf_clk cell_2675 ( .C (clk), .D (signal_5220), .Q (signal_5221) ) ;
    buf_clk cell_2691 ( .C (clk), .D (signal_5236), .Q (signal_5237) ) ;
    buf_clk cell_2707 ( .C (clk), .D (signal_5252), .Q (signal_5253) ) ;
    buf_clk cell_2723 ( .C (clk), .D (signal_5268), .Q (signal_5269) ) ;
    buf_clk cell_2739 ( .C (clk), .D (signal_5284), .Q (signal_5285) ) ;
    buf_clk cell_2755 ( .C (clk), .D (signal_5300), .Q (signal_5301) ) ;
    buf_clk cell_2771 ( .C (clk), .D (signal_5316), .Q (signal_5317) ) ;
    buf_clk cell_2787 ( .C (clk), .D (signal_5332), .Q (signal_5333) ) ;
    buf_clk cell_2803 ( .C (clk), .D (signal_5348), .Q (signal_5349) ) ;
    buf_clk cell_2819 ( .C (clk), .D (signal_5364), .Q (signal_5365) ) ;
    buf_clk cell_2835 ( .C (clk), .D (signal_5380), .Q (signal_5381) ) ;
    buf_clk cell_2851 ( .C (clk), .D (signal_5396), .Q (signal_5397) ) ;
    buf_clk cell_2867 ( .C (clk), .D (signal_5412), .Q (signal_5413) ) ;
    buf_clk cell_2883 ( .C (clk), .D (signal_5428), .Q (signal_5429) ) ;
    buf_clk cell_2899 ( .C (clk), .D (signal_5444), .Q (signal_5445) ) ;
    buf_clk cell_2915 ( .C (clk), .D (signal_5460), .Q (signal_5461) ) ;
    buf_clk cell_2931 ( .C (clk), .D (signal_5476), .Q (signal_5477) ) ;
    buf_clk cell_2947 ( .C (clk), .D (signal_5492), .Q (signal_5493) ) ;
    buf_clk cell_2963 ( .C (clk), .D (signal_5508), .Q (signal_5509) ) ;
    buf_clk cell_2979 ( .C (clk), .D (signal_5524), .Q (signal_5525) ) ;
    buf_clk cell_2995 ( .C (clk), .D (signal_5540), .Q (signal_5541) ) ;
    buf_clk cell_3011 ( .C (clk), .D (signal_5556), .Q (signal_5557) ) ;
    buf_clk cell_3027 ( .C (clk), .D (signal_5572), .Q (signal_5573) ) ;
    buf_clk cell_3043 ( .C (clk), .D (signal_5588), .Q (signal_5589) ) ;
    buf_clk cell_3059 ( .C (clk), .D (signal_5604), .Q (signal_5605) ) ;
    buf_clk cell_3075 ( .C (clk), .D (signal_5620), .Q (signal_5621) ) ;
    buf_clk cell_3091 ( .C (clk), .D (signal_5636), .Q (signal_5637) ) ;
    buf_clk cell_3107 ( .C (clk), .D (signal_5652), .Q (signal_5653) ) ;
    buf_clk cell_3123 ( .C (clk), .D (signal_5668), .Q (signal_5669) ) ;
    buf_clk cell_3139 ( .C (clk), .D (signal_5684), .Q (signal_5685) ) ;
    buf_clk cell_3155 ( .C (clk), .D (signal_5700), .Q (signal_5701) ) ;
    buf_clk cell_3171 ( .C (clk), .D (signal_5716), .Q (signal_5717) ) ;
    buf_clk cell_3187 ( .C (clk), .D (signal_5732), .Q (signal_5733) ) ;
    buf_clk cell_3203 ( .C (clk), .D (signal_5748), .Q (signal_5749) ) ;
    buf_clk cell_3219 ( .C (clk), .D (signal_5764), .Q (signal_5765) ) ;
    buf_clk cell_3235 ( .C (clk), .D (signal_5780), .Q (signal_5781) ) ;
    buf_clk cell_3251 ( .C (clk), .D (signal_5796), .Q (signal_5797) ) ;
    buf_clk cell_3267 ( .C (clk), .D (signal_5812), .Q (signal_5813) ) ;
    buf_clk cell_3283 ( .C (clk), .D (signal_5828), .Q (signal_5829) ) ;
    buf_clk cell_3299 ( .C (clk), .D (signal_5844), .Q (signal_5845) ) ;
    buf_clk cell_3315 ( .C (clk), .D (signal_5860), .Q (signal_5861) ) ;
    buf_clk cell_3331 ( .C (clk), .D (signal_5876), .Q (signal_5877) ) ;
    buf_clk cell_3347 ( .C (clk), .D (signal_5892), .Q (signal_5893) ) ;
    buf_clk cell_3363 ( .C (clk), .D (signal_5908), .Q (signal_5909) ) ;
    buf_clk cell_3379 ( .C (clk), .D (signal_5924), .Q (signal_5925) ) ;
    buf_clk cell_3395 ( .C (clk), .D (signal_5940), .Q (signal_5941) ) ;
    buf_clk cell_3411 ( .C (clk), .D (signal_5956), .Q (signal_5957) ) ;
    buf_clk cell_3427 ( .C (clk), .D (signal_5972), .Q (signal_5973) ) ;
    buf_clk cell_3443 ( .C (clk), .D (signal_5988), .Q (signal_5989) ) ;
    buf_clk cell_3459 ( .C (clk), .D (signal_6004), .Q (signal_6005) ) ;
    buf_clk cell_3475 ( .C (clk), .D (signal_6020), .Q (signal_6021) ) ;
    buf_clk cell_3491 ( .C (clk), .D (signal_6036), .Q (signal_6037) ) ;
    buf_clk cell_3507 ( .C (clk), .D (signal_6052), .Q (signal_6053) ) ;
    buf_clk cell_3523 ( .C (clk), .D (signal_6068), .Q (signal_6069) ) ;
    buf_clk cell_3539 ( .C (clk), .D (signal_6084), .Q (signal_6085) ) ;
    buf_clk cell_3555 ( .C (clk), .D (signal_6100), .Q (signal_6101) ) ;
    buf_clk cell_3571 ( .C (clk), .D (signal_6116), .Q (signal_6117) ) ;
    buf_clk cell_3587 ( .C (clk), .D (signal_6132), .Q (signal_6133) ) ;
    buf_clk cell_3603 ( .C (clk), .D (signal_6148), .Q (signal_6149) ) ;
    buf_clk cell_3619 ( .C (clk), .D (signal_6164), .Q (signal_6165) ) ;
    buf_clk cell_3635 ( .C (clk), .D (signal_6180), .Q (signal_6181) ) ;
    buf_clk cell_3651 ( .C (clk), .D (signal_6196), .Q (signal_6197) ) ;
    buf_clk cell_3667 ( .C (clk), .D (signal_6212), .Q (signal_6213) ) ;
    buf_clk cell_3683 ( .C (clk), .D (signal_6228), .Q (signal_6229) ) ;
    buf_clk cell_3699 ( .C (clk), .D (signal_6244), .Q (signal_6245) ) ;
    buf_clk cell_3715 ( .C (clk), .D (signal_6260), .Q (signal_6261) ) ;
    buf_clk cell_3731 ( .C (clk), .D (signal_6276), .Q (signal_6277) ) ;
    buf_clk cell_3747 ( .C (clk), .D (signal_6292), .Q (signal_6293) ) ;
    buf_clk cell_3763 ( .C (clk), .D (signal_6308), .Q (signal_6309) ) ;
    buf_clk cell_3779 ( .C (clk), .D (signal_6324), .Q (signal_6325) ) ;
    buf_clk cell_3795 ( .C (clk), .D (signal_6340), .Q (signal_6341) ) ;
    buf_clk cell_3811 ( .C (clk), .D (signal_6356), .Q (signal_6357) ) ;
    buf_clk cell_3827 ( .C (clk), .D (signal_6372), .Q (signal_6373) ) ;
    buf_clk cell_3843 ( .C (clk), .D (signal_6388), .Q (signal_6389) ) ;
    buf_clk cell_3859 ( .C (clk), .D (signal_6404), .Q (signal_6405) ) ;
    buf_clk cell_3875 ( .C (clk), .D (signal_6420), .Q (signal_6421) ) ;
    buf_clk cell_3891 ( .C (clk), .D (signal_6436), .Q (signal_6437) ) ;
    buf_clk cell_3907 ( .C (clk), .D (signal_6452), .Q (signal_6453) ) ;
    buf_clk cell_3923 ( .C (clk), .D (signal_6468), .Q (signal_6469) ) ;
    buf_clk cell_3939 ( .C (clk), .D (signal_6484), .Q (signal_6485) ) ;
    buf_clk cell_3955 ( .C (clk), .D (signal_6500), .Q (signal_6501) ) ;
    buf_clk cell_3971 ( .C (clk), .D (signal_6516), .Q (signal_6517) ) ;
    buf_clk cell_3987 ( .C (clk), .D (signal_6532), .Q (signal_6533) ) ;
    buf_clk cell_4003 ( .C (clk), .D (signal_6548), .Q (signal_6549) ) ;
    buf_clk cell_4019 ( .C (clk), .D (signal_6564), .Q (signal_6565) ) ;
    buf_clk cell_4035 ( .C (clk), .D (signal_6580), .Q (signal_6581) ) ;
    buf_clk cell_4051 ( .C (clk), .D (signal_6596), .Q (signal_6597) ) ;
    buf_clk cell_4067 ( .C (clk), .D (signal_6612), .Q (signal_6613) ) ;
    buf_clk cell_4083 ( .C (clk), .D (signal_6628), .Q (signal_6629) ) ;
    buf_clk cell_4099 ( .C (clk), .D (signal_6644), .Q (signal_6645) ) ;
    buf_clk cell_4115 ( .C (clk), .D (signal_6660), .Q (signal_6661) ) ;
    buf_clk cell_4131 ( .C (clk), .D (signal_6676), .Q (signal_6677) ) ;
    buf_clk cell_4147 ( .C (clk), .D (signal_6692), .Q (signal_6693) ) ;
    buf_clk cell_4163 ( .C (clk), .D (signal_6708), .Q (signal_6709) ) ;
    buf_clk cell_4179 ( .C (clk), .D (signal_6724), .Q (signal_6725) ) ;
    buf_clk cell_4195 ( .C (clk), .D (signal_6740), .Q (signal_6741) ) ;
    buf_clk cell_4211 ( .C (clk), .D (signal_6756), .Q (signal_6757) ) ;
    buf_clk cell_4227 ( .C (clk), .D (signal_6772), .Q (signal_6773) ) ;
    buf_clk cell_4243 ( .C (clk), .D (signal_6788), .Q (signal_6789) ) ;
    buf_clk cell_4259 ( .C (clk), .D (signal_6804), .Q (signal_6805) ) ;
    buf_clk cell_4275 ( .C (clk), .D (signal_6820), .Q (signal_6821) ) ;
    buf_clk cell_4291 ( .C (clk), .D (signal_6836), .Q (signal_6837) ) ;
    buf_clk cell_4307 ( .C (clk), .D (signal_6852), .Q (signal_6853) ) ;
    buf_clk cell_4323 ( .C (clk), .D (signal_6868), .Q (signal_6869) ) ;
    buf_clk cell_4339 ( .C (clk), .D (signal_6884), .Q (signal_6885) ) ;
    buf_clk cell_4355 ( .C (clk), .D (signal_6900), .Q (signal_6901) ) ;
    buf_clk cell_4371 ( .C (clk), .D (signal_6916), .Q (signal_6917) ) ;
    buf_clk cell_4387 ( .C (clk), .D (signal_6932), .Q (signal_6933) ) ;
    buf_clk cell_4403 ( .C (clk), .D (signal_6948), .Q (signal_6949) ) ;
    buf_clk cell_4417 ( .C (clk), .D (signal_6962), .Q (signal_6963) ) ;
    buf_clk cell_4431 ( .C (clk), .D (signal_6976), .Q (signal_6977) ) ;
    buf_clk cell_4447 ( .C (clk), .D (signal_6992), .Q (signal_6993) ) ;
    buf_clk cell_4463 ( .C (clk), .D (signal_7008), .Q (signal_7009) ) ;
    buf_clk cell_4479 ( .C (clk), .D (signal_7024), .Q (signal_7025) ) ;
    buf_clk cell_4495 ( .C (clk), .D (signal_7040), .Q (signal_7041) ) ;
    buf_clk cell_4511 ( .C (clk), .D (signal_7056), .Q (signal_7057) ) ;
    buf_clk cell_4527 ( .C (clk), .D (signal_7072), .Q (signal_7073) ) ;
    buf_clk cell_4543 ( .C (clk), .D (signal_7088), .Q (signal_7089) ) ;
    buf_clk cell_4559 ( .C (clk), .D (signal_7104), .Q (signal_7105) ) ;
    buf_clk cell_4575 ( .C (clk), .D (signal_7120), .Q (signal_7121) ) ;
    buf_clk cell_4591 ( .C (clk), .D (signal_7136), .Q (signal_7137) ) ;
    buf_clk cell_4607 ( .C (clk), .D (signal_7152), .Q (signal_7153) ) ;
    buf_clk cell_4623 ( .C (clk), .D (signal_7168), .Q (signal_7169) ) ;
    buf_clk cell_4639 ( .C (clk), .D (signal_7184), .Q (signal_7185) ) ;
    buf_clk cell_4655 ( .C (clk), .D (signal_7200), .Q (signal_7201) ) ;
    buf_clk cell_4671 ( .C (clk), .D (signal_7216), .Q (signal_7217) ) ;
    buf_clk cell_4687 ( .C (clk), .D (signal_7232), .Q (signal_7233) ) ;
    buf_clk cell_4703 ( .C (clk), .D (signal_7248), .Q (signal_7249) ) ;
    buf_clk cell_4719 ( .C (clk), .D (signal_7264), .Q (signal_7265) ) ;
    buf_clk cell_4735 ( .C (clk), .D (signal_7280), .Q (signal_7281) ) ;
    buf_clk cell_4751 ( .C (clk), .D (signal_7296), .Q (signal_7297) ) ;
    buf_clk cell_4767 ( .C (clk), .D (signal_7312), .Q (signal_7313) ) ;
    buf_clk cell_4783 ( .C (clk), .D (signal_7328), .Q (signal_7329) ) ;
    buf_clk cell_4799 ( .C (clk), .D (signal_7344), .Q (signal_7345) ) ;
    buf_clk cell_4815 ( .C (clk), .D (signal_7360), .Q (signal_7361) ) ;
    buf_clk cell_4831 ( .C (clk), .D (signal_7376), .Q (signal_7377) ) ;
    buf_clk cell_4847 ( .C (clk), .D (signal_7392), .Q (signal_7393) ) ;
    buf_clk cell_4863 ( .C (clk), .D (signal_7408), .Q (signal_7409) ) ;
    buf_clk cell_4879 ( .C (clk), .D (signal_7424), .Q (signal_7425) ) ;
    buf_clk cell_4895 ( .C (clk), .D (signal_7440), .Q (signal_7441) ) ;
    buf_clk cell_4911 ( .C (clk), .D (signal_7456), .Q (signal_7457) ) ;
    buf_clk cell_4927 ( .C (clk), .D (signal_7472), .Q (signal_7473) ) ;
    buf_clk cell_4943 ( .C (clk), .D (signal_7488), .Q (signal_7489) ) ;
    buf_clk cell_4959 ( .C (clk), .D (signal_7504), .Q (signal_7505) ) ;
    buf_clk cell_4975 ( .C (clk), .D (signal_7520), .Q (signal_7521) ) ;
    buf_clk cell_4991 ( .C (clk), .D (signal_7536), .Q (signal_7537) ) ;
    buf_clk cell_5007 ( .C (clk), .D (signal_7552), .Q (signal_7553) ) ;
    buf_clk cell_5023 ( .C (clk), .D (signal_7568), .Q (signal_7569) ) ;
    buf_clk cell_5039 ( .C (clk), .D (signal_7584), .Q (signal_7585) ) ;
    buf_clk cell_5055 ( .C (clk), .D (signal_7600), .Q (signal_7601) ) ;
    buf_clk cell_5071 ( .C (clk), .D (signal_7616), .Q (signal_7617) ) ;
    buf_clk cell_5087 ( .C (clk), .D (signal_7632), .Q (signal_7633) ) ;
    buf_clk cell_5103 ( .C (clk), .D (signal_7648), .Q (signal_7649) ) ;
    buf_clk cell_5119 ( .C (clk), .D (signal_7664), .Q (signal_7665) ) ;
    buf_clk cell_5135 ( .C (clk), .D (signal_7680), .Q (signal_7681) ) ;
    buf_clk cell_5151 ( .C (clk), .D (signal_7696), .Q (signal_7697) ) ;
    buf_clk cell_5167 ( .C (clk), .D (signal_7712), .Q (signal_7713) ) ;
    buf_clk cell_5183 ( .C (clk), .D (signal_7728), .Q (signal_7729) ) ;
    buf_clk cell_5199 ( .C (clk), .D (signal_7744), .Q (signal_7745) ) ;
    buf_clk cell_5215 ( .C (clk), .D (signal_7760), .Q (signal_7761) ) ;
    buf_clk cell_5231 ( .C (clk), .D (signal_7776), .Q (signal_7777) ) ;
    buf_clk cell_5247 ( .C (clk), .D (signal_7792), .Q (signal_7793) ) ;
    buf_clk cell_5263 ( .C (clk), .D (signal_7808), .Q (signal_7809) ) ;
    buf_clk cell_5279 ( .C (clk), .D (signal_7824), .Q (signal_7825) ) ;
    buf_clk cell_5295 ( .C (clk), .D (signal_7840), .Q (signal_7841) ) ;
    buf_clk cell_5311 ( .C (clk), .D (signal_7856), .Q (signal_7857) ) ;
    buf_clk cell_5327 ( .C (clk), .D (signal_7872), .Q (signal_7873) ) ;
    buf_clk cell_5343 ( .C (clk), .D (signal_7888), .Q (signal_7889) ) ;
    buf_clk cell_5359 ( .C (clk), .D (signal_7904), .Q (signal_7905) ) ;
    buf_clk cell_5375 ( .C (clk), .D (signal_7920), .Q (signal_7921) ) ;
    buf_clk cell_5391 ( .C (clk), .D (signal_7936), .Q (signal_7937) ) ;
    buf_clk cell_5407 ( .C (clk), .D (signal_7952), .Q (signal_7953) ) ;
    buf_clk cell_5423 ( .C (clk), .D (signal_7968), .Q (signal_7969) ) ;
    buf_clk cell_5439 ( .C (clk), .D (signal_7984), .Q (signal_7985) ) ;
    buf_clk cell_5455 ( .C (clk), .D (signal_8000), .Q (signal_8001) ) ;
    buf_clk cell_5471 ( .C (clk), .D (signal_8016), .Q (signal_8017) ) ;
    buf_clk cell_5487 ( .C (clk), .D (signal_8032), .Q (signal_8033) ) ;
    buf_clk cell_5503 ( .C (clk), .D (signal_8048), .Q (signal_8049) ) ;
    buf_clk cell_5519 ( .C (clk), .D (signal_8064), .Q (signal_8065) ) ;
    buf_clk cell_5535 ( .C (clk), .D (signal_8080), .Q (signal_8081) ) ;
    buf_clk cell_5551 ( .C (clk), .D (signal_8096), .Q (signal_8097) ) ;
    buf_clk cell_5567 ( .C (clk), .D (signal_8112), .Q (signal_8113) ) ;
    buf_clk cell_5583 ( .C (clk), .D (signal_8128), .Q (signal_8129) ) ;
    buf_clk cell_5599 ( .C (clk), .D (signal_8144), .Q (signal_8145) ) ;
    buf_clk cell_5615 ( .C (clk), .D (signal_8160), .Q (signal_8161) ) ;
    buf_clk cell_5631 ( .C (clk), .D (signal_8176), .Q (signal_8177) ) ;
    buf_clk cell_5647 ( .C (clk), .D (signal_8192), .Q (signal_8193) ) ;
    buf_clk cell_5663 ( .C (clk), .D (signal_8208), .Q (signal_8209) ) ;
    buf_clk cell_5679 ( .C (clk), .D (signal_8224), .Q (signal_8225) ) ;
    buf_clk cell_5695 ( .C (clk), .D (signal_8240), .Q (signal_8241) ) ;
    buf_clk cell_5711 ( .C (clk), .D (signal_8256), .Q (signal_8257) ) ;
    buf_clk cell_5727 ( .C (clk), .D (signal_8272), .Q (signal_8273) ) ;
    buf_clk cell_5743 ( .C (clk), .D (signal_8288), .Q (signal_8289) ) ;
    buf_clk cell_5759 ( .C (clk), .D (signal_8304), .Q (signal_8305) ) ;
    buf_clk cell_5775 ( .C (clk), .D (signal_8320), .Q (signal_8321) ) ;
    buf_clk cell_5791 ( .C (clk), .D (signal_8336), .Q (signal_8337) ) ;
    buf_clk cell_5807 ( .C (clk), .D (signal_8352), .Q (signal_8353) ) ;
    buf_clk cell_5823 ( .C (clk), .D (signal_8368), .Q (signal_8369) ) ;
    buf_clk cell_5839 ( .C (clk), .D (signal_8384), .Q (signal_8385) ) ;
    buf_clk cell_5855 ( .C (clk), .D (signal_8400), .Q (signal_8401) ) ;
    buf_clk cell_5871 ( .C (clk), .D (signal_8416), .Q (signal_8417) ) ;
    buf_clk cell_5887 ( .C (clk), .D (signal_8432), .Q (signal_8433) ) ;
    buf_clk cell_5903 ( .C (clk), .D (signal_8448), .Q (signal_8449) ) ;
    buf_clk cell_5919 ( .C (clk), .D (signal_8464), .Q (signal_8465) ) ;
    buf_clk cell_5935 ( .C (clk), .D (signal_8480), .Q (signal_8481) ) ;
    buf_clk cell_5951 ( .C (clk), .D (signal_8496), .Q (signal_8497) ) ;
    buf_clk cell_5967 ( .C (clk), .D (signal_8512), .Q (signal_8513) ) ;
    buf_clk cell_5983 ( .C (clk), .D (signal_8528), .Q (signal_8529) ) ;
    buf_clk cell_5999 ( .C (clk), .D (signal_8544), .Q (signal_8545) ) ;
    buf_clk cell_6015 ( .C (clk), .D (signal_8560), .Q (signal_8561) ) ;
    buf_clk cell_6031 ( .C (clk), .D (signal_8576), .Q (signal_8577) ) ;
    buf_clk cell_6047 ( .C (clk), .D (signal_8592), .Q (signal_8593) ) ;
    buf_clk cell_6063 ( .C (clk), .D (signal_8608), .Q (signal_8609) ) ;
    buf_clk cell_6079 ( .C (clk), .D (signal_8624), .Q (signal_8625) ) ;
    buf_clk cell_6095 ( .C (clk), .D (signal_8640), .Q (signal_8641) ) ;
    buf_clk cell_6111 ( .C (clk), .D (signal_8656), .Q (signal_8657) ) ;
    buf_clk cell_6127 ( .C (clk), .D (signal_8672), .Q (signal_8673) ) ;
    buf_clk cell_6143 ( .C (clk), .D (signal_8688), .Q (signal_8689) ) ;
    buf_clk cell_6159 ( .C (clk), .D (signal_8704), .Q (signal_8705) ) ;
    buf_clk cell_6175 ( .C (clk), .D (signal_8720), .Q (signal_8721) ) ;
    buf_clk cell_6191 ( .C (clk), .D (signal_8736), .Q (signal_8737) ) ;
    buf_clk cell_6207 ( .C (clk), .D (signal_8752), .Q (signal_8753) ) ;
    buf_clk cell_6223 ( .C (clk), .D (signal_8768), .Q (signal_8769) ) ;
    buf_clk cell_6239 ( .C (clk), .D (signal_8784), .Q (signal_8785) ) ;
    buf_clk cell_6255 ( .C (clk), .D (signal_8800), .Q (signal_8801) ) ;
    buf_clk cell_6271 ( .C (clk), .D (signal_8816), .Q (signal_8817) ) ;
    buf_clk cell_6287 ( .C (clk), .D (signal_8832), .Q (signal_8833) ) ;
    buf_clk cell_6303 ( .C (clk), .D (signal_8848), .Q (signal_8849) ) ;
    buf_clk cell_6319 ( .C (clk), .D (signal_8864), .Q (signal_8865) ) ;
    buf_clk cell_6335 ( .C (clk), .D (signal_8880), .Q (signal_8881) ) ;
    buf_clk cell_6351 ( .C (clk), .D (signal_8896), .Q (signal_8897) ) ;
    buf_clk cell_6367 ( .C (clk), .D (signal_8912), .Q (signal_8913) ) ;
    buf_clk cell_6383 ( .C (clk), .D (signal_8928), .Q (signal_8929) ) ;
    buf_clk cell_6399 ( .C (clk), .D (signal_8944), .Q (signal_8945) ) ;
    buf_clk cell_6415 ( .C (clk), .D (signal_8960), .Q (signal_8961) ) ;
    buf_clk cell_6431 ( .C (clk), .D (signal_8976), .Q (signal_8977) ) ;
    buf_clk cell_6447 ( .C (clk), .D (signal_8992), .Q (signal_8993) ) ;
    buf_clk cell_6463 ( .C (clk), .D (signal_9008), .Q (signal_9009) ) ;
    buf_clk cell_6479 ( .C (clk), .D (signal_9024), .Q (signal_9025) ) ;
    buf_clk cell_6495 ( .C (clk), .D (signal_9040), .Q (signal_9041) ) ;
    buf_clk cell_6511 ( .C (clk), .D (signal_9056), .Q (signal_9057) ) ;
    buf_clk cell_6527 ( .C (clk), .D (signal_9072), .Q (signal_9073) ) ;
    buf_clk cell_6543 ( .C (clk), .D (signal_9088), .Q (signal_9089) ) ;
    buf_clk cell_6559 ( .C (clk), .D (signal_9104), .Q (signal_9105) ) ;
    buf_clk cell_6575 ( .C (clk), .D (signal_9120), .Q (signal_9121) ) ;
    buf_clk cell_6591 ( .C (clk), .D (signal_9136), .Q (signal_9137) ) ;
    buf_clk cell_6607 ( .C (clk), .D (signal_9152), .Q (signal_9153) ) ;
    buf_clk cell_6623 ( .C (clk), .D (signal_9168), .Q (signal_9169) ) ;
    buf_clk cell_6639 ( .C (clk), .D (signal_9184), .Q (signal_9185) ) ;
    buf_clk cell_6655 ( .C (clk), .D (signal_9200), .Q (signal_9201) ) ;
    buf_clk cell_6671 ( .C (clk), .D (signal_9216), .Q (signal_9217) ) ;
    buf_clk cell_6687 ( .C (clk), .D (signal_9232), .Q (signal_9233) ) ;
    buf_clk cell_6703 ( .C (clk), .D (signal_9248), .Q (signal_9249) ) ;
    buf_clk cell_6719 ( .C (clk), .D (signal_9264), .Q (signal_9265) ) ;
    buf_clk cell_6735 ( .C (clk), .D (signal_9280), .Q (signal_9281) ) ;
    buf_clk cell_6751 ( .C (clk), .D (signal_9296), .Q (signal_9297) ) ;
    buf_clk cell_6767 ( .C (clk), .D (signal_9312), .Q (signal_9313) ) ;
    buf_clk cell_6783 ( .C (clk), .D (signal_9328), .Q (signal_9329) ) ;
    buf_clk cell_6799 ( .C (clk), .D (signal_9344), .Q (signal_9345) ) ;
    buf_clk cell_6815 ( .C (clk), .D (signal_9360), .Q (signal_9361) ) ;
    buf_clk cell_6831 ( .C (clk), .D (signal_9376), .Q (signal_9377) ) ;
    buf_clk cell_6847 ( .C (clk), .D (signal_9392), .Q (signal_9393) ) ;
    buf_clk cell_6863 ( .C (clk), .D (signal_9408), .Q (signal_9409) ) ;
    buf_clk cell_6879 ( .C (clk), .D (signal_9424), .Q (signal_9425) ) ;
    buf_clk cell_6895 ( .C (clk), .D (signal_9440), .Q (signal_9441) ) ;
    buf_clk cell_6911 ( .C (clk), .D (signal_9456), .Q (signal_9457) ) ;
    buf_clk cell_6927 ( .C (clk), .D (signal_9472), .Q (signal_9473) ) ;
    buf_clk cell_6943 ( .C (clk), .D (signal_9488), .Q (signal_9489) ) ;
    buf_clk cell_6959 ( .C (clk), .D (signal_9504), .Q (signal_9505) ) ;
    buf_clk cell_6975 ( .C (clk), .D (signal_9520), .Q (signal_9521) ) ;
    buf_clk cell_6991 ( .C (clk), .D (signal_9536), .Q (signal_9537) ) ;
    buf_clk cell_7007 ( .C (clk), .D (signal_9552), .Q (signal_9553) ) ;
    buf_clk cell_7023 ( .C (clk), .D (signal_9568), .Q (signal_9569) ) ;
    buf_clk cell_7039 ( .C (clk), .D (signal_9584), .Q (signal_9585) ) ;
    buf_clk cell_7055 ( .C (clk), .D (signal_9600), .Q (signal_9601) ) ;
    buf_clk cell_7071 ( .C (clk), .D (signal_9616), .Q (signal_9617) ) ;
    buf_clk cell_7087 ( .C (clk), .D (signal_9632), .Q (signal_9633) ) ;
    buf_clk cell_7103 ( .C (clk), .D (signal_9648), .Q (signal_9649) ) ;
    buf_clk cell_7119 ( .C (clk), .D (signal_9664), .Q (signal_9665) ) ;
    buf_clk cell_7135 ( .C (clk), .D (signal_9680), .Q (signal_9681) ) ;
    buf_clk cell_7151 ( .C (clk), .D (signal_9696), .Q (signal_9697) ) ;
    buf_clk cell_7167 ( .C (clk), .D (signal_9712), .Q (signal_9713) ) ;
    buf_clk cell_7183 ( .C (clk), .D (signal_9728), .Q (signal_9729) ) ;
    buf_clk cell_7199 ( .C (clk), .D (signal_9744), .Q (signal_9745) ) ;
    buf_clk cell_7215 ( .C (clk), .D (signal_9760), .Q (signal_9761) ) ;
    buf_clk cell_7231 ( .C (clk), .D (signal_9776), .Q (signal_9777) ) ;
    buf_clk cell_7247 ( .C (clk), .D (signal_9792), .Q (signal_9793) ) ;
    buf_clk cell_7263 ( .C (clk), .D (signal_9808), .Q (signal_9809) ) ;
    buf_clk cell_7279 ( .C (clk), .D (signal_9824), .Q (signal_9825) ) ;
    buf_clk cell_7295 ( .C (clk), .D (signal_9840), .Q (signal_9841) ) ;
    buf_clk cell_7311 ( .C (clk), .D (signal_9856), .Q (signal_9857) ) ;
    buf_clk cell_7327 ( .C (clk), .D (signal_9872), .Q (signal_9873) ) ;
    buf_clk cell_7343 ( .C (clk), .D (signal_9888), .Q (signal_9889) ) ;
    buf_clk cell_7359 ( .C (clk), .D (signal_9904), .Q (signal_9905) ) ;
    buf_clk cell_7375 ( .C (clk), .D (signal_9920), .Q (signal_9921) ) ;
    buf_clk cell_7391 ( .C (clk), .D (signal_9936), .Q (signal_9937) ) ;
    buf_clk cell_7407 ( .C (clk), .D (signal_9952), .Q (signal_9953) ) ;
    buf_clk cell_7423 ( .C (clk), .D (signal_9968), .Q (signal_9969) ) ;
    buf_clk cell_7439 ( .C (clk), .D (signal_9984), .Q (signal_9985) ) ;
    buf_clk cell_7455 ( .C (clk), .D (signal_10000), .Q (signal_10001) ) ;
    buf_clk cell_7471 ( .C (clk), .D (signal_10016), .Q (signal_10017) ) ;
    buf_clk cell_7487 ( .C (clk), .D (signal_10032), .Q (signal_10033) ) ;
    buf_clk cell_7503 ( .C (clk), .D (signal_10048), .Q (signal_10049) ) ;
    buf_clk cell_7519 ( .C (clk), .D (signal_10064), .Q (signal_10065) ) ;
    buf_clk cell_7535 ( .C (clk), .D (signal_10080), .Q (signal_10081) ) ;
    buf_clk cell_7551 ( .C (clk), .D (signal_10096), .Q (signal_10097) ) ;
    buf_clk cell_7567 ( .C (clk), .D (signal_10112), .Q (signal_10113) ) ;
    buf_clk cell_7583 ( .C (clk), .D (signal_10128), .Q (signal_10129) ) ;
    buf_clk cell_7599 ( .C (clk), .D (signal_10144), .Q (signal_10145) ) ;
    buf_clk cell_7615 ( .C (clk), .D (signal_10160), .Q (signal_10161) ) ;
    buf_clk cell_7631 ( .C (clk), .D (signal_10176), .Q (signal_10177) ) ;
    buf_clk cell_7647 ( .C (clk), .D (signal_10192), .Q (signal_10193) ) ;
    buf_clk cell_7663 ( .C (clk), .D (signal_10208), .Q (signal_10209) ) ;
    buf_clk cell_7679 ( .C (clk), .D (signal_10224), .Q (signal_10225) ) ;
    buf_clk cell_7695 ( .C (clk), .D (signal_10240), .Q (signal_10241) ) ;
    buf_clk cell_7711 ( .C (clk), .D (signal_10256), .Q (signal_10257) ) ;
    buf_clk cell_7727 ( .C (clk), .D (signal_10272), .Q (signal_10273) ) ;
    buf_clk cell_7743 ( .C (clk), .D (signal_10288), .Q (signal_10289) ) ;
    buf_clk cell_7759 ( .C (clk), .D (signal_10304), .Q (signal_10305) ) ;
    buf_clk cell_7775 ( .C (clk), .D (signal_10320), .Q (signal_10321) ) ;
    buf_clk cell_7791 ( .C (clk), .D (signal_10336), .Q (signal_10337) ) ;
    buf_clk cell_7807 ( .C (clk), .D (signal_10352), .Q (signal_10353) ) ;
    buf_clk cell_7823 ( .C (clk), .D (signal_10368), .Q (signal_10369) ) ;
    buf_clk cell_7839 ( .C (clk), .D (signal_10384), .Q (signal_10385) ) ;
    buf_clk cell_7855 ( .C (clk), .D (signal_10400), .Q (signal_10401) ) ;
    buf_clk cell_7871 ( .C (clk), .D (signal_10416), .Q (signal_10417) ) ;
    buf_clk cell_7887 ( .C (clk), .D (signal_10432), .Q (signal_10433) ) ;
    buf_clk cell_7903 ( .C (clk), .D (signal_10448), .Q (signal_10449) ) ;
    buf_clk cell_7919 ( .C (clk), .D (signal_10464), .Q (signal_10465) ) ;
    buf_clk cell_7935 ( .C (clk), .D (signal_10480), .Q (signal_10481) ) ;
    buf_clk cell_7951 ( .C (clk), .D (signal_10496), .Q (signal_10497) ) ;
    buf_clk cell_7967 ( .C (clk), .D (signal_10512), .Q (signal_10513) ) ;
    buf_clk cell_7983 ( .C (clk), .D (signal_10528), .Q (signal_10529) ) ;
    buf_clk cell_7999 ( .C (clk), .D (signal_10544), .Q (signal_10545) ) ;
    buf_clk cell_8015 ( .C (clk), .D (signal_10560), .Q (signal_10561) ) ;
    buf_clk cell_8031 ( .C (clk), .D (signal_10576), .Q (signal_10577) ) ;
    buf_clk cell_8047 ( .C (clk), .D (signal_10592), .Q (signal_10593) ) ;
    buf_clk cell_8063 ( .C (clk), .D (signal_10608), .Q (signal_10609) ) ;
    buf_clk cell_8079 ( .C (clk), .D (signal_10624), .Q (signal_10625) ) ;
    buf_clk cell_8095 ( .C (clk), .D (signal_10640), .Q (signal_10641) ) ;
    buf_clk cell_8111 ( .C (clk), .D (signal_10656), .Q (signal_10657) ) ;
    buf_clk cell_8127 ( .C (clk), .D (signal_10672), .Q (signal_10673) ) ;
    buf_clk cell_8143 ( .C (clk), .D (signal_10688), .Q (signal_10689) ) ;
    buf_clk cell_8159 ( .C (clk), .D (signal_10704), .Q (signal_10705) ) ;
    buf_clk cell_8175 ( .C (clk), .D (signal_10720), .Q (signal_10721) ) ;
    buf_clk cell_8191 ( .C (clk), .D (signal_10736), .Q (signal_10737) ) ;
    buf_clk cell_8207 ( .C (clk), .D (signal_10752), .Q (signal_10753) ) ;
    buf_clk cell_8223 ( .C (clk), .D (signal_10768), .Q (signal_10769) ) ;
    buf_clk cell_8239 ( .C (clk), .D (signal_10784), .Q (signal_10785) ) ;
    buf_clk cell_8255 ( .C (clk), .D (signal_10800), .Q (signal_10801) ) ;
    buf_clk cell_8271 ( .C (clk), .D (signal_10816), .Q (signal_10817) ) ;
    buf_clk cell_8287 ( .C (clk), .D (signal_10832), .Q (signal_10833) ) ;
    buf_clk cell_8303 ( .C (clk), .D (signal_10848), .Q (signal_10849) ) ;
    buf_clk cell_8319 ( .C (clk), .D (signal_10864), .Q (signal_10865) ) ;
    buf_clk cell_8335 ( .C (clk), .D (signal_10880), .Q (signal_10881) ) ;
    buf_clk cell_8351 ( .C (clk), .D (signal_10896), .Q (signal_10897) ) ;
    buf_clk cell_8367 ( .C (clk), .D (signal_10912), .Q (signal_10913) ) ;
    buf_clk cell_8383 ( .C (clk), .D (signal_10928), .Q (signal_10929) ) ;
    buf_clk cell_8399 ( .C (clk), .D (signal_10944), .Q (signal_10945) ) ;
    buf_clk cell_8415 ( .C (clk), .D (signal_10960), .Q (signal_10961) ) ;
    buf_clk cell_8431 ( .C (clk), .D (signal_10976), .Q (signal_10977) ) ;
    buf_clk cell_8447 ( .C (clk), .D (signal_10992), .Q (signal_10993) ) ;
    buf_clk cell_8463 ( .C (clk), .D (signal_11008), .Q (signal_11009) ) ;
    buf_clk cell_8479 ( .C (clk), .D (signal_11024), .Q (signal_11025) ) ;
    buf_clk cell_8495 ( .C (clk), .D (signal_11040), .Q (signal_11041) ) ;
    buf_clk cell_8511 ( .C (clk), .D (signal_11056), .Q (signal_11057) ) ;
    buf_clk cell_8527 ( .C (clk), .D (signal_11072), .Q (signal_11073) ) ;
    buf_clk cell_8543 ( .C (clk), .D (signal_11088), .Q (signal_11089) ) ;
    buf_clk cell_8559 ( .C (clk), .D (signal_11104), .Q (signal_11105) ) ;
    buf_clk cell_8575 ( .C (clk), .D (signal_11120), .Q (signal_11121) ) ;
    buf_clk cell_8591 ( .C (clk), .D (signal_11136), .Q (signal_11137) ) ;
    buf_clk cell_8607 ( .C (clk), .D (signal_11152), .Q (signal_11153) ) ;
    buf_clk cell_8623 ( .C (clk), .D (signal_11168), .Q (signal_11169) ) ;
    buf_clk cell_8639 ( .C (clk), .D (signal_11184), .Q (signal_11185) ) ;
    buf_clk cell_8655 ( .C (clk), .D (signal_11200), .Q (signal_11201) ) ;
    buf_clk cell_8671 ( .C (clk), .D (signal_11216), .Q (signal_11217) ) ;
    buf_clk cell_8687 ( .C (clk), .D (signal_11232), .Q (signal_11233) ) ;
    buf_clk cell_8703 ( .C (clk), .D (signal_11248), .Q (signal_11249) ) ;
    buf_clk cell_8719 ( .C (clk), .D (signal_11264), .Q (signal_11265) ) ;
    buf_clk cell_8735 ( .C (clk), .D (signal_11280), .Q (signal_11281) ) ;
    buf_clk cell_8751 ( .C (clk), .D (signal_11296), .Q (signal_11297) ) ;
    buf_clk cell_8767 ( .C (clk), .D (signal_11312), .Q (signal_11313) ) ;
    buf_clk cell_8783 ( .C (clk), .D (signal_11328), .Q (signal_11329) ) ;
    buf_clk cell_8799 ( .C (clk), .D (signal_11344), .Q (signal_11345) ) ;
    buf_clk cell_8815 ( .C (clk), .D (signal_11360), .Q (signal_11361) ) ;
    buf_clk cell_8831 ( .C (clk), .D (signal_11376), .Q (signal_11377) ) ;
    buf_clk cell_8847 ( .C (clk), .D (signal_11392), .Q (signal_11393) ) ;
    buf_clk cell_8863 ( .C (clk), .D (signal_11408), .Q (signal_11409) ) ;
    buf_clk cell_8879 ( .C (clk), .D (signal_11424), .Q (signal_11425) ) ;
    buf_clk cell_8895 ( .C (clk), .D (signal_11440), .Q (signal_11441) ) ;
    buf_clk cell_8911 ( .C (clk), .D (signal_11456), .Q (signal_11457) ) ;
    buf_clk cell_8927 ( .C (clk), .D (signal_11472), .Q (signal_11473) ) ;
    buf_clk cell_8943 ( .C (clk), .D (signal_11488), .Q (signal_11489) ) ;
    buf_clk cell_8959 ( .C (clk), .D (signal_11504), .Q (signal_11505) ) ;
    buf_clk cell_8975 ( .C (clk), .D (signal_11520), .Q (signal_11521) ) ;
    buf_clk cell_8991 ( .C (clk), .D (signal_11536), .Q (signal_11537) ) ;
    buf_clk cell_9007 ( .C (clk), .D (signal_11552), .Q (signal_11553) ) ;
    buf_clk cell_9023 ( .C (clk), .D (signal_11568), .Q (signal_11569) ) ;
    buf_clk cell_9039 ( .C (clk), .D (signal_11584), .Q (signal_11585) ) ;
    buf_clk cell_9055 ( .C (clk), .D (signal_11600), .Q (signal_11601) ) ;
    buf_clk cell_9071 ( .C (clk), .D (signal_11616), .Q (signal_11617) ) ;
    buf_clk cell_9087 ( .C (clk), .D (signal_11632), .Q (signal_11633) ) ;
    buf_clk cell_9103 ( .C (clk), .D (signal_11648), .Q (signal_11649) ) ;
    buf_clk cell_9119 ( .C (clk), .D (signal_11664), .Q (signal_11665) ) ;
    buf_clk cell_9135 ( .C (clk), .D (signal_11680), .Q (signal_11681) ) ;
    buf_clk cell_9151 ( .C (clk), .D (signal_11696), .Q (signal_11697) ) ;
    buf_clk cell_9167 ( .C (clk), .D (signal_11712), .Q (signal_11713) ) ;
    buf_clk cell_9183 ( .C (clk), .D (signal_11728), .Q (signal_11729) ) ;
    buf_clk cell_9199 ( .C (clk), .D (signal_11744), .Q (signal_11745) ) ;
    buf_clk cell_9215 ( .C (clk), .D (signal_11760), .Q (signal_11761) ) ;
    buf_clk cell_9231 ( .C (clk), .D (signal_11776), .Q (signal_11777) ) ;
    buf_clk cell_9247 ( .C (clk), .D (signal_11792), .Q (signal_11793) ) ;
    buf_clk cell_9263 ( .C (clk), .D (signal_11808), .Q (signal_11809) ) ;
    buf_clk cell_9279 ( .C (clk), .D (signal_11824), .Q (signal_11825) ) ;
    buf_clk cell_9295 ( .C (clk), .D (signal_11840), .Q (signal_11841) ) ;
    buf_clk cell_9311 ( .C (clk), .D (signal_11856), .Q (signal_11857) ) ;
    buf_clk cell_9327 ( .C (clk), .D (signal_11872), .Q (signal_11873) ) ;
    buf_clk cell_9343 ( .C (clk), .D (signal_11888), .Q (signal_11889) ) ;
    buf_clk cell_9359 ( .C (clk), .D (signal_11904), .Q (signal_11905) ) ;
    buf_clk cell_9375 ( .C (clk), .D (signal_11920), .Q (signal_11921) ) ;
    buf_clk cell_9391 ( .C (clk), .D (signal_11936), .Q (signal_11937) ) ;
    buf_clk cell_9407 ( .C (clk), .D (signal_11952), .Q (signal_11953) ) ;
    buf_clk cell_9423 ( .C (clk), .D (signal_11968), .Q (signal_11969) ) ;
    buf_clk cell_9439 ( .C (clk), .D (signal_11984), .Q (signal_11985) ) ;
    buf_clk cell_9455 ( .C (clk), .D (signal_12000), .Q (signal_12001) ) ;
    buf_clk cell_9471 ( .C (clk), .D (signal_12016), .Q (signal_12017) ) ;
    buf_clk cell_9487 ( .C (clk), .D (signal_12032), .Q (signal_12033) ) ;
    buf_clk cell_9503 ( .C (clk), .D (signal_12048), .Q (signal_12049) ) ;
    buf_clk cell_9519 ( .C (clk), .D (signal_12064), .Q (signal_12065) ) ;
    buf_clk cell_9535 ( .C (clk), .D (signal_12080), .Q (signal_12081) ) ;
    buf_clk cell_9551 ( .C (clk), .D (signal_12096), .Q (signal_12097) ) ;
    buf_clk cell_9567 ( .C (clk), .D (signal_12112), .Q (signal_12113) ) ;
    buf_clk cell_9583 ( .C (clk), .D (signal_12128), .Q (signal_12129) ) ;
    buf_clk cell_9599 ( .C (clk), .D (signal_12144), .Q (signal_12145) ) ;
    buf_clk cell_9615 ( .C (clk), .D (signal_12160), .Q (signal_12161) ) ;
    buf_clk cell_9631 ( .C (clk), .D (signal_12176), .Q (signal_12177) ) ;
    buf_clk cell_9647 ( .C (clk), .D (signal_12192), .Q (signal_12193) ) ;
    buf_clk cell_9663 ( .C (clk), .D (signal_12208), .Q (signal_12209) ) ;
    buf_clk cell_9679 ( .C (clk), .D (signal_12224), .Q (signal_12225) ) ;
    buf_clk cell_9695 ( .C (clk), .D (signal_12240), .Q (signal_12241) ) ;
    buf_clk cell_9711 ( .C (clk), .D (signal_12256), .Q (signal_12257) ) ;
    buf_clk cell_9727 ( .C (clk), .D (signal_12272), .Q (signal_12273) ) ;
    buf_clk cell_9743 ( .C (clk), .D (signal_12288), .Q (signal_12289) ) ;
    buf_clk cell_9759 ( .C (clk), .D (signal_12304), .Q (signal_12305) ) ;
    buf_clk cell_9775 ( .C (clk), .D (signal_12320), .Q (signal_12321) ) ;
    buf_clk cell_9791 ( .C (clk), .D (signal_12336), .Q (signal_12337) ) ;
    buf_clk cell_9807 ( .C (clk), .D (signal_12352), .Q (signal_12353) ) ;
    buf_clk cell_9823 ( .C (clk), .D (signal_12368), .Q (signal_12369) ) ;
    buf_clk cell_9839 ( .C (clk), .D (signal_12384), .Q (signal_12385) ) ;
    buf_clk cell_9855 ( .C (clk), .D (signal_12400), .Q (signal_12401) ) ;
    buf_clk cell_9871 ( .C (clk), .D (signal_12416), .Q (signal_12417) ) ;
    buf_clk cell_9887 ( .C (clk), .D (signal_12432), .Q (signal_12433) ) ;
    buf_clk cell_9903 ( .C (clk), .D (signal_12448), .Q (signal_12449) ) ;
    buf_clk cell_9919 ( .C (clk), .D (signal_12464), .Q (signal_12465) ) ;
    buf_clk cell_9935 ( .C (clk), .D (signal_12480), .Q (signal_12481) ) ;
    buf_clk cell_9951 ( .C (clk), .D (signal_12496), .Q (signal_12497) ) ;
    buf_clk cell_9967 ( .C (clk), .D (signal_12512), .Q (signal_12513) ) ;
    buf_clk cell_9983 ( .C (clk), .D (signal_12528), .Q (signal_12529) ) ;
    buf_clk cell_9999 ( .C (clk), .D (signal_12544), .Q (signal_12545) ) ;
    buf_clk cell_10015 ( .C (clk), .D (signal_12560), .Q (signal_12561) ) ;
    buf_clk cell_10031 ( .C (clk), .D (signal_12576), .Q (signal_12577) ) ;
    buf_clk cell_10047 ( .C (clk), .D (signal_12592), .Q (signal_12593) ) ;
    buf_clk cell_10063 ( .C (clk), .D (signal_12608), .Q (signal_12609) ) ;
    buf_clk cell_10079 ( .C (clk), .D (signal_12624), .Q (signal_12625) ) ;
    buf_clk cell_10095 ( .C (clk), .D (signal_12640), .Q (signal_12641) ) ;
    buf_clk cell_10111 ( .C (clk), .D (signal_12656), .Q (signal_12657) ) ;
    buf_clk cell_10127 ( .C (clk), .D (signal_12672), .Q (signal_12673) ) ;
    buf_clk cell_10143 ( .C (clk), .D (signal_12688), .Q (signal_12689) ) ;
    buf_clk cell_10159 ( .C (clk), .D (signal_12704), .Q (signal_12705) ) ;
    buf_clk cell_10175 ( .C (clk), .D (signal_12720), .Q (signal_12721) ) ;
    buf_clk cell_10191 ( .C (clk), .D (signal_12736), .Q (signal_12737) ) ;
    buf_clk cell_10207 ( .C (clk), .D (signal_12752), .Q (signal_12753) ) ;
    buf_clk cell_10223 ( .C (clk), .D (signal_12768), .Q (signal_12769) ) ;
    buf_clk cell_10239 ( .C (clk), .D (signal_12784), .Q (signal_12785) ) ;
    buf_clk cell_10255 ( .C (clk), .D (signal_12800), .Q (signal_12801) ) ;
    buf_clk cell_10271 ( .C (clk), .D (signal_12816), .Q (signal_12817) ) ;
    buf_clk cell_10287 ( .C (clk), .D (signal_12832), .Q (signal_12833) ) ;
    buf_clk cell_10303 ( .C (clk), .D (signal_12848), .Q (signal_12849) ) ;
    buf_clk cell_10319 ( .C (clk), .D (signal_12864), .Q (signal_12865) ) ;
    buf_clk cell_10335 ( .C (clk), .D (signal_12880), .Q (signal_12881) ) ;
    buf_clk cell_10351 ( .C (clk), .D (signal_12896), .Q (signal_12897) ) ;
    buf_clk cell_10367 ( .C (clk), .D (signal_12912), .Q (signal_12913) ) ;
    buf_clk cell_10383 ( .C (clk), .D (signal_12928), .Q (signal_12929) ) ;
    buf_clk cell_10399 ( .C (clk), .D (signal_12944), .Q (signal_12945) ) ;
    buf_clk cell_10415 ( .C (clk), .D (signal_12960), .Q (signal_12961) ) ;
    buf_clk cell_10431 ( .C (clk), .D (signal_12976), .Q (signal_12977) ) ;
    buf_clk cell_10447 ( .C (clk), .D (signal_12992), .Q (signal_12993) ) ;
    buf_clk cell_10463 ( .C (clk), .D (signal_13008), .Q (signal_13009) ) ;
    buf_clk cell_10479 ( .C (clk), .D (signal_13024), .Q (signal_13025) ) ;
    buf_clk cell_10495 ( .C (clk), .D (signal_13040), .Q (signal_13041) ) ;
    buf_clk cell_10511 ( .C (clk), .D (signal_13056), .Q (signal_13057) ) ;
    buf_clk cell_10527 ( .C (clk), .D (signal_13072), .Q (signal_13073) ) ;
    buf_clk cell_10543 ( .C (clk), .D (signal_13088), .Q (signal_13089) ) ;
    buf_clk cell_10559 ( .C (clk), .D (signal_13104), .Q (signal_13105) ) ;
    buf_clk cell_10575 ( .C (clk), .D (signal_13120), .Q (signal_13121) ) ;
    buf_clk cell_10591 ( .C (clk), .D (signal_13136), .Q (signal_13137) ) ;
    buf_clk cell_10607 ( .C (clk), .D (signal_13152), .Q (signal_13153) ) ;
    buf_clk cell_10623 ( .C (clk), .D (signal_13168), .Q (signal_13169) ) ;
    buf_clk cell_10639 ( .C (clk), .D (signal_13184), .Q (signal_13185) ) ;
    buf_clk cell_10655 ( .C (clk), .D (signal_13200), .Q (signal_13201) ) ;
    buf_clk cell_10671 ( .C (clk), .D (signal_13216), .Q (signal_13217) ) ;
    buf_clk cell_10687 ( .C (clk), .D (signal_13232), .Q (signal_13233) ) ;
    buf_clk cell_10703 ( .C (clk), .D (signal_13248), .Q (signal_13249) ) ;
    buf_clk cell_10719 ( .C (clk), .D (signal_13264), .Q (signal_13265) ) ;
    buf_clk cell_10735 ( .C (clk), .D (signal_13280), .Q (signal_13281) ) ;
    buf_clk cell_10751 ( .C (clk), .D (signal_13296), .Q (signal_13297) ) ;
    buf_clk cell_10767 ( .C (clk), .D (signal_13312), .Q (signal_13313) ) ;
    buf_clk cell_10783 ( .C (clk), .D (signal_13328), .Q (signal_13329) ) ;
    buf_clk cell_10799 ( .C (clk), .D (signal_13344), .Q (signal_13345) ) ;
    buf_clk cell_10815 ( .C (clk), .D (signal_13360), .Q (signal_13361) ) ;
    buf_clk cell_10831 ( .C (clk), .D (signal_13376), .Q (signal_13377) ) ;
    buf_clk cell_10847 ( .C (clk), .D (signal_13392), .Q (signal_13393) ) ;
    buf_clk cell_10863 ( .C (clk), .D (signal_13408), .Q (signal_13409) ) ;
    buf_clk cell_10879 ( .C (clk), .D (signal_13424), .Q (signal_13425) ) ;
    buf_clk cell_10895 ( .C (clk), .D (signal_13440), .Q (signal_13441) ) ;
    buf_clk cell_10911 ( .C (clk), .D (signal_13456), .Q (signal_13457) ) ;
    buf_clk cell_10927 ( .C (clk), .D (signal_13472), .Q (signal_13473) ) ;
    buf_clk cell_10943 ( .C (clk), .D (signal_13488), .Q (signal_13489) ) ;
    buf_clk cell_10959 ( .C (clk), .D (signal_13504), .Q (signal_13505) ) ;
    buf_clk cell_10975 ( .C (clk), .D (signal_13520), .Q (signal_13521) ) ;
    buf_clk cell_10991 ( .C (clk), .D (signal_13536), .Q (signal_13537) ) ;
    buf_clk cell_11007 ( .C (clk), .D (signal_13552), .Q (signal_13553) ) ;
    buf_clk cell_11023 ( .C (clk), .D (signal_13568), .Q (signal_13569) ) ;
    buf_clk cell_11039 ( .C (clk), .D (signal_13584), .Q (signal_13585) ) ;
    buf_clk cell_11055 ( .C (clk), .D (signal_13600), .Q (signal_13601) ) ;
    buf_clk cell_11071 ( .C (clk), .D (signal_13616), .Q (signal_13617) ) ;
    buf_clk cell_11087 ( .C (clk), .D (signal_13632), .Q (signal_13633) ) ;
    buf_clk cell_11103 ( .C (clk), .D (signal_13648), .Q (signal_13649) ) ;
    buf_clk cell_11119 ( .C (clk), .D (signal_13664), .Q (signal_13665) ) ;
    buf_clk cell_11135 ( .C (clk), .D (signal_13680), .Q (signal_13681) ) ;
    buf_clk cell_11151 ( .C (clk), .D (signal_13696), .Q (signal_13697) ) ;
    buf_clk cell_11167 ( .C (clk), .D (signal_13712), .Q (signal_13713) ) ;
    buf_clk cell_11183 ( .C (clk), .D (signal_13728), .Q (signal_13729) ) ;
    buf_clk cell_11199 ( .C (clk), .D (signal_13744), .Q (signal_13745) ) ;
    buf_clk cell_11215 ( .C (clk), .D (signal_13760), .Q (signal_13761) ) ;
    buf_clk cell_11231 ( .C (clk), .D (signal_13776), .Q (signal_13777) ) ;
    buf_clk cell_11247 ( .C (clk), .D (signal_13792), .Q (signal_13793) ) ;
    buf_clk cell_11263 ( .C (clk), .D (signal_13808), .Q (signal_13809) ) ;
    buf_clk cell_11279 ( .C (clk), .D (signal_13824), .Q (signal_13825) ) ;
    buf_clk cell_11295 ( .C (clk), .D (signal_13840), .Q (signal_13841) ) ;
    buf_clk cell_11311 ( .C (clk), .D (signal_13856), .Q (signal_13857) ) ;
    buf_clk cell_11327 ( .C (clk), .D (signal_13872), .Q (signal_13873) ) ;
    buf_clk cell_11343 ( .C (clk), .D (signal_13888), .Q (signal_13889) ) ;
    buf_clk cell_11359 ( .C (clk), .D (signal_13904), .Q (signal_13905) ) ;
    buf_clk cell_11375 ( .C (clk), .D (signal_13920), .Q (signal_13921) ) ;
    buf_clk cell_11391 ( .C (clk), .D (signal_13936), .Q (signal_13937) ) ;
    buf_clk cell_11407 ( .C (clk), .D (signal_13952), .Q (signal_13953) ) ;
    buf_clk cell_11423 ( .C (clk), .D (signal_13968), .Q (signal_13969) ) ;
    buf_clk cell_11439 ( .C (clk), .D (signal_13984), .Q (signal_13985) ) ;
    buf_clk cell_11455 ( .C (clk), .D (signal_14000), .Q (signal_14001) ) ;
    buf_clk cell_11471 ( .C (clk), .D (signal_14016), .Q (signal_14017) ) ;
    buf_clk cell_11487 ( .C (clk), .D (signal_14032), .Q (signal_14033) ) ;
    buf_clk cell_11503 ( .C (clk), .D (signal_14048), .Q (signal_14049) ) ;
    buf_clk cell_11519 ( .C (clk), .D (signal_14064), .Q (signal_14065) ) ;
    buf_clk cell_11535 ( .C (clk), .D (signal_14080), .Q (signal_14081) ) ;
    buf_clk cell_11551 ( .C (clk), .D (signal_14096), .Q (signal_14097) ) ;
    buf_clk cell_11567 ( .C (clk), .D (signal_14112), .Q (signal_14113) ) ;
    buf_clk cell_11583 ( .C (clk), .D (signal_14128), .Q (signal_14129) ) ;
    buf_clk cell_11599 ( .C (clk), .D (signal_14144), .Q (signal_14145) ) ;
    buf_clk cell_11615 ( .C (clk), .D (signal_14160), .Q (signal_14161) ) ;
    buf_clk cell_11631 ( .C (clk), .D (signal_14176), .Q (signal_14177) ) ;
    buf_clk cell_11647 ( .C (clk), .D (signal_14192), .Q (signal_14193) ) ;
    buf_clk cell_11663 ( .C (clk), .D (signal_14208), .Q (signal_14209) ) ;
    buf_clk cell_11679 ( .C (clk), .D (signal_14224), .Q (signal_14225) ) ;
    buf_clk cell_11695 ( .C (clk), .D (signal_14240), .Q (signal_14241) ) ;
    buf_clk cell_11711 ( .C (clk), .D (signal_14256), .Q (signal_14257) ) ;
    buf_clk cell_11727 ( .C (clk), .D (signal_14272), .Q (signal_14273) ) ;
    buf_clk cell_11743 ( .C (clk), .D (signal_14288), .Q (signal_14289) ) ;
    buf_clk cell_11759 ( .C (clk), .D (signal_14304), .Q (signal_14305) ) ;
    buf_clk cell_11775 ( .C (clk), .D (signal_14320), .Q (signal_14321) ) ;
    buf_clk cell_11791 ( .C (clk), .D (signal_14336), .Q (signal_14337) ) ;
    buf_clk cell_11807 ( .C (clk), .D (signal_14352), .Q (signal_14353) ) ;
    buf_clk cell_11823 ( .C (clk), .D (signal_14368), .Q (signal_14369) ) ;
    buf_clk cell_11839 ( .C (clk), .D (signal_14384), .Q (signal_14385) ) ;
    buf_clk cell_11855 ( .C (clk), .D (signal_14400), .Q (signal_14401) ) ;
    buf_clk cell_11871 ( .C (clk), .D (signal_14416), .Q (signal_14417) ) ;
    buf_clk cell_11887 ( .C (clk), .D (signal_14432), .Q (signal_14433) ) ;
    buf_clk cell_11903 ( .C (clk), .D (signal_14448), .Q (signal_14449) ) ;
    buf_clk cell_11919 ( .C (clk), .D (signal_14464), .Q (signal_14465) ) ;
    buf_clk cell_11935 ( .C (clk), .D (signal_14480), .Q (signal_14481) ) ;
    buf_clk cell_11951 ( .C (clk), .D (signal_14496), .Q (signal_14497) ) ;
    buf_clk cell_11967 ( .C (clk), .D (signal_14512), .Q (signal_14513) ) ;
    buf_clk cell_11983 ( .C (clk), .D (signal_14528), .Q (signal_14529) ) ;
    buf_clk cell_11999 ( .C (clk), .D (signal_14544), .Q (signal_14545) ) ;
    buf_clk cell_12015 ( .C (clk), .D (signal_14560), .Q (signal_14561) ) ;
    buf_clk cell_12031 ( .C (clk), .D (signal_14576), .Q (signal_14577) ) ;
    buf_clk cell_12047 ( .C (clk), .D (signal_14592), .Q (signal_14593) ) ;
    buf_clk cell_12063 ( .C (clk), .D (signal_14608), .Q (signal_14609) ) ;
    buf_clk cell_12079 ( .C (clk), .D (signal_14624), .Q (signal_14625) ) ;
    buf_clk cell_12095 ( .C (clk), .D (signal_14640), .Q (signal_14641) ) ;
    buf_clk cell_12111 ( .C (clk), .D (signal_14656), .Q (signal_14657) ) ;
    buf_clk cell_12127 ( .C (clk), .D (signal_14672), .Q (signal_14673) ) ;
    buf_clk cell_12143 ( .C (clk), .D (signal_14688), .Q (signal_14689) ) ;
    buf_clk cell_12159 ( .C (clk), .D (signal_14704), .Q (signal_14705) ) ;
    buf_clk cell_12175 ( .C (clk), .D (signal_14720), .Q (signal_14721) ) ;
    buf_clk cell_12191 ( .C (clk), .D (signal_14736), .Q (signal_14737) ) ;
    buf_clk cell_12207 ( .C (clk), .D (signal_14752), .Q (signal_14753) ) ;
    buf_clk cell_12223 ( .C (clk), .D (signal_14768), .Q (signal_14769) ) ;
    buf_clk cell_12239 ( .C (clk), .D (signal_14784), .Q (signal_14785) ) ;
    buf_clk cell_12255 ( .C (clk), .D (signal_14800), .Q (signal_14801) ) ;
    buf_clk cell_12271 ( .C (clk), .D (signal_14816), .Q (signal_14817) ) ;
    buf_clk cell_12287 ( .C (clk), .D (signal_14832), .Q (signal_14833) ) ;
    buf_clk cell_12303 ( .C (clk), .D (signal_14848), .Q (signal_14849) ) ;
    buf_clk cell_12319 ( .C (clk), .D (signal_14864), .Q (signal_14865) ) ;
    buf_clk cell_12335 ( .C (clk), .D (signal_14880), .Q (signal_14881) ) ;
    buf_clk cell_12351 ( .C (clk), .D (signal_14896), .Q (signal_14897) ) ;
    buf_clk cell_12367 ( .C (clk), .D (signal_14912), .Q (signal_14913) ) ;
    buf_clk cell_12383 ( .C (clk), .D (signal_14928), .Q (signal_14929) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1719 ( .s ({signal_4694, signal_4692}), .b ({signal_3273, signal_1982}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[5]), .c ({signal_3418, signal_1987}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1720 ( .s ({signal_4694, signal_4692}), .b ({signal_3274, signal_1983}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[6]), .c ({signal_3419, signal_1988}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1721 ( .s ({signal_4694, signal_4692}), .b ({1'b0, 1'b1}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[7]), .c ({signal_3420, signal_1989}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1722 ( .s ({signal_4694, signal_4692}), .b ({signal_3274, signal_1983}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[8]), .c ({signal_3421, signal_1990}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1723 ( .s ({signal_4694, signal_4692}), .b ({1'b0, 1'b0}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[9]), .c ({signal_3422, signal_1991}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1724 ( .s ({signal_4694, signal_4692}), .b ({signal_3273, signal_1982}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[10]), .c ({signal_3423, signal_1992}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1725 ( .s ({signal_4698, signal_4696}), .b ({signal_3273, signal_1982}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[11]), .c ({signal_3424, signal_1993}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1726 ( .s ({signal_4694, signal_4692}), .b ({1'b0, 1'b0}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[12]), .c ({signal_3425, signal_1994}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1727 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b1}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[13]), .c ({signal_3426, signal_1995}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1728 ( .s ({signal_4694, signal_4692}), .b ({signal_3273, signal_1982}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[14]), .c ({signal_3427, signal_1996}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1729 ( .s ({signal_4694, signal_4692}), .b ({1'b0, 1'b1}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[15]), .c ({signal_3428, signal_1997}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1730 ( .s ({signal_4698, signal_4696}), .b ({signal_3274, signal_1983}), .a ({signal_3276, signal_1985}), .clk (clk), .r (Fresh[16]), .c ({signal_3429, signal_1998}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1731 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b1}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[17]), .c ({signal_3430, signal_1999}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1732 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b0}), .a ({signal_3275, signal_1984}), .clk (clk), .r (Fresh[18]), .c ({signal_3431, signal_2000}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1733 ( .s ({signal_4698, signal_4696}), .b ({signal_3276, signal_1985}), .a ({signal_3275, signal_1984}), .clk (clk), .r (Fresh[19]), .c ({signal_3432, signal_2001}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1734 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b0}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[20]), .c ({signal_3433, signal_2002}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1735 ( .s ({signal_4694, signal_4692}), .b ({signal_3274, signal_1983}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[21]), .c ({signal_3434, signal_2003}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1736 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b0}), .a ({signal_3276, signal_1985}), .clk (clk), .r (Fresh[22]), .c ({signal_3435, signal_2004}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1737 ( .s ({signal_4698, signal_4696}), .b ({signal_3274, signal_1983}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[23]), .c ({signal_3436, signal_2005}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1738 ( .s ({signal_4698, signal_4696}), .b ({signal_3273, signal_1982}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[24]), .c ({signal_3437, signal_2006}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1739 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b1}), .a ({signal_3275, signal_1984}), .clk (clk), .r (Fresh[25]), .c ({signal_3438, signal_2007}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1740 ( .s ({signal_4698, signal_4696}), .b ({signal_3275, signal_1984}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[26]), .c ({signal_3439, signal_2008}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1741 ( .s ({signal_4698, signal_4696}), .b ({signal_3275, signal_1984}), .a ({signal_3276, signal_1985}), .clk (clk), .r (Fresh[27]), .c ({signal_3440, signal_2009}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1742 ( .s ({signal_4698, signal_4696}), .b ({signal_3275, signal_1984}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[28]), .c ({signal_3441, signal_2010}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1743 ( .s ({signal_4698, signal_4696}), .b ({signal_3276, signal_1985}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[29]), .c ({signal_3442, signal_2011}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1744 ( .s ({signal_4698, signal_4696}), .b ({signal_3274, signal_1983}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[30]), .c ({signal_3443, signal_2012}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1745 ( .s ({signal_4698, signal_4696}), .b ({1'b0, 1'b1}), .a ({signal_3276, signal_1985}), .clk (clk), .r (Fresh[31]), .c ({signal_3444, signal_2013}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1746 ( .s ({signal_4698, signal_4696}), .b ({signal_3275, signal_1984}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[32]), .c ({signal_3445, signal_2014}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1747 ( .s ({signal_4698, signal_4696}), .b ({signal_3273, signal_1982}), .a ({signal_3276, signal_1985}), .clk (clk), .r (Fresh[33]), .c ({signal_3446, signal_2015}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1748 ( .s ({signal_4698, signal_4696}), .b ({signal_3276, signal_1985}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[34]), .c ({signal_3447, signal_2016}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1749 ( .s ({signal_4698, signal_4696}), .b ({signal_3276, signal_1985}), .a ({signal_3273, signal_1982}), .clk (clk), .r (Fresh[35]), .c ({signal_3448, signal_2017}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1750 ( .s ({signal_4698, signal_4696}), .b ({signal_3275, signal_1984}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[36]), .c ({signal_3449, signal_2018}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1751 ( .s ({signal_4698, signal_4696}), .b ({signal_3273, signal_1982}), .a ({signal_3274, signal_1983}), .clk (clk), .r (Fresh[37]), .c ({signal_3450, signal_2019}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1752 ( .s ({signal_4698, signal_4696}), .b ({signal_3274, signal_1983}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[38]), .c ({signal_3451, signal_2020}) ) ;
    buf_clk cell_2154 ( .C (clk), .D (signal_4699), .Q (signal_4700) ) ;
    buf_clk cell_2156 ( .C (clk), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_2158 ( .C (clk), .D (signal_4703), .Q (signal_4704) ) ;
    buf_clk cell_2160 ( .C (clk), .D (signal_4705), .Q (signal_4706) ) ;
    buf_clk cell_2162 ( .C (clk), .D (signal_4707), .Q (signal_4708) ) ;
    buf_clk cell_2164 ( .C (clk), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_2166 ( .C (clk), .D (signal_4711), .Q (signal_4712) ) ;
    buf_clk cell_2168 ( .C (clk), .D (signal_4713), .Q (signal_4714) ) ;
    buf_clk cell_2172 ( .C (clk), .D (signal_4717), .Q (signal_4718) ) ;
    buf_clk cell_2176 ( .C (clk), .D (signal_4721), .Q (signal_4722) ) ;
    buf_clk cell_2178 ( .C (clk), .D (signal_4723), .Q (signal_4724) ) ;
    buf_clk cell_2180 ( .C (clk), .D (signal_4725), .Q (signal_4726) ) ;
    buf_clk cell_2182 ( .C (clk), .D (signal_4727), .Q (signal_4728) ) ;
    buf_clk cell_2184 ( .C (clk), .D (signal_4729), .Q (signal_4730) ) ;
    buf_clk cell_2300 ( .C (clk), .D (signal_4845), .Q (signal_4846) ) ;
    buf_clk cell_2308 ( .C (clk), .D (signal_4853), .Q (signal_4854) ) ;
    buf_clk cell_2344 ( .C (clk), .D (signal_4889), .Q (signal_4890) ) ;
    buf_clk cell_2354 ( .C (clk), .D (signal_4899), .Q (signal_4900) ) ;
    buf_clk cell_2364 ( .C (clk), .D (signal_4909), .Q (signal_4910) ) ;
    buf_clk cell_2376 ( .C (clk), .D (signal_4921), .Q (signal_4922) ) ;
    buf_clk cell_2388 ( .C (clk), .D (signal_4933), .Q (signal_4934) ) ;
    buf_clk cell_2404 ( .C (clk), .D (signal_4949), .Q (signal_4950) ) ;
    buf_clk cell_2420 ( .C (clk), .D (signal_4965), .Q (signal_4966) ) ;
    buf_clk cell_2436 ( .C (clk), .D (signal_4981), .Q (signal_4982) ) ;
    buf_clk cell_2452 ( .C (clk), .D (signal_4997), .Q (signal_4998) ) ;
    buf_clk cell_2468 ( .C (clk), .D (signal_5013), .Q (signal_5014) ) ;
    buf_clk cell_2484 ( .C (clk), .D (signal_5029), .Q (signal_5030) ) ;
    buf_clk cell_2500 ( .C (clk), .D (signal_5045), .Q (signal_5046) ) ;
    buf_clk cell_2516 ( .C (clk), .D (signal_5061), .Q (signal_5062) ) ;
    buf_clk cell_2532 ( .C (clk), .D (signal_5077), .Q (signal_5078) ) ;
    buf_clk cell_2548 ( .C (clk), .D (signal_5093), .Q (signal_5094) ) ;
    buf_clk cell_2564 ( .C (clk), .D (signal_5109), .Q (signal_5110) ) ;
    buf_clk cell_2580 ( .C (clk), .D (signal_5125), .Q (signal_5126) ) ;
    buf_clk cell_2596 ( .C (clk), .D (signal_5141), .Q (signal_5142) ) ;
    buf_clk cell_2612 ( .C (clk), .D (signal_5157), .Q (signal_5158) ) ;
    buf_clk cell_2628 ( .C (clk), .D (signal_5173), .Q (signal_5174) ) ;
    buf_clk cell_2644 ( .C (clk), .D (signal_5189), .Q (signal_5190) ) ;
    buf_clk cell_2660 ( .C (clk), .D (signal_5205), .Q (signal_5206) ) ;
    buf_clk cell_2676 ( .C (clk), .D (signal_5221), .Q (signal_5222) ) ;
    buf_clk cell_2692 ( .C (clk), .D (signal_5237), .Q (signal_5238) ) ;
    buf_clk cell_2708 ( .C (clk), .D (signal_5253), .Q (signal_5254) ) ;
    buf_clk cell_2724 ( .C (clk), .D (signal_5269), .Q (signal_5270) ) ;
    buf_clk cell_2740 ( .C (clk), .D (signal_5285), .Q (signal_5286) ) ;
    buf_clk cell_2756 ( .C (clk), .D (signal_5301), .Q (signal_5302) ) ;
    buf_clk cell_2772 ( .C (clk), .D (signal_5317), .Q (signal_5318) ) ;
    buf_clk cell_2788 ( .C (clk), .D (signal_5333), .Q (signal_5334) ) ;
    buf_clk cell_2804 ( .C (clk), .D (signal_5349), .Q (signal_5350) ) ;
    buf_clk cell_2820 ( .C (clk), .D (signal_5365), .Q (signal_5366) ) ;
    buf_clk cell_2836 ( .C (clk), .D (signal_5381), .Q (signal_5382) ) ;
    buf_clk cell_2852 ( .C (clk), .D (signal_5397), .Q (signal_5398) ) ;
    buf_clk cell_2868 ( .C (clk), .D (signal_5413), .Q (signal_5414) ) ;
    buf_clk cell_2884 ( .C (clk), .D (signal_5429), .Q (signal_5430) ) ;
    buf_clk cell_2900 ( .C (clk), .D (signal_5445), .Q (signal_5446) ) ;
    buf_clk cell_2916 ( .C (clk), .D (signal_5461), .Q (signal_5462) ) ;
    buf_clk cell_2932 ( .C (clk), .D (signal_5477), .Q (signal_5478) ) ;
    buf_clk cell_2948 ( .C (clk), .D (signal_5493), .Q (signal_5494) ) ;
    buf_clk cell_2964 ( .C (clk), .D (signal_5509), .Q (signal_5510) ) ;
    buf_clk cell_2980 ( .C (clk), .D (signal_5525), .Q (signal_5526) ) ;
    buf_clk cell_2996 ( .C (clk), .D (signal_5541), .Q (signal_5542) ) ;
    buf_clk cell_3012 ( .C (clk), .D (signal_5557), .Q (signal_5558) ) ;
    buf_clk cell_3028 ( .C (clk), .D (signal_5573), .Q (signal_5574) ) ;
    buf_clk cell_3044 ( .C (clk), .D (signal_5589), .Q (signal_5590) ) ;
    buf_clk cell_3060 ( .C (clk), .D (signal_5605), .Q (signal_5606) ) ;
    buf_clk cell_3076 ( .C (clk), .D (signal_5621), .Q (signal_5622) ) ;
    buf_clk cell_3092 ( .C (clk), .D (signal_5637), .Q (signal_5638) ) ;
    buf_clk cell_3108 ( .C (clk), .D (signal_5653), .Q (signal_5654) ) ;
    buf_clk cell_3124 ( .C (clk), .D (signal_5669), .Q (signal_5670) ) ;
    buf_clk cell_3140 ( .C (clk), .D (signal_5685), .Q (signal_5686) ) ;
    buf_clk cell_3156 ( .C (clk), .D (signal_5701), .Q (signal_5702) ) ;
    buf_clk cell_3172 ( .C (clk), .D (signal_5717), .Q (signal_5718) ) ;
    buf_clk cell_3188 ( .C (clk), .D (signal_5733), .Q (signal_5734) ) ;
    buf_clk cell_3204 ( .C (clk), .D (signal_5749), .Q (signal_5750) ) ;
    buf_clk cell_3220 ( .C (clk), .D (signal_5765), .Q (signal_5766) ) ;
    buf_clk cell_3236 ( .C (clk), .D (signal_5781), .Q (signal_5782) ) ;
    buf_clk cell_3252 ( .C (clk), .D (signal_5797), .Q (signal_5798) ) ;
    buf_clk cell_3268 ( .C (clk), .D (signal_5813), .Q (signal_5814) ) ;
    buf_clk cell_3284 ( .C (clk), .D (signal_5829), .Q (signal_5830) ) ;
    buf_clk cell_3300 ( .C (clk), .D (signal_5845), .Q (signal_5846) ) ;
    buf_clk cell_3316 ( .C (clk), .D (signal_5861), .Q (signal_5862) ) ;
    buf_clk cell_3332 ( .C (clk), .D (signal_5877), .Q (signal_5878) ) ;
    buf_clk cell_3348 ( .C (clk), .D (signal_5893), .Q (signal_5894) ) ;
    buf_clk cell_3364 ( .C (clk), .D (signal_5909), .Q (signal_5910) ) ;
    buf_clk cell_3380 ( .C (clk), .D (signal_5925), .Q (signal_5926) ) ;
    buf_clk cell_3396 ( .C (clk), .D (signal_5941), .Q (signal_5942) ) ;
    buf_clk cell_3412 ( .C (clk), .D (signal_5957), .Q (signal_5958) ) ;
    buf_clk cell_3428 ( .C (clk), .D (signal_5973), .Q (signal_5974) ) ;
    buf_clk cell_3444 ( .C (clk), .D (signal_5989), .Q (signal_5990) ) ;
    buf_clk cell_3460 ( .C (clk), .D (signal_6005), .Q (signal_6006) ) ;
    buf_clk cell_3476 ( .C (clk), .D (signal_6021), .Q (signal_6022) ) ;
    buf_clk cell_3492 ( .C (clk), .D (signal_6037), .Q (signal_6038) ) ;
    buf_clk cell_3508 ( .C (clk), .D (signal_6053), .Q (signal_6054) ) ;
    buf_clk cell_3524 ( .C (clk), .D (signal_6069), .Q (signal_6070) ) ;
    buf_clk cell_3540 ( .C (clk), .D (signal_6085), .Q (signal_6086) ) ;
    buf_clk cell_3556 ( .C (clk), .D (signal_6101), .Q (signal_6102) ) ;
    buf_clk cell_3572 ( .C (clk), .D (signal_6117), .Q (signal_6118) ) ;
    buf_clk cell_3588 ( .C (clk), .D (signal_6133), .Q (signal_6134) ) ;
    buf_clk cell_3604 ( .C (clk), .D (signal_6149), .Q (signal_6150) ) ;
    buf_clk cell_3620 ( .C (clk), .D (signal_6165), .Q (signal_6166) ) ;
    buf_clk cell_3636 ( .C (clk), .D (signal_6181), .Q (signal_6182) ) ;
    buf_clk cell_3652 ( .C (clk), .D (signal_6197), .Q (signal_6198) ) ;
    buf_clk cell_3668 ( .C (clk), .D (signal_6213), .Q (signal_6214) ) ;
    buf_clk cell_3684 ( .C (clk), .D (signal_6229), .Q (signal_6230) ) ;
    buf_clk cell_3700 ( .C (clk), .D (signal_6245), .Q (signal_6246) ) ;
    buf_clk cell_3716 ( .C (clk), .D (signal_6261), .Q (signal_6262) ) ;
    buf_clk cell_3732 ( .C (clk), .D (signal_6277), .Q (signal_6278) ) ;
    buf_clk cell_3748 ( .C (clk), .D (signal_6293), .Q (signal_6294) ) ;
    buf_clk cell_3764 ( .C (clk), .D (signal_6309), .Q (signal_6310) ) ;
    buf_clk cell_3780 ( .C (clk), .D (signal_6325), .Q (signal_6326) ) ;
    buf_clk cell_3796 ( .C (clk), .D (signal_6341), .Q (signal_6342) ) ;
    buf_clk cell_3812 ( .C (clk), .D (signal_6357), .Q (signal_6358) ) ;
    buf_clk cell_3828 ( .C (clk), .D (signal_6373), .Q (signal_6374) ) ;
    buf_clk cell_3844 ( .C (clk), .D (signal_6389), .Q (signal_6390) ) ;
    buf_clk cell_3860 ( .C (clk), .D (signal_6405), .Q (signal_6406) ) ;
    buf_clk cell_3876 ( .C (clk), .D (signal_6421), .Q (signal_6422) ) ;
    buf_clk cell_3892 ( .C (clk), .D (signal_6437), .Q (signal_6438) ) ;
    buf_clk cell_3908 ( .C (clk), .D (signal_6453), .Q (signal_6454) ) ;
    buf_clk cell_3924 ( .C (clk), .D (signal_6469), .Q (signal_6470) ) ;
    buf_clk cell_3940 ( .C (clk), .D (signal_6485), .Q (signal_6486) ) ;
    buf_clk cell_3956 ( .C (clk), .D (signal_6501), .Q (signal_6502) ) ;
    buf_clk cell_3972 ( .C (clk), .D (signal_6517), .Q (signal_6518) ) ;
    buf_clk cell_3988 ( .C (clk), .D (signal_6533), .Q (signal_6534) ) ;
    buf_clk cell_4004 ( .C (clk), .D (signal_6549), .Q (signal_6550) ) ;
    buf_clk cell_4020 ( .C (clk), .D (signal_6565), .Q (signal_6566) ) ;
    buf_clk cell_4036 ( .C (clk), .D (signal_6581), .Q (signal_6582) ) ;
    buf_clk cell_4052 ( .C (clk), .D (signal_6597), .Q (signal_6598) ) ;
    buf_clk cell_4068 ( .C (clk), .D (signal_6613), .Q (signal_6614) ) ;
    buf_clk cell_4084 ( .C (clk), .D (signal_6629), .Q (signal_6630) ) ;
    buf_clk cell_4100 ( .C (clk), .D (signal_6645), .Q (signal_6646) ) ;
    buf_clk cell_4116 ( .C (clk), .D (signal_6661), .Q (signal_6662) ) ;
    buf_clk cell_4132 ( .C (clk), .D (signal_6677), .Q (signal_6678) ) ;
    buf_clk cell_4148 ( .C (clk), .D (signal_6693), .Q (signal_6694) ) ;
    buf_clk cell_4164 ( .C (clk), .D (signal_6709), .Q (signal_6710) ) ;
    buf_clk cell_4180 ( .C (clk), .D (signal_6725), .Q (signal_6726) ) ;
    buf_clk cell_4196 ( .C (clk), .D (signal_6741), .Q (signal_6742) ) ;
    buf_clk cell_4212 ( .C (clk), .D (signal_6757), .Q (signal_6758) ) ;
    buf_clk cell_4228 ( .C (clk), .D (signal_6773), .Q (signal_6774) ) ;
    buf_clk cell_4244 ( .C (clk), .D (signal_6789), .Q (signal_6790) ) ;
    buf_clk cell_4260 ( .C (clk), .D (signal_6805), .Q (signal_6806) ) ;
    buf_clk cell_4276 ( .C (clk), .D (signal_6821), .Q (signal_6822) ) ;
    buf_clk cell_4292 ( .C (clk), .D (signal_6837), .Q (signal_6838) ) ;
    buf_clk cell_4308 ( .C (clk), .D (signal_6853), .Q (signal_6854) ) ;
    buf_clk cell_4324 ( .C (clk), .D (signal_6869), .Q (signal_6870) ) ;
    buf_clk cell_4340 ( .C (clk), .D (signal_6885), .Q (signal_6886) ) ;
    buf_clk cell_4356 ( .C (clk), .D (signal_6901), .Q (signal_6902) ) ;
    buf_clk cell_4372 ( .C (clk), .D (signal_6917), .Q (signal_6918) ) ;
    buf_clk cell_4388 ( .C (clk), .D (signal_6933), .Q (signal_6934) ) ;
    buf_clk cell_4404 ( .C (clk), .D (signal_6949), .Q (signal_6950) ) ;
    buf_clk cell_4418 ( .C (clk), .D (signal_6963), .Q (signal_6964) ) ;
    buf_clk cell_4432 ( .C (clk), .D (signal_6977), .Q (signal_6978) ) ;
    buf_clk cell_4448 ( .C (clk), .D (signal_6993), .Q (signal_6994) ) ;
    buf_clk cell_4464 ( .C (clk), .D (signal_7009), .Q (signal_7010) ) ;
    buf_clk cell_4480 ( .C (clk), .D (signal_7025), .Q (signal_7026) ) ;
    buf_clk cell_4496 ( .C (clk), .D (signal_7041), .Q (signal_7042) ) ;
    buf_clk cell_4512 ( .C (clk), .D (signal_7057), .Q (signal_7058) ) ;
    buf_clk cell_4528 ( .C (clk), .D (signal_7073), .Q (signal_7074) ) ;
    buf_clk cell_4544 ( .C (clk), .D (signal_7089), .Q (signal_7090) ) ;
    buf_clk cell_4560 ( .C (clk), .D (signal_7105), .Q (signal_7106) ) ;
    buf_clk cell_4576 ( .C (clk), .D (signal_7121), .Q (signal_7122) ) ;
    buf_clk cell_4592 ( .C (clk), .D (signal_7137), .Q (signal_7138) ) ;
    buf_clk cell_4608 ( .C (clk), .D (signal_7153), .Q (signal_7154) ) ;
    buf_clk cell_4624 ( .C (clk), .D (signal_7169), .Q (signal_7170) ) ;
    buf_clk cell_4640 ( .C (clk), .D (signal_7185), .Q (signal_7186) ) ;
    buf_clk cell_4656 ( .C (clk), .D (signal_7201), .Q (signal_7202) ) ;
    buf_clk cell_4672 ( .C (clk), .D (signal_7217), .Q (signal_7218) ) ;
    buf_clk cell_4688 ( .C (clk), .D (signal_7233), .Q (signal_7234) ) ;
    buf_clk cell_4704 ( .C (clk), .D (signal_7249), .Q (signal_7250) ) ;
    buf_clk cell_4720 ( .C (clk), .D (signal_7265), .Q (signal_7266) ) ;
    buf_clk cell_4736 ( .C (clk), .D (signal_7281), .Q (signal_7282) ) ;
    buf_clk cell_4752 ( .C (clk), .D (signal_7297), .Q (signal_7298) ) ;
    buf_clk cell_4768 ( .C (clk), .D (signal_7313), .Q (signal_7314) ) ;
    buf_clk cell_4784 ( .C (clk), .D (signal_7329), .Q (signal_7330) ) ;
    buf_clk cell_4800 ( .C (clk), .D (signal_7345), .Q (signal_7346) ) ;
    buf_clk cell_4816 ( .C (clk), .D (signal_7361), .Q (signal_7362) ) ;
    buf_clk cell_4832 ( .C (clk), .D (signal_7377), .Q (signal_7378) ) ;
    buf_clk cell_4848 ( .C (clk), .D (signal_7393), .Q (signal_7394) ) ;
    buf_clk cell_4864 ( .C (clk), .D (signal_7409), .Q (signal_7410) ) ;
    buf_clk cell_4880 ( .C (clk), .D (signal_7425), .Q (signal_7426) ) ;
    buf_clk cell_4896 ( .C (clk), .D (signal_7441), .Q (signal_7442) ) ;
    buf_clk cell_4912 ( .C (clk), .D (signal_7457), .Q (signal_7458) ) ;
    buf_clk cell_4928 ( .C (clk), .D (signal_7473), .Q (signal_7474) ) ;
    buf_clk cell_4944 ( .C (clk), .D (signal_7489), .Q (signal_7490) ) ;
    buf_clk cell_4960 ( .C (clk), .D (signal_7505), .Q (signal_7506) ) ;
    buf_clk cell_4976 ( .C (clk), .D (signal_7521), .Q (signal_7522) ) ;
    buf_clk cell_4992 ( .C (clk), .D (signal_7537), .Q (signal_7538) ) ;
    buf_clk cell_5008 ( .C (clk), .D (signal_7553), .Q (signal_7554) ) ;
    buf_clk cell_5024 ( .C (clk), .D (signal_7569), .Q (signal_7570) ) ;
    buf_clk cell_5040 ( .C (clk), .D (signal_7585), .Q (signal_7586) ) ;
    buf_clk cell_5056 ( .C (clk), .D (signal_7601), .Q (signal_7602) ) ;
    buf_clk cell_5072 ( .C (clk), .D (signal_7617), .Q (signal_7618) ) ;
    buf_clk cell_5088 ( .C (clk), .D (signal_7633), .Q (signal_7634) ) ;
    buf_clk cell_5104 ( .C (clk), .D (signal_7649), .Q (signal_7650) ) ;
    buf_clk cell_5120 ( .C (clk), .D (signal_7665), .Q (signal_7666) ) ;
    buf_clk cell_5136 ( .C (clk), .D (signal_7681), .Q (signal_7682) ) ;
    buf_clk cell_5152 ( .C (clk), .D (signal_7697), .Q (signal_7698) ) ;
    buf_clk cell_5168 ( .C (clk), .D (signal_7713), .Q (signal_7714) ) ;
    buf_clk cell_5184 ( .C (clk), .D (signal_7729), .Q (signal_7730) ) ;
    buf_clk cell_5200 ( .C (clk), .D (signal_7745), .Q (signal_7746) ) ;
    buf_clk cell_5216 ( .C (clk), .D (signal_7761), .Q (signal_7762) ) ;
    buf_clk cell_5232 ( .C (clk), .D (signal_7777), .Q (signal_7778) ) ;
    buf_clk cell_5248 ( .C (clk), .D (signal_7793), .Q (signal_7794) ) ;
    buf_clk cell_5264 ( .C (clk), .D (signal_7809), .Q (signal_7810) ) ;
    buf_clk cell_5280 ( .C (clk), .D (signal_7825), .Q (signal_7826) ) ;
    buf_clk cell_5296 ( .C (clk), .D (signal_7841), .Q (signal_7842) ) ;
    buf_clk cell_5312 ( .C (clk), .D (signal_7857), .Q (signal_7858) ) ;
    buf_clk cell_5328 ( .C (clk), .D (signal_7873), .Q (signal_7874) ) ;
    buf_clk cell_5344 ( .C (clk), .D (signal_7889), .Q (signal_7890) ) ;
    buf_clk cell_5360 ( .C (clk), .D (signal_7905), .Q (signal_7906) ) ;
    buf_clk cell_5376 ( .C (clk), .D (signal_7921), .Q (signal_7922) ) ;
    buf_clk cell_5392 ( .C (clk), .D (signal_7937), .Q (signal_7938) ) ;
    buf_clk cell_5408 ( .C (clk), .D (signal_7953), .Q (signal_7954) ) ;
    buf_clk cell_5424 ( .C (clk), .D (signal_7969), .Q (signal_7970) ) ;
    buf_clk cell_5440 ( .C (clk), .D (signal_7985), .Q (signal_7986) ) ;
    buf_clk cell_5456 ( .C (clk), .D (signal_8001), .Q (signal_8002) ) ;
    buf_clk cell_5472 ( .C (clk), .D (signal_8017), .Q (signal_8018) ) ;
    buf_clk cell_5488 ( .C (clk), .D (signal_8033), .Q (signal_8034) ) ;
    buf_clk cell_5504 ( .C (clk), .D (signal_8049), .Q (signal_8050) ) ;
    buf_clk cell_5520 ( .C (clk), .D (signal_8065), .Q (signal_8066) ) ;
    buf_clk cell_5536 ( .C (clk), .D (signal_8081), .Q (signal_8082) ) ;
    buf_clk cell_5552 ( .C (clk), .D (signal_8097), .Q (signal_8098) ) ;
    buf_clk cell_5568 ( .C (clk), .D (signal_8113), .Q (signal_8114) ) ;
    buf_clk cell_5584 ( .C (clk), .D (signal_8129), .Q (signal_8130) ) ;
    buf_clk cell_5600 ( .C (clk), .D (signal_8145), .Q (signal_8146) ) ;
    buf_clk cell_5616 ( .C (clk), .D (signal_8161), .Q (signal_8162) ) ;
    buf_clk cell_5632 ( .C (clk), .D (signal_8177), .Q (signal_8178) ) ;
    buf_clk cell_5648 ( .C (clk), .D (signal_8193), .Q (signal_8194) ) ;
    buf_clk cell_5664 ( .C (clk), .D (signal_8209), .Q (signal_8210) ) ;
    buf_clk cell_5680 ( .C (clk), .D (signal_8225), .Q (signal_8226) ) ;
    buf_clk cell_5696 ( .C (clk), .D (signal_8241), .Q (signal_8242) ) ;
    buf_clk cell_5712 ( .C (clk), .D (signal_8257), .Q (signal_8258) ) ;
    buf_clk cell_5728 ( .C (clk), .D (signal_8273), .Q (signal_8274) ) ;
    buf_clk cell_5744 ( .C (clk), .D (signal_8289), .Q (signal_8290) ) ;
    buf_clk cell_5760 ( .C (clk), .D (signal_8305), .Q (signal_8306) ) ;
    buf_clk cell_5776 ( .C (clk), .D (signal_8321), .Q (signal_8322) ) ;
    buf_clk cell_5792 ( .C (clk), .D (signal_8337), .Q (signal_8338) ) ;
    buf_clk cell_5808 ( .C (clk), .D (signal_8353), .Q (signal_8354) ) ;
    buf_clk cell_5824 ( .C (clk), .D (signal_8369), .Q (signal_8370) ) ;
    buf_clk cell_5840 ( .C (clk), .D (signal_8385), .Q (signal_8386) ) ;
    buf_clk cell_5856 ( .C (clk), .D (signal_8401), .Q (signal_8402) ) ;
    buf_clk cell_5872 ( .C (clk), .D (signal_8417), .Q (signal_8418) ) ;
    buf_clk cell_5888 ( .C (clk), .D (signal_8433), .Q (signal_8434) ) ;
    buf_clk cell_5904 ( .C (clk), .D (signal_8449), .Q (signal_8450) ) ;
    buf_clk cell_5920 ( .C (clk), .D (signal_8465), .Q (signal_8466) ) ;
    buf_clk cell_5936 ( .C (clk), .D (signal_8481), .Q (signal_8482) ) ;
    buf_clk cell_5952 ( .C (clk), .D (signal_8497), .Q (signal_8498) ) ;
    buf_clk cell_5968 ( .C (clk), .D (signal_8513), .Q (signal_8514) ) ;
    buf_clk cell_5984 ( .C (clk), .D (signal_8529), .Q (signal_8530) ) ;
    buf_clk cell_6000 ( .C (clk), .D (signal_8545), .Q (signal_8546) ) ;
    buf_clk cell_6016 ( .C (clk), .D (signal_8561), .Q (signal_8562) ) ;
    buf_clk cell_6032 ( .C (clk), .D (signal_8577), .Q (signal_8578) ) ;
    buf_clk cell_6048 ( .C (clk), .D (signal_8593), .Q (signal_8594) ) ;
    buf_clk cell_6064 ( .C (clk), .D (signal_8609), .Q (signal_8610) ) ;
    buf_clk cell_6080 ( .C (clk), .D (signal_8625), .Q (signal_8626) ) ;
    buf_clk cell_6096 ( .C (clk), .D (signal_8641), .Q (signal_8642) ) ;
    buf_clk cell_6112 ( .C (clk), .D (signal_8657), .Q (signal_8658) ) ;
    buf_clk cell_6128 ( .C (clk), .D (signal_8673), .Q (signal_8674) ) ;
    buf_clk cell_6144 ( .C (clk), .D (signal_8689), .Q (signal_8690) ) ;
    buf_clk cell_6160 ( .C (clk), .D (signal_8705), .Q (signal_8706) ) ;
    buf_clk cell_6176 ( .C (clk), .D (signal_8721), .Q (signal_8722) ) ;
    buf_clk cell_6192 ( .C (clk), .D (signal_8737), .Q (signal_8738) ) ;
    buf_clk cell_6208 ( .C (clk), .D (signal_8753), .Q (signal_8754) ) ;
    buf_clk cell_6224 ( .C (clk), .D (signal_8769), .Q (signal_8770) ) ;
    buf_clk cell_6240 ( .C (clk), .D (signal_8785), .Q (signal_8786) ) ;
    buf_clk cell_6256 ( .C (clk), .D (signal_8801), .Q (signal_8802) ) ;
    buf_clk cell_6272 ( .C (clk), .D (signal_8817), .Q (signal_8818) ) ;
    buf_clk cell_6288 ( .C (clk), .D (signal_8833), .Q (signal_8834) ) ;
    buf_clk cell_6304 ( .C (clk), .D (signal_8849), .Q (signal_8850) ) ;
    buf_clk cell_6320 ( .C (clk), .D (signal_8865), .Q (signal_8866) ) ;
    buf_clk cell_6336 ( .C (clk), .D (signal_8881), .Q (signal_8882) ) ;
    buf_clk cell_6352 ( .C (clk), .D (signal_8897), .Q (signal_8898) ) ;
    buf_clk cell_6368 ( .C (clk), .D (signal_8913), .Q (signal_8914) ) ;
    buf_clk cell_6384 ( .C (clk), .D (signal_8929), .Q (signal_8930) ) ;
    buf_clk cell_6400 ( .C (clk), .D (signal_8945), .Q (signal_8946) ) ;
    buf_clk cell_6416 ( .C (clk), .D (signal_8961), .Q (signal_8962) ) ;
    buf_clk cell_6432 ( .C (clk), .D (signal_8977), .Q (signal_8978) ) ;
    buf_clk cell_6448 ( .C (clk), .D (signal_8993), .Q (signal_8994) ) ;
    buf_clk cell_6464 ( .C (clk), .D (signal_9009), .Q (signal_9010) ) ;
    buf_clk cell_6480 ( .C (clk), .D (signal_9025), .Q (signal_9026) ) ;
    buf_clk cell_6496 ( .C (clk), .D (signal_9041), .Q (signal_9042) ) ;
    buf_clk cell_6512 ( .C (clk), .D (signal_9057), .Q (signal_9058) ) ;
    buf_clk cell_6528 ( .C (clk), .D (signal_9073), .Q (signal_9074) ) ;
    buf_clk cell_6544 ( .C (clk), .D (signal_9089), .Q (signal_9090) ) ;
    buf_clk cell_6560 ( .C (clk), .D (signal_9105), .Q (signal_9106) ) ;
    buf_clk cell_6576 ( .C (clk), .D (signal_9121), .Q (signal_9122) ) ;
    buf_clk cell_6592 ( .C (clk), .D (signal_9137), .Q (signal_9138) ) ;
    buf_clk cell_6608 ( .C (clk), .D (signal_9153), .Q (signal_9154) ) ;
    buf_clk cell_6624 ( .C (clk), .D (signal_9169), .Q (signal_9170) ) ;
    buf_clk cell_6640 ( .C (clk), .D (signal_9185), .Q (signal_9186) ) ;
    buf_clk cell_6656 ( .C (clk), .D (signal_9201), .Q (signal_9202) ) ;
    buf_clk cell_6672 ( .C (clk), .D (signal_9217), .Q (signal_9218) ) ;
    buf_clk cell_6688 ( .C (clk), .D (signal_9233), .Q (signal_9234) ) ;
    buf_clk cell_6704 ( .C (clk), .D (signal_9249), .Q (signal_9250) ) ;
    buf_clk cell_6720 ( .C (clk), .D (signal_9265), .Q (signal_9266) ) ;
    buf_clk cell_6736 ( .C (clk), .D (signal_9281), .Q (signal_9282) ) ;
    buf_clk cell_6752 ( .C (clk), .D (signal_9297), .Q (signal_9298) ) ;
    buf_clk cell_6768 ( .C (clk), .D (signal_9313), .Q (signal_9314) ) ;
    buf_clk cell_6784 ( .C (clk), .D (signal_9329), .Q (signal_9330) ) ;
    buf_clk cell_6800 ( .C (clk), .D (signal_9345), .Q (signal_9346) ) ;
    buf_clk cell_6816 ( .C (clk), .D (signal_9361), .Q (signal_9362) ) ;
    buf_clk cell_6832 ( .C (clk), .D (signal_9377), .Q (signal_9378) ) ;
    buf_clk cell_6848 ( .C (clk), .D (signal_9393), .Q (signal_9394) ) ;
    buf_clk cell_6864 ( .C (clk), .D (signal_9409), .Q (signal_9410) ) ;
    buf_clk cell_6880 ( .C (clk), .D (signal_9425), .Q (signal_9426) ) ;
    buf_clk cell_6896 ( .C (clk), .D (signal_9441), .Q (signal_9442) ) ;
    buf_clk cell_6912 ( .C (clk), .D (signal_9457), .Q (signal_9458) ) ;
    buf_clk cell_6928 ( .C (clk), .D (signal_9473), .Q (signal_9474) ) ;
    buf_clk cell_6944 ( .C (clk), .D (signal_9489), .Q (signal_9490) ) ;
    buf_clk cell_6960 ( .C (clk), .D (signal_9505), .Q (signal_9506) ) ;
    buf_clk cell_6976 ( .C (clk), .D (signal_9521), .Q (signal_9522) ) ;
    buf_clk cell_6992 ( .C (clk), .D (signal_9537), .Q (signal_9538) ) ;
    buf_clk cell_7008 ( .C (clk), .D (signal_9553), .Q (signal_9554) ) ;
    buf_clk cell_7024 ( .C (clk), .D (signal_9569), .Q (signal_9570) ) ;
    buf_clk cell_7040 ( .C (clk), .D (signal_9585), .Q (signal_9586) ) ;
    buf_clk cell_7056 ( .C (clk), .D (signal_9601), .Q (signal_9602) ) ;
    buf_clk cell_7072 ( .C (clk), .D (signal_9617), .Q (signal_9618) ) ;
    buf_clk cell_7088 ( .C (clk), .D (signal_9633), .Q (signal_9634) ) ;
    buf_clk cell_7104 ( .C (clk), .D (signal_9649), .Q (signal_9650) ) ;
    buf_clk cell_7120 ( .C (clk), .D (signal_9665), .Q (signal_9666) ) ;
    buf_clk cell_7136 ( .C (clk), .D (signal_9681), .Q (signal_9682) ) ;
    buf_clk cell_7152 ( .C (clk), .D (signal_9697), .Q (signal_9698) ) ;
    buf_clk cell_7168 ( .C (clk), .D (signal_9713), .Q (signal_9714) ) ;
    buf_clk cell_7184 ( .C (clk), .D (signal_9729), .Q (signal_9730) ) ;
    buf_clk cell_7200 ( .C (clk), .D (signal_9745), .Q (signal_9746) ) ;
    buf_clk cell_7216 ( .C (clk), .D (signal_9761), .Q (signal_9762) ) ;
    buf_clk cell_7232 ( .C (clk), .D (signal_9777), .Q (signal_9778) ) ;
    buf_clk cell_7248 ( .C (clk), .D (signal_9793), .Q (signal_9794) ) ;
    buf_clk cell_7264 ( .C (clk), .D (signal_9809), .Q (signal_9810) ) ;
    buf_clk cell_7280 ( .C (clk), .D (signal_9825), .Q (signal_9826) ) ;
    buf_clk cell_7296 ( .C (clk), .D (signal_9841), .Q (signal_9842) ) ;
    buf_clk cell_7312 ( .C (clk), .D (signal_9857), .Q (signal_9858) ) ;
    buf_clk cell_7328 ( .C (clk), .D (signal_9873), .Q (signal_9874) ) ;
    buf_clk cell_7344 ( .C (clk), .D (signal_9889), .Q (signal_9890) ) ;
    buf_clk cell_7360 ( .C (clk), .D (signal_9905), .Q (signal_9906) ) ;
    buf_clk cell_7376 ( .C (clk), .D (signal_9921), .Q (signal_9922) ) ;
    buf_clk cell_7392 ( .C (clk), .D (signal_9937), .Q (signal_9938) ) ;
    buf_clk cell_7408 ( .C (clk), .D (signal_9953), .Q (signal_9954) ) ;
    buf_clk cell_7424 ( .C (clk), .D (signal_9969), .Q (signal_9970) ) ;
    buf_clk cell_7440 ( .C (clk), .D (signal_9985), .Q (signal_9986) ) ;
    buf_clk cell_7456 ( .C (clk), .D (signal_10001), .Q (signal_10002) ) ;
    buf_clk cell_7472 ( .C (clk), .D (signal_10017), .Q (signal_10018) ) ;
    buf_clk cell_7488 ( .C (clk), .D (signal_10033), .Q (signal_10034) ) ;
    buf_clk cell_7504 ( .C (clk), .D (signal_10049), .Q (signal_10050) ) ;
    buf_clk cell_7520 ( .C (clk), .D (signal_10065), .Q (signal_10066) ) ;
    buf_clk cell_7536 ( .C (clk), .D (signal_10081), .Q (signal_10082) ) ;
    buf_clk cell_7552 ( .C (clk), .D (signal_10097), .Q (signal_10098) ) ;
    buf_clk cell_7568 ( .C (clk), .D (signal_10113), .Q (signal_10114) ) ;
    buf_clk cell_7584 ( .C (clk), .D (signal_10129), .Q (signal_10130) ) ;
    buf_clk cell_7600 ( .C (clk), .D (signal_10145), .Q (signal_10146) ) ;
    buf_clk cell_7616 ( .C (clk), .D (signal_10161), .Q (signal_10162) ) ;
    buf_clk cell_7632 ( .C (clk), .D (signal_10177), .Q (signal_10178) ) ;
    buf_clk cell_7648 ( .C (clk), .D (signal_10193), .Q (signal_10194) ) ;
    buf_clk cell_7664 ( .C (clk), .D (signal_10209), .Q (signal_10210) ) ;
    buf_clk cell_7680 ( .C (clk), .D (signal_10225), .Q (signal_10226) ) ;
    buf_clk cell_7696 ( .C (clk), .D (signal_10241), .Q (signal_10242) ) ;
    buf_clk cell_7712 ( .C (clk), .D (signal_10257), .Q (signal_10258) ) ;
    buf_clk cell_7728 ( .C (clk), .D (signal_10273), .Q (signal_10274) ) ;
    buf_clk cell_7744 ( .C (clk), .D (signal_10289), .Q (signal_10290) ) ;
    buf_clk cell_7760 ( .C (clk), .D (signal_10305), .Q (signal_10306) ) ;
    buf_clk cell_7776 ( .C (clk), .D (signal_10321), .Q (signal_10322) ) ;
    buf_clk cell_7792 ( .C (clk), .D (signal_10337), .Q (signal_10338) ) ;
    buf_clk cell_7808 ( .C (clk), .D (signal_10353), .Q (signal_10354) ) ;
    buf_clk cell_7824 ( .C (clk), .D (signal_10369), .Q (signal_10370) ) ;
    buf_clk cell_7840 ( .C (clk), .D (signal_10385), .Q (signal_10386) ) ;
    buf_clk cell_7856 ( .C (clk), .D (signal_10401), .Q (signal_10402) ) ;
    buf_clk cell_7872 ( .C (clk), .D (signal_10417), .Q (signal_10418) ) ;
    buf_clk cell_7888 ( .C (clk), .D (signal_10433), .Q (signal_10434) ) ;
    buf_clk cell_7904 ( .C (clk), .D (signal_10449), .Q (signal_10450) ) ;
    buf_clk cell_7920 ( .C (clk), .D (signal_10465), .Q (signal_10466) ) ;
    buf_clk cell_7936 ( .C (clk), .D (signal_10481), .Q (signal_10482) ) ;
    buf_clk cell_7952 ( .C (clk), .D (signal_10497), .Q (signal_10498) ) ;
    buf_clk cell_7968 ( .C (clk), .D (signal_10513), .Q (signal_10514) ) ;
    buf_clk cell_7984 ( .C (clk), .D (signal_10529), .Q (signal_10530) ) ;
    buf_clk cell_8000 ( .C (clk), .D (signal_10545), .Q (signal_10546) ) ;
    buf_clk cell_8016 ( .C (clk), .D (signal_10561), .Q (signal_10562) ) ;
    buf_clk cell_8032 ( .C (clk), .D (signal_10577), .Q (signal_10578) ) ;
    buf_clk cell_8048 ( .C (clk), .D (signal_10593), .Q (signal_10594) ) ;
    buf_clk cell_8064 ( .C (clk), .D (signal_10609), .Q (signal_10610) ) ;
    buf_clk cell_8080 ( .C (clk), .D (signal_10625), .Q (signal_10626) ) ;
    buf_clk cell_8096 ( .C (clk), .D (signal_10641), .Q (signal_10642) ) ;
    buf_clk cell_8112 ( .C (clk), .D (signal_10657), .Q (signal_10658) ) ;
    buf_clk cell_8128 ( .C (clk), .D (signal_10673), .Q (signal_10674) ) ;
    buf_clk cell_8144 ( .C (clk), .D (signal_10689), .Q (signal_10690) ) ;
    buf_clk cell_8160 ( .C (clk), .D (signal_10705), .Q (signal_10706) ) ;
    buf_clk cell_8176 ( .C (clk), .D (signal_10721), .Q (signal_10722) ) ;
    buf_clk cell_8192 ( .C (clk), .D (signal_10737), .Q (signal_10738) ) ;
    buf_clk cell_8208 ( .C (clk), .D (signal_10753), .Q (signal_10754) ) ;
    buf_clk cell_8224 ( .C (clk), .D (signal_10769), .Q (signal_10770) ) ;
    buf_clk cell_8240 ( .C (clk), .D (signal_10785), .Q (signal_10786) ) ;
    buf_clk cell_8256 ( .C (clk), .D (signal_10801), .Q (signal_10802) ) ;
    buf_clk cell_8272 ( .C (clk), .D (signal_10817), .Q (signal_10818) ) ;
    buf_clk cell_8288 ( .C (clk), .D (signal_10833), .Q (signal_10834) ) ;
    buf_clk cell_8304 ( .C (clk), .D (signal_10849), .Q (signal_10850) ) ;
    buf_clk cell_8320 ( .C (clk), .D (signal_10865), .Q (signal_10866) ) ;
    buf_clk cell_8336 ( .C (clk), .D (signal_10881), .Q (signal_10882) ) ;
    buf_clk cell_8352 ( .C (clk), .D (signal_10897), .Q (signal_10898) ) ;
    buf_clk cell_8368 ( .C (clk), .D (signal_10913), .Q (signal_10914) ) ;
    buf_clk cell_8384 ( .C (clk), .D (signal_10929), .Q (signal_10930) ) ;
    buf_clk cell_8400 ( .C (clk), .D (signal_10945), .Q (signal_10946) ) ;
    buf_clk cell_8416 ( .C (clk), .D (signal_10961), .Q (signal_10962) ) ;
    buf_clk cell_8432 ( .C (clk), .D (signal_10977), .Q (signal_10978) ) ;
    buf_clk cell_8448 ( .C (clk), .D (signal_10993), .Q (signal_10994) ) ;
    buf_clk cell_8464 ( .C (clk), .D (signal_11009), .Q (signal_11010) ) ;
    buf_clk cell_8480 ( .C (clk), .D (signal_11025), .Q (signal_11026) ) ;
    buf_clk cell_8496 ( .C (clk), .D (signal_11041), .Q (signal_11042) ) ;
    buf_clk cell_8512 ( .C (clk), .D (signal_11057), .Q (signal_11058) ) ;
    buf_clk cell_8528 ( .C (clk), .D (signal_11073), .Q (signal_11074) ) ;
    buf_clk cell_8544 ( .C (clk), .D (signal_11089), .Q (signal_11090) ) ;
    buf_clk cell_8560 ( .C (clk), .D (signal_11105), .Q (signal_11106) ) ;
    buf_clk cell_8576 ( .C (clk), .D (signal_11121), .Q (signal_11122) ) ;
    buf_clk cell_8592 ( .C (clk), .D (signal_11137), .Q (signal_11138) ) ;
    buf_clk cell_8608 ( .C (clk), .D (signal_11153), .Q (signal_11154) ) ;
    buf_clk cell_8624 ( .C (clk), .D (signal_11169), .Q (signal_11170) ) ;
    buf_clk cell_8640 ( .C (clk), .D (signal_11185), .Q (signal_11186) ) ;
    buf_clk cell_8656 ( .C (clk), .D (signal_11201), .Q (signal_11202) ) ;
    buf_clk cell_8672 ( .C (clk), .D (signal_11217), .Q (signal_11218) ) ;
    buf_clk cell_8688 ( .C (clk), .D (signal_11233), .Q (signal_11234) ) ;
    buf_clk cell_8704 ( .C (clk), .D (signal_11249), .Q (signal_11250) ) ;
    buf_clk cell_8720 ( .C (clk), .D (signal_11265), .Q (signal_11266) ) ;
    buf_clk cell_8736 ( .C (clk), .D (signal_11281), .Q (signal_11282) ) ;
    buf_clk cell_8752 ( .C (clk), .D (signal_11297), .Q (signal_11298) ) ;
    buf_clk cell_8768 ( .C (clk), .D (signal_11313), .Q (signal_11314) ) ;
    buf_clk cell_8784 ( .C (clk), .D (signal_11329), .Q (signal_11330) ) ;
    buf_clk cell_8800 ( .C (clk), .D (signal_11345), .Q (signal_11346) ) ;
    buf_clk cell_8816 ( .C (clk), .D (signal_11361), .Q (signal_11362) ) ;
    buf_clk cell_8832 ( .C (clk), .D (signal_11377), .Q (signal_11378) ) ;
    buf_clk cell_8848 ( .C (clk), .D (signal_11393), .Q (signal_11394) ) ;
    buf_clk cell_8864 ( .C (clk), .D (signal_11409), .Q (signal_11410) ) ;
    buf_clk cell_8880 ( .C (clk), .D (signal_11425), .Q (signal_11426) ) ;
    buf_clk cell_8896 ( .C (clk), .D (signal_11441), .Q (signal_11442) ) ;
    buf_clk cell_8912 ( .C (clk), .D (signal_11457), .Q (signal_11458) ) ;
    buf_clk cell_8928 ( .C (clk), .D (signal_11473), .Q (signal_11474) ) ;
    buf_clk cell_8944 ( .C (clk), .D (signal_11489), .Q (signal_11490) ) ;
    buf_clk cell_8960 ( .C (clk), .D (signal_11505), .Q (signal_11506) ) ;
    buf_clk cell_8976 ( .C (clk), .D (signal_11521), .Q (signal_11522) ) ;
    buf_clk cell_8992 ( .C (clk), .D (signal_11537), .Q (signal_11538) ) ;
    buf_clk cell_9008 ( .C (clk), .D (signal_11553), .Q (signal_11554) ) ;
    buf_clk cell_9024 ( .C (clk), .D (signal_11569), .Q (signal_11570) ) ;
    buf_clk cell_9040 ( .C (clk), .D (signal_11585), .Q (signal_11586) ) ;
    buf_clk cell_9056 ( .C (clk), .D (signal_11601), .Q (signal_11602) ) ;
    buf_clk cell_9072 ( .C (clk), .D (signal_11617), .Q (signal_11618) ) ;
    buf_clk cell_9088 ( .C (clk), .D (signal_11633), .Q (signal_11634) ) ;
    buf_clk cell_9104 ( .C (clk), .D (signal_11649), .Q (signal_11650) ) ;
    buf_clk cell_9120 ( .C (clk), .D (signal_11665), .Q (signal_11666) ) ;
    buf_clk cell_9136 ( .C (clk), .D (signal_11681), .Q (signal_11682) ) ;
    buf_clk cell_9152 ( .C (clk), .D (signal_11697), .Q (signal_11698) ) ;
    buf_clk cell_9168 ( .C (clk), .D (signal_11713), .Q (signal_11714) ) ;
    buf_clk cell_9184 ( .C (clk), .D (signal_11729), .Q (signal_11730) ) ;
    buf_clk cell_9200 ( .C (clk), .D (signal_11745), .Q (signal_11746) ) ;
    buf_clk cell_9216 ( .C (clk), .D (signal_11761), .Q (signal_11762) ) ;
    buf_clk cell_9232 ( .C (clk), .D (signal_11777), .Q (signal_11778) ) ;
    buf_clk cell_9248 ( .C (clk), .D (signal_11793), .Q (signal_11794) ) ;
    buf_clk cell_9264 ( .C (clk), .D (signal_11809), .Q (signal_11810) ) ;
    buf_clk cell_9280 ( .C (clk), .D (signal_11825), .Q (signal_11826) ) ;
    buf_clk cell_9296 ( .C (clk), .D (signal_11841), .Q (signal_11842) ) ;
    buf_clk cell_9312 ( .C (clk), .D (signal_11857), .Q (signal_11858) ) ;
    buf_clk cell_9328 ( .C (clk), .D (signal_11873), .Q (signal_11874) ) ;
    buf_clk cell_9344 ( .C (clk), .D (signal_11889), .Q (signal_11890) ) ;
    buf_clk cell_9360 ( .C (clk), .D (signal_11905), .Q (signal_11906) ) ;
    buf_clk cell_9376 ( .C (clk), .D (signal_11921), .Q (signal_11922) ) ;
    buf_clk cell_9392 ( .C (clk), .D (signal_11937), .Q (signal_11938) ) ;
    buf_clk cell_9408 ( .C (clk), .D (signal_11953), .Q (signal_11954) ) ;
    buf_clk cell_9424 ( .C (clk), .D (signal_11969), .Q (signal_11970) ) ;
    buf_clk cell_9440 ( .C (clk), .D (signal_11985), .Q (signal_11986) ) ;
    buf_clk cell_9456 ( .C (clk), .D (signal_12001), .Q (signal_12002) ) ;
    buf_clk cell_9472 ( .C (clk), .D (signal_12017), .Q (signal_12018) ) ;
    buf_clk cell_9488 ( .C (clk), .D (signal_12033), .Q (signal_12034) ) ;
    buf_clk cell_9504 ( .C (clk), .D (signal_12049), .Q (signal_12050) ) ;
    buf_clk cell_9520 ( .C (clk), .D (signal_12065), .Q (signal_12066) ) ;
    buf_clk cell_9536 ( .C (clk), .D (signal_12081), .Q (signal_12082) ) ;
    buf_clk cell_9552 ( .C (clk), .D (signal_12097), .Q (signal_12098) ) ;
    buf_clk cell_9568 ( .C (clk), .D (signal_12113), .Q (signal_12114) ) ;
    buf_clk cell_9584 ( .C (clk), .D (signal_12129), .Q (signal_12130) ) ;
    buf_clk cell_9600 ( .C (clk), .D (signal_12145), .Q (signal_12146) ) ;
    buf_clk cell_9616 ( .C (clk), .D (signal_12161), .Q (signal_12162) ) ;
    buf_clk cell_9632 ( .C (clk), .D (signal_12177), .Q (signal_12178) ) ;
    buf_clk cell_9648 ( .C (clk), .D (signal_12193), .Q (signal_12194) ) ;
    buf_clk cell_9664 ( .C (clk), .D (signal_12209), .Q (signal_12210) ) ;
    buf_clk cell_9680 ( .C (clk), .D (signal_12225), .Q (signal_12226) ) ;
    buf_clk cell_9696 ( .C (clk), .D (signal_12241), .Q (signal_12242) ) ;
    buf_clk cell_9712 ( .C (clk), .D (signal_12257), .Q (signal_12258) ) ;
    buf_clk cell_9728 ( .C (clk), .D (signal_12273), .Q (signal_12274) ) ;
    buf_clk cell_9744 ( .C (clk), .D (signal_12289), .Q (signal_12290) ) ;
    buf_clk cell_9760 ( .C (clk), .D (signal_12305), .Q (signal_12306) ) ;
    buf_clk cell_9776 ( .C (clk), .D (signal_12321), .Q (signal_12322) ) ;
    buf_clk cell_9792 ( .C (clk), .D (signal_12337), .Q (signal_12338) ) ;
    buf_clk cell_9808 ( .C (clk), .D (signal_12353), .Q (signal_12354) ) ;
    buf_clk cell_9824 ( .C (clk), .D (signal_12369), .Q (signal_12370) ) ;
    buf_clk cell_9840 ( .C (clk), .D (signal_12385), .Q (signal_12386) ) ;
    buf_clk cell_9856 ( .C (clk), .D (signal_12401), .Q (signal_12402) ) ;
    buf_clk cell_9872 ( .C (clk), .D (signal_12417), .Q (signal_12418) ) ;
    buf_clk cell_9888 ( .C (clk), .D (signal_12433), .Q (signal_12434) ) ;
    buf_clk cell_9904 ( .C (clk), .D (signal_12449), .Q (signal_12450) ) ;
    buf_clk cell_9920 ( .C (clk), .D (signal_12465), .Q (signal_12466) ) ;
    buf_clk cell_9936 ( .C (clk), .D (signal_12481), .Q (signal_12482) ) ;
    buf_clk cell_9952 ( .C (clk), .D (signal_12497), .Q (signal_12498) ) ;
    buf_clk cell_9968 ( .C (clk), .D (signal_12513), .Q (signal_12514) ) ;
    buf_clk cell_9984 ( .C (clk), .D (signal_12529), .Q (signal_12530) ) ;
    buf_clk cell_10000 ( .C (clk), .D (signal_12545), .Q (signal_12546) ) ;
    buf_clk cell_10016 ( .C (clk), .D (signal_12561), .Q (signal_12562) ) ;
    buf_clk cell_10032 ( .C (clk), .D (signal_12577), .Q (signal_12578) ) ;
    buf_clk cell_10048 ( .C (clk), .D (signal_12593), .Q (signal_12594) ) ;
    buf_clk cell_10064 ( .C (clk), .D (signal_12609), .Q (signal_12610) ) ;
    buf_clk cell_10080 ( .C (clk), .D (signal_12625), .Q (signal_12626) ) ;
    buf_clk cell_10096 ( .C (clk), .D (signal_12641), .Q (signal_12642) ) ;
    buf_clk cell_10112 ( .C (clk), .D (signal_12657), .Q (signal_12658) ) ;
    buf_clk cell_10128 ( .C (clk), .D (signal_12673), .Q (signal_12674) ) ;
    buf_clk cell_10144 ( .C (clk), .D (signal_12689), .Q (signal_12690) ) ;
    buf_clk cell_10160 ( .C (clk), .D (signal_12705), .Q (signal_12706) ) ;
    buf_clk cell_10176 ( .C (clk), .D (signal_12721), .Q (signal_12722) ) ;
    buf_clk cell_10192 ( .C (clk), .D (signal_12737), .Q (signal_12738) ) ;
    buf_clk cell_10208 ( .C (clk), .D (signal_12753), .Q (signal_12754) ) ;
    buf_clk cell_10224 ( .C (clk), .D (signal_12769), .Q (signal_12770) ) ;
    buf_clk cell_10240 ( .C (clk), .D (signal_12785), .Q (signal_12786) ) ;
    buf_clk cell_10256 ( .C (clk), .D (signal_12801), .Q (signal_12802) ) ;
    buf_clk cell_10272 ( .C (clk), .D (signal_12817), .Q (signal_12818) ) ;
    buf_clk cell_10288 ( .C (clk), .D (signal_12833), .Q (signal_12834) ) ;
    buf_clk cell_10304 ( .C (clk), .D (signal_12849), .Q (signal_12850) ) ;
    buf_clk cell_10320 ( .C (clk), .D (signal_12865), .Q (signal_12866) ) ;
    buf_clk cell_10336 ( .C (clk), .D (signal_12881), .Q (signal_12882) ) ;
    buf_clk cell_10352 ( .C (clk), .D (signal_12897), .Q (signal_12898) ) ;
    buf_clk cell_10368 ( .C (clk), .D (signal_12913), .Q (signal_12914) ) ;
    buf_clk cell_10384 ( .C (clk), .D (signal_12929), .Q (signal_12930) ) ;
    buf_clk cell_10400 ( .C (clk), .D (signal_12945), .Q (signal_12946) ) ;
    buf_clk cell_10416 ( .C (clk), .D (signal_12961), .Q (signal_12962) ) ;
    buf_clk cell_10432 ( .C (clk), .D (signal_12977), .Q (signal_12978) ) ;
    buf_clk cell_10448 ( .C (clk), .D (signal_12993), .Q (signal_12994) ) ;
    buf_clk cell_10464 ( .C (clk), .D (signal_13009), .Q (signal_13010) ) ;
    buf_clk cell_10480 ( .C (clk), .D (signal_13025), .Q (signal_13026) ) ;
    buf_clk cell_10496 ( .C (clk), .D (signal_13041), .Q (signal_13042) ) ;
    buf_clk cell_10512 ( .C (clk), .D (signal_13057), .Q (signal_13058) ) ;
    buf_clk cell_10528 ( .C (clk), .D (signal_13073), .Q (signal_13074) ) ;
    buf_clk cell_10544 ( .C (clk), .D (signal_13089), .Q (signal_13090) ) ;
    buf_clk cell_10560 ( .C (clk), .D (signal_13105), .Q (signal_13106) ) ;
    buf_clk cell_10576 ( .C (clk), .D (signal_13121), .Q (signal_13122) ) ;
    buf_clk cell_10592 ( .C (clk), .D (signal_13137), .Q (signal_13138) ) ;
    buf_clk cell_10608 ( .C (clk), .D (signal_13153), .Q (signal_13154) ) ;
    buf_clk cell_10624 ( .C (clk), .D (signal_13169), .Q (signal_13170) ) ;
    buf_clk cell_10640 ( .C (clk), .D (signal_13185), .Q (signal_13186) ) ;
    buf_clk cell_10656 ( .C (clk), .D (signal_13201), .Q (signal_13202) ) ;
    buf_clk cell_10672 ( .C (clk), .D (signal_13217), .Q (signal_13218) ) ;
    buf_clk cell_10688 ( .C (clk), .D (signal_13233), .Q (signal_13234) ) ;
    buf_clk cell_10704 ( .C (clk), .D (signal_13249), .Q (signal_13250) ) ;
    buf_clk cell_10720 ( .C (clk), .D (signal_13265), .Q (signal_13266) ) ;
    buf_clk cell_10736 ( .C (clk), .D (signal_13281), .Q (signal_13282) ) ;
    buf_clk cell_10752 ( .C (clk), .D (signal_13297), .Q (signal_13298) ) ;
    buf_clk cell_10768 ( .C (clk), .D (signal_13313), .Q (signal_13314) ) ;
    buf_clk cell_10784 ( .C (clk), .D (signal_13329), .Q (signal_13330) ) ;
    buf_clk cell_10800 ( .C (clk), .D (signal_13345), .Q (signal_13346) ) ;
    buf_clk cell_10816 ( .C (clk), .D (signal_13361), .Q (signal_13362) ) ;
    buf_clk cell_10832 ( .C (clk), .D (signal_13377), .Q (signal_13378) ) ;
    buf_clk cell_10848 ( .C (clk), .D (signal_13393), .Q (signal_13394) ) ;
    buf_clk cell_10864 ( .C (clk), .D (signal_13409), .Q (signal_13410) ) ;
    buf_clk cell_10880 ( .C (clk), .D (signal_13425), .Q (signal_13426) ) ;
    buf_clk cell_10896 ( .C (clk), .D (signal_13441), .Q (signal_13442) ) ;
    buf_clk cell_10912 ( .C (clk), .D (signal_13457), .Q (signal_13458) ) ;
    buf_clk cell_10928 ( .C (clk), .D (signal_13473), .Q (signal_13474) ) ;
    buf_clk cell_10944 ( .C (clk), .D (signal_13489), .Q (signal_13490) ) ;
    buf_clk cell_10960 ( .C (clk), .D (signal_13505), .Q (signal_13506) ) ;
    buf_clk cell_10976 ( .C (clk), .D (signal_13521), .Q (signal_13522) ) ;
    buf_clk cell_10992 ( .C (clk), .D (signal_13537), .Q (signal_13538) ) ;
    buf_clk cell_11008 ( .C (clk), .D (signal_13553), .Q (signal_13554) ) ;
    buf_clk cell_11024 ( .C (clk), .D (signal_13569), .Q (signal_13570) ) ;
    buf_clk cell_11040 ( .C (clk), .D (signal_13585), .Q (signal_13586) ) ;
    buf_clk cell_11056 ( .C (clk), .D (signal_13601), .Q (signal_13602) ) ;
    buf_clk cell_11072 ( .C (clk), .D (signal_13617), .Q (signal_13618) ) ;
    buf_clk cell_11088 ( .C (clk), .D (signal_13633), .Q (signal_13634) ) ;
    buf_clk cell_11104 ( .C (clk), .D (signal_13649), .Q (signal_13650) ) ;
    buf_clk cell_11120 ( .C (clk), .D (signal_13665), .Q (signal_13666) ) ;
    buf_clk cell_11136 ( .C (clk), .D (signal_13681), .Q (signal_13682) ) ;
    buf_clk cell_11152 ( .C (clk), .D (signal_13697), .Q (signal_13698) ) ;
    buf_clk cell_11168 ( .C (clk), .D (signal_13713), .Q (signal_13714) ) ;
    buf_clk cell_11184 ( .C (clk), .D (signal_13729), .Q (signal_13730) ) ;
    buf_clk cell_11200 ( .C (clk), .D (signal_13745), .Q (signal_13746) ) ;
    buf_clk cell_11216 ( .C (clk), .D (signal_13761), .Q (signal_13762) ) ;
    buf_clk cell_11232 ( .C (clk), .D (signal_13777), .Q (signal_13778) ) ;
    buf_clk cell_11248 ( .C (clk), .D (signal_13793), .Q (signal_13794) ) ;
    buf_clk cell_11264 ( .C (clk), .D (signal_13809), .Q (signal_13810) ) ;
    buf_clk cell_11280 ( .C (clk), .D (signal_13825), .Q (signal_13826) ) ;
    buf_clk cell_11296 ( .C (clk), .D (signal_13841), .Q (signal_13842) ) ;
    buf_clk cell_11312 ( .C (clk), .D (signal_13857), .Q (signal_13858) ) ;
    buf_clk cell_11328 ( .C (clk), .D (signal_13873), .Q (signal_13874) ) ;
    buf_clk cell_11344 ( .C (clk), .D (signal_13889), .Q (signal_13890) ) ;
    buf_clk cell_11360 ( .C (clk), .D (signal_13905), .Q (signal_13906) ) ;
    buf_clk cell_11376 ( .C (clk), .D (signal_13921), .Q (signal_13922) ) ;
    buf_clk cell_11392 ( .C (clk), .D (signal_13937), .Q (signal_13938) ) ;
    buf_clk cell_11408 ( .C (clk), .D (signal_13953), .Q (signal_13954) ) ;
    buf_clk cell_11424 ( .C (clk), .D (signal_13969), .Q (signal_13970) ) ;
    buf_clk cell_11440 ( .C (clk), .D (signal_13985), .Q (signal_13986) ) ;
    buf_clk cell_11456 ( .C (clk), .D (signal_14001), .Q (signal_14002) ) ;
    buf_clk cell_11472 ( .C (clk), .D (signal_14017), .Q (signal_14018) ) ;
    buf_clk cell_11488 ( .C (clk), .D (signal_14033), .Q (signal_14034) ) ;
    buf_clk cell_11504 ( .C (clk), .D (signal_14049), .Q (signal_14050) ) ;
    buf_clk cell_11520 ( .C (clk), .D (signal_14065), .Q (signal_14066) ) ;
    buf_clk cell_11536 ( .C (clk), .D (signal_14081), .Q (signal_14082) ) ;
    buf_clk cell_11552 ( .C (clk), .D (signal_14097), .Q (signal_14098) ) ;
    buf_clk cell_11568 ( .C (clk), .D (signal_14113), .Q (signal_14114) ) ;
    buf_clk cell_11584 ( .C (clk), .D (signal_14129), .Q (signal_14130) ) ;
    buf_clk cell_11600 ( .C (clk), .D (signal_14145), .Q (signal_14146) ) ;
    buf_clk cell_11616 ( .C (clk), .D (signal_14161), .Q (signal_14162) ) ;
    buf_clk cell_11632 ( .C (clk), .D (signal_14177), .Q (signal_14178) ) ;
    buf_clk cell_11648 ( .C (clk), .D (signal_14193), .Q (signal_14194) ) ;
    buf_clk cell_11664 ( .C (clk), .D (signal_14209), .Q (signal_14210) ) ;
    buf_clk cell_11680 ( .C (clk), .D (signal_14225), .Q (signal_14226) ) ;
    buf_clk cell_11696 ( .C (clk), .D (signal_14241), .Q (signal_14242) ) ;
    buf_clk cell_11712 ( .C (clk), .D (signal_14257), .Q (signal_14258) ) ;
    buf_clk cell_11728 ( .C (clk), .D (signal_14273), .Q (signal_14274) ) ;
    buf_clk cell_11744 ( .C (clk), .D (signal_14289), .Q (signal_14290) ) ;
    buf_clk cell_11760 ( .C (clk), .D (signal_14305), .Q (signal_14306) ) ;
    buf_clk cell_11776 ( .C (clk), .D (signal_14321), .Q (signal_14322) ) ;
    buf_clk cell_11792 ( .C (clk), .D (signal_14337), .Q (signal_14338) ) ;
    buf_clk cell_11808 ( .C (clk), .D (signal_14353), .Q (signal_14354) ) ;
    buf_clk cell_11824 ( .C (clk), .D (signal_14369), .Q (signal_14370) ) ;
    buf_clk cell_11840 ( .C (clk), .D (signal_14385), .Q (signal_14386) ) ;
    buf_clk cell_11856 ( .C (clk), .D (signal_14401), .Q (signal_14402) ) ;
    buf_clk cell_11872 ( .C (clk), .D (signal_14417), .Q (signal_14418) ) ;
    buf_clk cell_11888 ( .C (clk), .D (signal_14433), .Q (signal_14434) ) ;
    buf_clk cell_11904 ( .C (clk), .D (signal_14449), .Q (signal_14450) ) ;
    buf_clk cell_11920 ( .C (clk), .D (signal_14465), .Q (signal_14466) ) ;
    buf_clk cell_11936 ( .C (clk), .D (signal_14481), .Q (signal_14482) ) ;
    buf_clk cell_11952 ( .C (clk), .D (signal_14497), .Q (signal_14498) ) ;
    buf_clk cell_11968 ( .C (clk), .D (signal_14513), .Q (signal_14514) ) ;
    buf_clk cell_11984 ( .C (clk), .D (signal_14529), .Q (signal_14530) ) ;
    buf_clk cell_12000 ( .C (clk), .D (signal_14545), .Q (signal_14546) ) ;
    buf_clk cell_12016 ( .C (clk), .D (signal_14561), .Q (signal_14562) ) ;
    buf_clk cell_12032 ( .C (clk), .D (signal_14577), .Q (signal_14578) ) ;
    buf_clk cell_12048 ( .C (clk), .D (signal_14593), .Q (signal_14594) ) ;
    buf_clk cell_12064 ( .C (clk), .D (signal_14609), .Q (signal_14610) ) ;
    buf_clk cell_12080 ( .C (clk), .D (signal_14625), .Q (signal_14626) ) ;
    buf_clk cell_12096 ( .C (clk), .D (signal_14641), .Q (signal_14642) ) ;
    buf_clk cell_12112 ( .C (clk), .D (signal_14657), .Q (signal_14658) ) ;
    buf_clk cell_12128 ( .C (clk), .D (signal_14673), .Q (signal_14674) ) ;
    buf_clk cell_12144 ( .C (clk), .D (signal_14689), .Q (signal_14690) ) ;
    buf_clk cell_12160 ( .C (clk), .D (signal_14705), .Q (signal_14706) ) ;
    buf_clk cell_12176 ( .C (clk), .D (signal_14721), .Q (signal_14722) ) ;
    buf_clk cell_12192 ( .C (clk), .D (signal_14737), .Q (signal_14738) ) ;
    buf_clk cell_12208 ( .C (clk), .D (signal_14753), .Q (signal_14754) ) ;
    buf_clk cell_12224 ( .C (clk), .D (signal_14769), .Q (signal_14770) ) ;
    buf_clk cell_12240 ( .C (clk), .D (signal_14785), .Q (signal_14786) ) ;
    buf_clk cell_12256 ( .C (clk), .D (signal_14801), .Q (signal_14802) ) ;
    buf_clk cell_12272 ( .C (clk), .D (signal_14817), .Q (signal_14818) ) ;
    buf_clk cell_12288 ( .C (clk), .D (signal_14833), .Q (signal_14834) ) ;
    buf_clk cell_12304 ( .C (clk), .D (signal_14849), .Q (signal_14850) ) ;
    buf_clk cell_12320 ( .C (clk), .D (signal_14865), .Q (signal_14866) ) ;
    buf_clk cell_12336 ( .C (clk), .D (signal_14881), .Q (signal_14882) ) ;
    buf_clk cell_12352 ( .C (clk), .D (signal_14897), .Q (signal_14898) ) ;
    buf_clk cell_12368 ( .C (clk), .D (signal_14913), .Q (signal_14914) ) ;
    buf_clk cell_12384 ( .C (clk), .D (signal_14929), .Q (signal_14930) ) ;

    /* cells in depth 5 */
    buf_clk cell_2185 ( .C (clk), .D (signal_4718), .Q (signal_4731) ) ;
    buf_clk cell_2187 ( .C (clk), .D (signal_4722), .Q (signal_4733) ) ;
    buf_clk cell_2189 ( .C (clk), .D (signal_1993), .Q (signal_4735) ) ;
    buf_clk cell_2191 ( .C (clk), .D (signal_3424), .Q (signal_4737) ) ;
    buf_clk cell_2193 ( .C (clk), .D (signal_1995), .Q (signal_4739) ) ;
    buf_clk cell_2195 ( .C (clk), .D (signal_3426), .Q (signal_4741) ) ;
    buf_clk cell_2197 ( .C (clk), .D (signal_1994), .Q (signal_4743) ) ;
    buf_clk cell_2199 ( .C (clk), .D (signal_3425), .Q (signal_4745) ) ;
    buf_clk cell_2201 ( .C (clk), .D (signal_1989), .Q (signal_4747) ) ;
    buf_clk cell_2203 ( .C (clk), .D (signal_3420), .Q (signal_4749) ) ;
    buf_clk cell_2205 ( .C (clk), .D (signal_2002), .Q (signal_4751) ) ;
    buf_clk cell_2207 ( .C (clk), .D (signal_3433), .Q (signal_4753) ) ;
    buf_clk cell_2209 ( .C (clk), .D (signal_2005), .Q (signal_4755) ) ;
    buf_clk cell_2211 ( .C (clk), .D (signal_3436), .Q (signal_4757) ) ;
    buf_clk cell_2213 ( .C (clk), .D (signal_2006), .Q (signal_4759) ) ;
    buf_clk cell_2215 ( .C (clk), .D (signal_3437), .Q (signal_4761) ) ;
    buf_clk cell_2217 ( .C (clk), .D (signal_2007), .Q (signal_4763) ) ;
    buf_clk cell_2219 ( .C (clk), .D (signal_3438), .Q (signal_4765) ) ;
    buf_clk cell_2221 ( .C (clk), .D (signal_2008), .Q (signal_4767) ) ;
    buf_clk cell_2223 ( .C (clk), .D (signal_3439), .Q (signal_4769) ) ;
    buf_clk cell_2225 ( .C (clk), .D (signal_2009), .Q (signal_4771) ) ;
    buf_clk cell_2227 ( .C (clk), .D (signal_3440), .Q (signal_4773) ) ;
    buf_clk cell_2229 ( .C (clk), .D (signal_2010), .Q (signal_4775) ) ;
    buf_clk cell_2231 ( .C (clk), .D (signal_3441), .Q (signal_4777) ) ;
    buf_clk cell_2233 ( .C (clk), .D (signal_2011), .Q (signal_4779) ) ;
    buf_clk cell_2235 ( .C (clk), .D (signal_3442), .Q (signal_4781) ) ;
    buf_clk cell_2237 ( .C (clk), .D (signal_2000), .Q (signal_4783) ) ;
    buf_clk cell_2239 ( .C (clk), .D (signal_3431), .Q (signal_4785) ) ;
    buf_clk cell_2241 ( .C (clk), .D (signal_4708), .Q (signal_4787) ) ;
    buf_clk cell_2243 ( .C (clk), .D (signal_4710), .Q (signal_4789) ) ;
    buf_clk cell_2245 ( .C (clk), .D (signal_2013), .Q (signal_4791) ) ;
    buf_clk cell_2247 ( .C (clk), .D (signal_3444), .Q (signal_4793) ) ;
    buf_clk cell_2249 ( .C (clk), .D (signal_1990), .Q (signal_4795) ) ;
    buf_clk cell_2251 ( .C (clk), .D (signal_3421), .Q (signal_4797) ) ;
    buf_clk cell_2253 ( .C (clk), .D (signal_4712), .Q (signal_4799) ) ;
    buf_clk cell_2255 ( .C (clk), .D (signal_4714), .Q (signal_4801) ) ;
    buf_clk cell_2257 ( .C (clk), .D (signal_2016), .Q (signal_4803) ) ;
    buf_clk cell_2259 ( .C (clk), .D (signal_3447), .Q (signal_4805) ) ;
    buf_clk cell_2261 ( .C (clk), .D (signal_1992), .Q (signal_4807) ) ;
    buf_clk cell_2263 ( .C (clk), .D (signal_3423), .Q (signal_4809) ) ;
    buf_clk cell_2265 ( .C (clk), .D (signal_2017), .Q (signal_4811) ) ;
    buf_clk cell_2267 ( .C (clk), .D (signal_3448), .Q (signal_4813) ) ;
    buf_clk cell_2269 ( .C (clk), .D (signal_2018), .Q (signal_4815) ) ;
    buf_clk cell_2271 ( .C (clk), .D (signal_3449), .Q (signal_4817) ) ;
    buf_clk cell_2273 ( .C (clk), .D (signal_2015), .Q (signal_4819) ) ;
    buf_clk cell_2275 ( .C (clk), .D (signal_3446), .Q (signal_4821) ) ;
    buf_clk cell_2277 ( .C (clk), .D (signal_2003), .Q (signal_4823) ) ;
    buf_clk cell_2279 ( .C (clk), .D (signal_3434), .Q (signal_4825) ) ;
    buf_clk cell_2281 ( .C (clk), .D (signal_4728), .Q (signal_4827) ) ;
    buf_clk cell_2283 ( .C (clk), .D (signal_4730), .Q (signal_4829) ) ;
    buf_clk cell_2285 ( .C (clk), .D (signal_1997), .Q (signal_4831) ) ;
    buf_clk cell_2287 ( .C (clk), .D (signal_3428), .Q (signal_4833) ) ;
    buf_clk cell_2289 ( .C (clk), .D (signal_4724), .Q (signal_4835) ) ;
    buf_clk cell_2291 ( .C (clk), .D (signal_4726), .Q (signal_4837) ) ;
    buf_clk cell_2293 ( .C (clk), .D (signal_2020), .Q (signal_4839) ) ;
    buf_clk cell_2295 ( .C (clk), .D (signal_3451), .Q (signal_4841) ) ;
    buf_clk cell_2301 ( .C (clk), .D (signal_4846), .Q (signal_4847) ) ;
    buf_clk cell_2309 ( .C (clk), .D (signal_4854), .Q (signal_4855) ) ;
    buf_clk cell_2345 ( .C (clk), .D (signal_4890), .Q (signal_4891) ) ;
    buf_clk cell_2355 ( .C (clk), .D (signal_4900), .Q (signal_4901) ) ;
    buf_clk cell_2365 ( .C (clk), .D (signal_4910), .Q (signal_4911) ) ;
    buf_clk cell_2377 ( .C (clk), .D (signal_4922), .Q (signal_4923) ) ;
    buf_clk cell_2389 ( .C (clk), .D (signal_4934), .Q (signal_4935) ) ;
    buf_clk cell_2405 ( .C (clk), .D (signal_4950), .Q (signal_4951) ) ;
    buf_clk cell_2421 ( .C (clk), .D (signal_4966), .Q (signal_4967) ) ;
    buf_clk cell_2437 ( .C (clk), .D (signal_4982), .Q (signal_4983) ) ;
    buf_clk cell_2453 ( .C (clk), .D (signal_4998), .Q (signal_4999) ) ;
    buf_clk cell_2469 ( .C (clk), .D (signal_5014), .Q (signal_5015) ) ;
    buf_clk cell_2485 ( .C (clk), .D (signal_5030), .Q (signal_5031) ) ;
    buf_clk cell_2501 ( .C (clk), .D (signal_5046), .Q (signal_5047) ) ;
    buf_clk cell_2517 ( .C (clk), .D (signal_5062), .Q (signal_5063) ) ;
    buf_clk cell_2533 ( .C (clk), .D (signal_5078), .Q (signal_5079) ) ;
    buf_clk cell_2549 ( .C (clk), .D (signal_5094), .Q (signal_5095) ) ;
    buf_clk cell_2565 ( .C (clk), .D (signal_5110), .Q (signal_5111) ) ;
    buf_clk cell_2581 ( .C (clk), .D (signal_5126), .Q (signal_5127) ) ;
    buf_clk cell_2597 ( .C (clk), .D (signal_5142), .Q (signal_5143) ) ;
    buf_clk cell_2613 ( .C (clk), .D (signal_5158), .Q (signal_5159) ) ;
    buf_clk cell_2629 ( .C (clk), .D (signal_5174), .Q (signal_5175) ) ;
    buf_clk cell_2645 ( .C (clk), .D (signal_5190), .Q (signal_5191) ) ;
    buf_clk cell_2661 ( .C (clk), .D (signal_5206), .Q (signal_5207) ) ;
    buf_clk cell_2677 ( .C (clk), .D (signal_5222), .Q (signal_5223) ) ;
    buf_clk cell_2693 ( .C (clk), .D (signal_5238), .Q (signal_5239) ) ;
    buf_clk cell_2709 ( .C (clk), .D (signal_5254), .Q (signal_5255) ) ;
    buf_clk cell_2725 ( .C (clk), .D (signal_5270), .Q (signal_5271) ) ;
    buf_clk cell_2741 ( .C (clk), .D (signal_5286), .Q (signal_5287) ) ;
    buf_clk cell_2757 ( .C (clk), .D (signal_5302), .Q (signal_5303) ) ;
    buf_clk cell_2773 ( .C (clk), .D (signal_5318), .Q (signal_5319) ) ;
    buf_clk cell_2789 ( .C (clk), .D (signal_5334), .Q (signal_5335) ) ;
    buf_clk cell_2805 ( .C (clk), .D (signal_5350), .Q (signal_5351) ) ;
    buf_clk cell_2821 ( .C (clk), .D (signal_5366), .Q (signal_5367) ) ;
    buf_clk cell_2837 ( .C (clk), .D (signal_5382), .Q (signal_5383) ) ;
    buf_clk cell_2853 ( .C (clk), .D (signal_5398), .Q (signal_5399) ) ;
    buf_clk cell_2869 ( .C (clk), .D (signal_5414), .Q (signal_5415) ) ;
    buf_clk cell_2885 ( .C (clk), .D (signal_5430), .Q (signal_5431) ) ;
    buf_clk cell_2901 ( .C (clk), .D (signal_5446), .Q (signal_5447) ) ;
    buf_clk cell_2917 ( .C (clk), .D (signal_5462), .Q (signal_5463) ) ;
    buf_clk cell_2933 ( .C (clk), .D (signal_5478), .Q (signal_5479) ) ;
    buf_clk cell_2949 ( .C (clk), .D (signal_5494), .Q (signal_5495) ) ;
    buf_clk cell_2965 ( .C (clk), .D (signal_5510), .Q (signal_5511) ) ;
    buf_clk cell_2981 ( .C (clk), .D (signal_5526), .Q (signal_5527) ) ;
    buf_clk cell_2997 ( .C (clk), .D (signal_5542), .Q (signal_5543) ) ;
    buf_clk cell_3013 ( .C (clk), .D (signal_5558), .Q (signal_5559) ) ;
    buf_clk cell_3029 ( .C (clk), .D (signal_5574), .Q (signal_5575) ) ;
    buf_clk cell_3045 ( .C (clk), .D (signal_5590), .Q (signal_5591) ) ;
    buf_clk cell_3061 ( .C (clk), .D (signal_5606), .Q (signal_5607) ) ;
    buf_clk cell_3077 ( .C (clk), .D (signal_5622), .Q (signal_5623) ) ;
    buf_clk cell_3093 ( .C (clk), .D (signal_5638), .Q (signal_5639) ) ;
    buf_clk cell_3109 ( .C (clk), .D (signal_5654), .Q (signal_5655) ) ;
    buf_clk cell_3125 ( .C (clk), .D (signal_5670), .Q (signal_5671) ) ;
    buf_clk cell_3141 ( .C (clk), .D (signal_5686), .Q (signal_5687) ) ;
    buf_clk cell_3157 ( .C (clk), .D (signal_5702), .Q (signal_5703) ) ;
    buf_clk cell_3173 ( .C (clk), .D (signal_5718), .Q (signal_5719) ) ;
    buf_clk cell_3189 ( .C (clk), .D (signal_5734), .Q (signal_5735) ) ;
    buf_clk cell_3205 ( .C (clk), .D (signal_5750), .Q (signal_5751) ) ;
    buf_clk cell_3221 ( .C (clk), .D (signal_5766), .Q (signal_5767) ) ;
    buf_clk cell_3237 ( .C (clk), .D (signal_5782), .Q (signal_5783) ) ;
    buf_clk cell_3253 ( .C (clk), .D (signal_5798), .Q (signal_5799) ) ;
    buf_clk cell_3269 ( .C (clk), .D (signal_5814), .Q (signal_5815) ) ;
    buf_clk cell_3285 ( .C (clk), .D (signal_5830), .Q (signal_5831) ) ;
    buf_clk cell_3301 ( .C (clk), .D (signal_5846), .Q (signal_5847) ) ;
    buf_clk cell_3317 ( .C (clk), .D (signal_5862), .Q (signal_5863) ) ;
    buf_clk cell_3333 ( .C (clk), .D (signal_5878), .Q (signal_5879) ) ;
    buf_clk cell_3349 ( .C (clk), .D (signal_5894), .Q (signal_5895) ) ;
    buf_clk cell_3365 ( .C (clk), .D (signal_5910), .Q (signal_5911) ) ;
    buf_clk cell_3381 ( .C (clk), .D (signal_5926), .Q (signal_5927) ) ;
    buf_clk cell_3397 ( .C (clk), .D (signal_5942), .Q (signal_5943) ) ;
    buf_clk cell_3413 ( .C (clk), .D (signal_5958), .Q (signal_5959) ) ;
    buf_clk cell_3429 ( .C (clk), .D (signal_5974), .Q (signal_5975) ) ;
    buf_clk cell_3445 ( .C (clk), .D (signal_5990), .Q (signal_5991) ) ;
    buf_clk cell_3461 ( .C (clk), .D (signal_6006), .Q (signal_6007) ) ;
    buf_clk cell_3477 ( .C (clk), .D (signal_6022), .Q (signal_6023) ) ;
    buf_clk cell_3493 ( .C (clk), .D (signal_6038), .Q (signal_6039) ) ;
    buf_clk cell_3509 ( .C (clk), .D (signal_6054), .Q (signal_6055) ) ;
    buf_clk cell_3525 ( .C (clk), .D (signal_6070), .Q (signal_6071) ) ;
    buf_clk cell_3541 ( .C (clk), .D (signal_6086), .Q (signal_6087) ) ;
    buf_clk cell_3557 ( .C (clk), .D (signal_6102), .Q (signal_6103) ) ;
    buf_clk cell_3573 ( .C (clk), .D (signal_6118), .Q (signal_6119) ) ;
    buf_clk cell_3589 ( .C (clk), .D (signal_6134), .Q (signal_6135) ) ;
    buf_clk cell_3605 ( .C (clk), .D (signal_6150), .Q (signal_6151) ) ;
    buf_clk cell_3621 ( .C (clk), .D (signal_6166), .Q (signal_6167) ) ;
    buf_clk cell_3637 ( .C (clk), .D (signal_6182), .Q (signal_6183) ) ;
    buf_clk cell_3653 ( .C (clk), .D (signal_6198), .Q (signal_6199) ) ;
    buf_clk cell_3669 ( .C (clk), .D (signal_6214), .Q (signal_6215) ) ;
    buf_clk cell_3685 ( .C (clk), .D (signal_6230), .Q (signal_6231) ) ;
    buf_clk cell_3701 ( .C (clk), .D (signal_6246), .Q (signal_6247) ) ;
    buf_clk cell_3717 ( .C (clk), .D (signal_6262), .Q (signal_6263) ) ;
    buf_clk cell_3733 ( .C (clk), .D (signal_6278), .Q (signal_6279) ) ;
    buf_clk cell_3749 ( .C (clk), .D (signal_6294), .Q (signal_6295) ) ;
    buf_clk cell_3765 ( .C (clk), .D (signal_6310), .Q (signal_6311) ) ;
    buf_clk cell_3781 ( .C (clk), .D (signal_6326), .Q (signal_6327) ) ;
    buf_clk cell_3797 ( .C (clk), .D (signal_6342), .Q (signal_6343) ) ;
    buf_clk cell_3813 ( .C (clk), .D (signal_6358), .Q (signal_6359) ) ;
    buf_clk cell_3829 ( .C (clk), .D (signal_6374), .Q (signal_6375) ) ;
    buf_clk cell_3845 ( .C (clk), .D (signal_6390), .Q (signal_6391) ) ;
    buf_clk cell_3861 ( .C (clk), .D (signal_6406), .Q (signal_6407) ) ;
    buf_clk cell_3877 ( .C (clk), .D (signal_6422), .Q (signal_6423) ) ;
    buf_clk cell_3893 ( .C (clk), .D (signal_6438), .Q (signal_6439) ) ;
    buf_clk cell_3909 ( .C (clk), .D (signal_6454), .Q (signal_6455) ) ;
    buf_clk cell_3925 ( .C (clk), .D (signal_6470), .Q (signal_6471) ) ;
    buf_clk cell_3941 ( .C (clk), .D (signal_6486), .Q (signal_6487) ) ;
    buf_clk cell_3957 ( .C (clk), .D (signal_6502), .Q (signal_6503) ) ;
    buf_clk cell_3973 ( .C (clk), .D (signal_6518), .Q (signal_6519) ) ;
    buf_clk cell_3989 ( .C (clk), .D (signal_6534), .Q (signal_6535) ) ;
    buf_clk cell_4005 ( .C (clk), .D (signal_6550), .Q (signal_6551) ) ;
    buf_clk cell_4021 ( .C (clk), .D (signal_6566), .Q (signal_6567) ) ;
    buf_clk cell_4037 ( .C (clk), .D (signal_6582), .Q (signal_6583) ) ;
    buf_clk cell_4053 ( .C (clk), .D (signal_6598), .Q (signal_6599) ) ;
    buf_clk cell_4069 ( .C (clk), .D (signal_6614), .Q (signal_6615) ) ;
    buf_clk cell_4085 ( .C (clk), .D (signal_6630), .Q (signal_6631) ) ;
    buf_clk cell_4101 ( .C (clk), .D (signal_6646), .Q (signal_6647) ) ;
    buf_clk cell_4117 ( .C (clk), .D (signal_6662), .Q (signal_6663) ) ;
    buf_clk cell_4133 ( .C (clk), .D (signal_6678), .Q (signal_6679) ) ;
    buf_clk cell_4149 ( .C (clk), .D (signal_6694), .Q (signal_6695) ) ;
    buf_clk cell_4165 ( .C (clk), .D (signal_6710), .Q (signal_6711) ) ;
    buf_clk cell_4181 ( .C (clk), .D (signal_6726), .Q (signal_6727) ) ;
    buf_clk cell_4197 ( .C (clk), .D (signal_6742), .Q (signal_6743) ) ;
    buf_clk cell_4213 ( .C (clk), .D (signal_6758), .Q (signal_6759) ) ;
    buf_clk cell_4229 ( .C (clk), .D (signal_6774), .Q (signal_6775) ) ;
    buf_clk cell_4245 ( .C (clk), .D (signal_6790), .Q (signal_6791) ) ;
    buf_clk cell_4261 ( .C (clk), .D (signal_6806), .Q (signal_6807) ) ;
    buf_clk cell_4277 ( .C (clk), .D (signal_6822), .Q (signal_6823) ) ;
    buf_clk cell_4293 ( .C (clk), .D (signal_6838), .Q (signal_6839) ) ;
    buf_clk cell_4309 ( .C (clk), .D (signal_6854), .Q (signal_6855) ) ;
    buf_clk cell_4325 ( .C (clk), .D (signal_6870), .Q (signal_6871) ) ;
    buf_clk cell_4341 ( .C (clk), .D (signal_6886), .Q (signal_6887) ) ;
    buf_clk cell_4357 ( .C (clk), .D (signal_6902), .Q (signal_6903) ) ;
    buf_clk cell_4373 ( .C (clk), .D (signal_6918), .Q (signal_6919) ) ;
    buf_clk cell_4389 ( .C (clk), .D (signal_6934), .Q (signal_6935) ) ;
    buf_clk cell_4405 ( .C (clk), .D (signal_6950), .Q (signal_6951) ) ;
    buf_clk cell_4419 ( .C (clk), .D (signal_6964), .Q (signal_6965) ) ;
    buf_clk cell_4433 ( .C (clk), .D (signal_6978), .Q (signal_6979) ) ;
    buf_clk cell_4449 ( .C (clk), .D (signal_6994), .Q (signal_6995) ) ;
    buf_clk cell_4465 ( .C (clk), .D (signal_7010), .Q (signal_7011) ) ;
    buf_clk cell_4481 ( .C (clk), .D (signal_7026), .Q (signal_7027) ) ;
    buf_clk cell_4497 ( .C (clk), .D (signal_7042), .Q (signal_7043) ) ;
    buf_clk cell_4513 ( .C (clk), .D (signal_7058), .Q (signal_7059) ) ;
    buf_clk cell_4529 ( .C (clk), .D (signal_7074), .Q (signal_7075) ) ;
    buf_clk cell_4545 ( .C (clk), .D (signal_7090), .Q (signal_7091) ) ;
    buf_clk cell_4561 ( .C (clk), .D (signal_7106), .Q (signal_7107) ) ;
    buf_clk cell_4577 ( .C (clk), .D (signal_7122), .Q (signal_7123) ) ;
    buf_clk cell_4593 ( .C (clk), .D (signal_7138), .Q (signal_7139) ) ;
    buf_clk cell_4609 ( .C (clk), .D (signal_7154), .Q (signal_7155) ) ;
    buf_clk cell_4625 ( .C (clk), .D (signal_7170), .Q (signal_7171) ) ;
    buf_clk cell_4641 ( .C (clk), .D (signal_7186), .Q (signal_7187) ) ;
    buf_clk cell_4657 ( .C (clk), .D (signal_7202), .Q (signal_7203) ) ;
    buf_clk cell_4673 ( .C (clk), .D (signal_7218), .Q (signal_7219) ) ;
    buf_clk cell_4689 ( .C (clk), .D (signal_7234), .Q (signal_7235) ) ;
    buf_clk cell_4705 ( .C (clk), .D (signal_7250), .Q (signal_7251) ) ;
    buf_clk cell_4721 ( .C (clk), .D (signal_7266), .Q (signal_7267) ) ;
    buf_clk cell_4737 ( .C (clk), .D (signal_7282), .Q (signal_7283) ) ;
    buf_clk cell_4753 ( .C (clk), .D (signal_7298), .Q (signal_7299) ) ;
    buf_clk cell_4769 ( .C (clk), .D (signal_7314), .Q (signal_7315) ) ;
    buf_clk cell_4785 ( .C (clk), .D (signal_7330), .Q (signal_7331) ) ;
    buf_clk cell_4801 ( .C (clk), .D (signal_7346), .Q (signal_7347) ) ;
    buf_clk cell_4817 ( .C (clk), .D (signal_7362), .Q (signal_7363) ) ;
    buf_clk cell_4833 ( .C (clk), .D (signal_7378), .Q (signal_7379) ) ;
    buf_clk cell_4849 ( .C (clk), .D (signal_7394), .Q (signal_7395) ) ;
    buf_clk cell_4865 ( .C (clk), .D (signal_7410), .Q (signal_7411) ) ;
    buf_clk cell_4881 ( .C (clk), .D (signal_7426), .Q (signal_7427) ) ;
    buf_clk cell_4897 ( .C (clk), .D (signal_7442), .Q (signal_7443) ) ;
    buf_clk cell_4913 ( .C (clk), .D (signal_7458), .Q (signal_7459) ) ;
    buf_clk cell_4929 ( .C (clk), .D (signal_7474), .Q (signal_7475) ) ;
    buf_clk cell_4945 ( .C (clk), .D (signal_7490), .Q (signal_7491) ) ;
    buf_clk cell_4961 ( .C (clk), .D (signal_7506), .Q (signal_7507) ) ;
    buf_clk cell_4977 ( .C (clk), .D (signal_7522), .Q (signal_7523) ) ;
    buf_clk cell_4993 ( .C (clk), .D (signal_7538), .Q (signal_7539) ) ;
    buf_clk cell_5009 ( .C (clk), .D (signal_7554), .Q (signal_7555) ) ;
    buf_clk cell_5025 ( .C (clk), .D (signal_7570), .Q (signal_7571) ) ;
    buf_clk cell_5041 ( .C (clk), .D (signal_7586), .Q (signal_7587) ) ;
    buf_clk cell_5057 ( .C (clk), .D (signal_7602), .Q (signal_7603) ) ;
    buf_clk cell_5073 ( .C (clk), .D (signal_7618), .Q (signal_7619) ) ;
    buf_clk cell_5089 ( .C (clk), .D (signal_7634), .Q (signal_7635) ) ;
    buf_clk cell_5105 ( .C (clk), .D (signal_7650), .Q (signal_7651) ) ;
    buf_clk cell_5121 ( .C (clk), .D (signal_7666), .Q (signal_7667) ) ;
    buf_clk cell_5137 ( .C (clk), .D (signal_7682), .Q (signal_7683) ) ;
    buf_clk cell_5153 ( .C (clk), .D (signal_7698), .Q (signal_7699) ) ;
    buf_clk cell_5169 ( .C (clk), .D (signal_7714), .Q (signal_7715) ) ;
    buf_clk cell_5185 ( .C (clk), .D (signal_7730), .Q (signal_7731) ) ;
    buf_clk cell_5201 ( .C (clk), .D (signal_7746), .Q (signal_7747) ) ;
    buf_clk cell_5217 ( .C (clk), .D (signal_7762), .Q (signal_7763) ) ;
    buf_clk cell_5233 ( .C (clk), .D (signal_7778), .Q (signal_7779) ) ;
    buf_clk cell_5249 ( .C (clk), .D (signal_7794), .Q (signal_7795) ) ;
    buf_clk cell_5265 ( .C (clk), .D (signal_7810), .Q (signal_7811) ) ;
    buf_clk cell_5281 ( .C (clk), .D (signal_7826), .Q (signal_7827) ) ;
    buf_clk cell_5297 ( .C (clk), .D (signal_7842), .Q (signal_7843) ) ;
    buf_clk cell_5313 ( .C (clk), .D (signal_7858), .Q (signal_7859) ) ;
    buf_clk cell_5329 ( .C (clk), .D (signal_7874), .Q (signal_7875) ) ;
    buf_clk cell_5345 ( .C (clk), .D (signal_7890), .Q (signal_7891) ) ;
    buf_clk cell_5361 ( .C (clk), .D (signal_7906), .Q (signal_7907) ) ;
    buf_clk cell_5377 ( .C (clk), .D (signal_7922), .Q (signal_7923) ) ;
    buf_clk cell_5393 ( .C (clk), .D (signal_7938), .Q (signal_7939) ) ;
    buf_clk cell_5409 ( .C (clk), .D (signal_7954), .Q (signal_7955) ) ;
    buf_clk cell_5425 ( .C (clk), .D (signal_7970), .Q (signal_7971) ) ;
    buf_clk cell_5441 ( .C (clk), .D (signal_7986), .Q (signal_7987) ) ;
    buf_clk cell_5457 ( .C (clk), .D (signal_8002), .Q (signal_8003) ) ;
    buf_clk cell_5473 ( .C (clk), .D (signal_8018), .Q (signal_8019) ) ;
    buf_clk cell_5489 ( .C (clk), .D (signal_8034), .Q (signal_8035) ) ;
    buf_clk cell_5505 ( .C (clk), .D (signal_8050), .Q (signal_8051) ) ;
    buf_clk cell_5521 ( .C (clk), .D (signal_8066), .Q (signal_8067) ) ;
    buf_clk cell_5537 ( .C (clk), .D (signal_8082), .Q (signal_8083) ) ;
    buf_clk cell_5553 ( .C (clk), .D (signal_8098), .Q (signal_8099) ) ;
    buf_clk cell_5569 ( .C (clk), .D (signal_8114), .Q (signal_8115) ) ;
    buf_clk cell_5585 ( .C (clk), .D (signal_8130), .Q (signal_8131) ) ;
    buf_clk cell_5601 ( .C (clk), .D (signal_8146), .Q (signal_8147) ) ;
    buf_clk cell_5617 ( .C (clk), .D (signal_8162), .Q (signal_8163) ) ;
    buf_clk cell_5633 ( .C (clk), .D (signal_8178), .Q (signal_8179) ) ;
    buf_clk cell_5649 ( .C (clk), .D (signal_8194), .Q (signal_8195) ) ;
    buf_clk cell_5665 ( .C (clk), .D (signal_8210), .Q (signal_8211) ) ;
    buf_clk cell_5681 ( .C (clk), .D (signal_8226), .Q (signal_8227) ) ;
    buf_clk cell_5697 ( .C (clk), .D (signal_8242), .Q (signal_8243) ) ;
    buf_clk cell_5713 ( .C (clk), .D (signal_8258), .Q (signal_8259) ) ;
    buf_clk cell_5729 ( .C (clk), .D (signal_8274), .Q (signal_8275) ) ;
    buf_clk cell_5745 ( .C (clk), .D (signal_8290), .Q (signal_8291) ) ;
    buf_clk cell_5761 ( .C (clk), .D (signal_8306), .Q (signal_8307) ) ;
    buf_clk cell_5777 ( .C (clk), .D (signal_8322), .Q (signal_8323) ) ;
    buf_clk cell_5793 ( .C (clk), .D (signal_8338), .Q (signal_8339) ) ;
    buf_clk cell_5809 ( .C (clk), .D (signal_8354), .Q (signal_8355) ) ;
    buf_clk cell_5825 ( .C (clk), .D (signal_8370), .Q (signal_8371) ) ;
    buf_clk cell_5841 ( .C (clk), .D (signal_8386), .Q (signal_8387) ) ;
    buf_clk cell_5857 ( .C (clk), .D (signal_8402), .Q (signal_8403) ) ;
    buf_clk cell_5873 ( .C (clk), .D (signal_8418), .Q (signal_8419) ) ;
    buf_clk cell_5889 ( .C (clk), .D (signal_8434), .Q (signal_8435) ) ;
    buf_clk cell_5905 ( .C (clk), .D (signal_8450), .Q (signal_8451) ) ;
    buf_clk cell_5921 ( .C (clk), .D (signal_8466), .Q (signal_8467) ) ;
    buf_clk cell_5937 ( .C (clk), .D (signal_8482), .Q (signal_8483) ) ;
    buf_clk cell_5953 ( .C (clk), .D (signal_8498), .Q (signal_8499) ) ;
    buf_clk cell_5969 ( .C (clk), .D (signal_8514), .Q (signal_8515) ) ;
    buf_clk cell_5985 ( .C (clk), .D (signal_8530), .Q (signal_8531) ) ;
    buf_clk cell_6001 ( .C (clk), .D (signal_8546), .Q (signal_8547) ) ;
    buf_clk cell_6017 ( .C (clk), .D (signal_8562), .Q (signal_8563) ) ;
    buf_clk cell_6033 ( .C (clk), .D (signal_8578), .Q (signal_8579) ) ;
    buf_clk cell_6049 ( .C (clk), .D (signal_8594), .Q (signal_8595) ) ;
    buf_clk cell_6065 ( .C (clk), .D (signal_8610), .Q (signal_8611) ) ;
    buf_clk cell_6081 ( .C (clk), .D (signal_8626), .Q (signal_8627) ) ;
    buf_clk cell_6097 ( .C (clk), .D (signal_8642), .Q (signal_8643) ) ;
    buf_clk cell_6113 ( .C (clk), .D (signal_8658), .Q (signal_8659) ) ;
    buf_clk cell_6129 ( .C (clk), .D (signal_8674), .Q (signal_8675) ) ;
    buf_clk cell_6145 ( .C (clk), .D (signal_8690), .Q (signal_8691) ) ;
    buf_clk cell_6161 ( .C (clk), .D (signal_8706), .Q (signal_8707) ) ;
    buf_clk cell_6177 ( .C (clk), .D (signal_8722), .Q (signal_8723) ) ;
    buf_clk cell_6193 ( .C (clk), .D (signal_8738), .Q (signal_8739) ) ;
    buf_clk cell_6209 ( .C (clk), .D (signal_8754), .Q (signal_8755) ) ;
    buf_clk cell_6225 ( .C (clk), .D (signal_8770), .Q (signal_8771) ) ;
    buf_clk cell_6241 ( .C (clk), .D (signal_8786), .Q (signal_8787) ) ;
    buf_clk cell_6257 ( .C (clk), .D (signal_8802), .Q (signal_8803) ) ;
    buf_clk cell_6273 ( .C (clk), .D (signal_8818), .Q (signal_8819) ) ;
    buf_clk cell_6289 ( .C (clk), .D (signal_8834), .Q (signal_8835) ) ;
    buf_clk cell_6305 ( .C (clk), .D (signal_8850), .Q (signal_8851) ) ;
    buf_clk cell_6321 ( .C (clk), .D (signal_8866), .Q (signal_8867) ) ;
    buf_clk cell_6337 ( .C (clk), .D (signal_8882), .Q (signal_8883) ) ;
    buf_clk cell_6353 ( .C (clk), .D (signal_8898), .Q (signal_8899) ) ;
    buf_clk cell_6369 ( .C (clk), .D (signal_8914), .Q (signal_8915) ) ;
    buf_clk cell_6385 ( .C (clk), .D (signal_8930), .Q (signal_8931) ) ;
    buf_clk cell_6401 ( .C (clk), .D (signal_8946), .Q (signal_8947) ) ;
    buf_clk cell_6417 ( .C (clk), .D (signal_8962), .Q (signal_8963) ) ;
    buf_clk cell_6433 ( .C (clk), .D (signal_8978), .Q (signal_8979) ) ;
    buf_clk cell_6449 ( .C (clk), .D (signal_8994), .Q (signal_8995) ) ;
    buf_clk cell_6465 ( .C (clk), .D (signal_9010), .Q (signal_9011) ) ;
    buf_clk cell_6481 ( .C (clk), .D (signal_9026), .Q (signal_9027) ) ;
    buf_clk cell_6497 ( .C (clk), .D (signal_9042), .Q (signal_9043) ) ;
    buf_clk cell_6513 ( .C (clk), .D (signal_9058), .Q (signal_9059) ) ;
    buf_clk cell_6529 ( .C (clk), .D (signal_9074), .Q (signal_9075) ) ;
    buf_clk cell_6545 ( .C (clk), .D (signal_9090), .Q (signal_9091) ) ;
    buf_clk cell_6561 ( .C (clk), .D (signal_9106), .Q (signal_9107) ) ;
    buf_clk cell_6577 ( .C (clk), .D (signal_9122), .Q (signal_9123) ) ;
    buf_clk cell_6593 ( .C (clk), .D (signal_9138), .Q (signal_9139) ) ;
    buf_clk cell_6609 ( .C (clk), .D (signal_9154), .Q (signal_9155) ) ;
    buf_clk cell_6625 ( .C (clk), .D (signal_9170), .Q (signal_9171) ) ;
    buf_clk cell_6641 ( .C (clk), .D (signal_9186), .Q (signal_9187) ) ;
    buf_clk cell_6657 ( .C (clk), .D (signal_9202), .Q (signal_9203) ) ;
    buf_clk cell_6673 ( .C (clk), .D (signal_9218), .Q (signal_9219) ) ;
    buf_clk cell_6689 ( .C (clk), .D (signal_9234), .Q (signal_9235) ) ;
    buf_clk cell_6705 ( .C (clk), .D (signal_9250), .Q (signal_9251) ) ;
    buf_clk cell_6721 ( .C (clk), .D (signal_9266), .Q (signal_9267) ) ;
    buf_clk cell_6737 ( .C (clk), .D (signal_9282), .Q (signal_9283) ) ;
    buf_clk cell_6753 ( .C (clk), .D (signal_9298), .Q (signal_9299) ) ;
    buf_clk cell_6769 ( .C (clk), .D (signal_9314), .Q (signal_9315) ) ;
    buf_clk cell_6785 ( .C (clk), .D (signal_9330), .Q (signal_9331) ) ;
    buf_clk cell_6801 ( .C (clk), .D (signal_9346), .Q (signal_9347) ) ;
    buf_clk cell_6817 ( .C (clk), .D (signal_9362), .Q (signal_9363) ) ;
    buf_clk cell_6833 ( .C (clk), .D (signal_9378), .Q (signal_9379) ) ;
    buf_clk cell_6849 ( .C (clk), .D (signal_9394), .Q (signal_9395) ) ;
    buf_clk cell_6865 ( .C (clk), .D (signal_9410), .Q (signal_9411) ) ;
    buf_clk cell_6881 ( .C (clk), .D (signal_9426), .Q (signal_9427) ) ;
    buf_clk cell_6897 ( .C (clk), .D (signal_9442), .Q (signal_9443) ) ;
    buf_clk cell_6913 ( .C (clk), .D (signal_9458), .Q (signal_9459) ) ;
    buf_clk cell_6929 ( .C (clk), .D (signal_9474), .Q (signal_9475) ) ;
    buf_clk cell_6945 ( .C (clk), .D (signal_9490), .Q (signal_9491) ) ;
    buf_clk cell_6961 ( .C (clk), .D (signal_9506), .Q (signal_9507) ) ;
    buf_clk cell_6977 ( .C (clk), .D (signal_9522), .Q (signal_9523) ) ;
    buf_clk cell_6993 ( .C (clk), .D (signal_9538), .Q (signal_9539) ) ;
    buf_clk cell_7009 ( .C (clk), .D (signal_9554), .Q (signal_9555) ) ;
    buf_clk cell_7025 ( .C (clk), .D (signal_9570), .Q (signal_9571) ) ;
    buf_clk cell_7041 ( .C (clk), .D (signal_9586), .Q (signal_9587) ) ;
    buf_clk cell_7057 ( .C (clk), .D (signal_9602), .Q (signal_9603) ) ;
    buf_clk cell_7073 ( .C (clk), .D (signal_9618), .Q (signal_9619) ) ;
    buf_clk cell_7089 ( .C (clk), .D (signal_9634), .Q (signal_9635) ) ;
    buf_clk cell_7105 ( .C (clk), .D (signal_9650), .Q (signal_9651) ) ;
    buf_clk cell_7121 ( .C (clk), .D (signal_9666), .Q (signal_9667) ) ;
    buf_clk cell_7137 ( .C (clk), .D (signal_9682), .Q (signal_9683) ) ;
    buf_clk cell_7153 ( .C (clk), .D (signal_9698), .Q (signal_9699) ) ;
    buf_clk cell_7169 ( .C (clk), .D (signal_9714), .Q (signal_9715) ) ;
    buf_clk cell_7185 ( .C (clk), .D (signal_9730), .Q (signal_9731) ) ;
    buf_clk cell_7201 ( .C (clk), .D (signal_9746), .Q (signal_9747) ) ;
    buf_clk cell_7217 ( .C (clk), .D (signal_9762), .Q (signal_9763) ) ;
    buf_clk cell_7233 ( .C (clk), .D (signal_9778), .Q (signal_9779) ) ;
    buf_clk cell_7249 ( .C (clk), .D (signal_9794), .Q (signal_9795) ) ;
    buf_clk cell_7265 ( .C (clk), .D (signal_9810), .Q (signal_9811) ) ;
    buf_clk cell_7281 ( .C (clk), .D (signal_9826), .Q (signal_9827) ) ;
    buf_clk cell_7297 ( .C (clk), .D (signal_9842), .Q (signal_9843) ) ;
    buf_clk cell_7313 ( .C (clk), .D (signal_9858), .Q (signal_9859) ) ;
    buf_clk cell_7329 ( .C (clk), .D (signal_9874), .Q (signal_9875) ) ;
    buf_clk cell_7345 ( .C (clk), .D (signal_9890), .Q (signal_9891) ) ;
    buf_clk cell_7361 ( .C (clk), .D (signal_9906), .Q (signal_9907) ) ;
    buf_clk cell_7377 ( .C (clk), .D (signal_9922), .Q (signal_9923) ) ;
    buf_clk cell_7393 ( .C (clk), .D (signal_9938), .Q (signal_9939) ) ;
    buf_clk cell_7409 ( .C (clk), .D (signal_9954), .Q (signal_9955) ) ;
    buf_clk cell_7425 ( .C (clk), .D (signal_9970), .Q (signal_9971) ) ;
    buf_clk cell_7441 ( .C (clk), .D (signal_9986), .Q (signal_9987) ) ;
    buf_clk cell_7457 ( .C (clk), .D (signal_10002), .Q (signal_10003) ) ;
    buf_clk cell_7473 ( .C (clk), .D (signal_10018), .Q (signal_10019) ) ;
    buf_clk cell_7489 ( .C (clk), .D (signal_10034), .Q (signal_10035) ) ;
    buf_clk cell_7505 ( .C (clk), .D (signal_10050), .Q (signal_10051) ) ;
    buf_clk cell_7521 ( .C (clk), .D (signal_10066), .Q (signal_10067) ) ;
    buf_clk cell_7537 ( .C (clk), .D (signal_10082), .Q (signal_10083) ) ;
    buf_clk cell_7553 ( .C (clk), .D (signal_10098), .Q (signal_10099) ) ;
    buf_clk cell_7569 ( .C (clk), .D (signal_10114), .Q (signal_10115) ) ;
    buf_clk cell_7585 ( .C (clk), .D (signal_10130), .Q (signal_10131) ) ;
    buf_clk cell_7601 ( .C (clk), .D (signal_10146), .Q (signal_10147) ) ;
    buf_clk cell_7617 ( .C (clk), .D (signal_10162), .Q (signal_10163) ) ;
    buf_clk cell_7633 ( .C (clk), .D (signal_10178), .Q (signal_10179) ) ;
    buf_clk cell_7649 ( .C (clk), .D (signal_10194), .Q (signal_10195) ) ;
    buf_clk cell_7665 ( .C (clk), .D (signal_10210), .Q (signal_10211) ) ;
    buf_clk cell_7681 ( .C (clk), .D (signal_10226), .Q (signal_10227) ) ;
    buf_clk cell_7697 ( .C (clk), .D (signal_10242), .Q (signal_10243) ) ;
    buf_clk cell_7713 ( .C (clk), .D (signal_10258), .Q (signal_10259) ) ;
    buf_clk cell_7729 ( .C (clk), .D (signal_10274), .Q (signal_10275) ) ;
    buf_clk cell_7745 ( .C (clk), .D (signal_10290), .Q (signal_10291) ) ;
    buf_clk cell_7761 ( .C (clk), .D (signal_10306), .Q (signal_10307) ) ;
    buf_clk cell_7777 ( .C (clk), .D (signal_10322), .Q (signal_10323) ) ;
    buf_clk cell_7793 ( .C (clk), .D (signal_10338), .Q (signal_10339) ) ;
    buf_clk cell_7809 ( .C (clk), .D (signal_10354), .Q (signal_10355) ) ;
    buf_clk cell_7825 ( .C (clk), .D (signal_10370), .Q (signal_10371) ) ;
    buf_clk cell_7841 ( .C (clk), .D (signal_10386), .Q (signal_10387) ) ;
    buf_clk cell_7857 ( .C (clk), .D (signal_10402), .Q (signal_10403) ) ;
    buf_clk cell_7873 ( .C (clk), .D (signal_10418), .Q (signal_10419) ) ;
    buf_clk cell_7889 ( .C (clk), .D (signal_10434), .Q (signal_10435) ) ;
    buf_clk cell_7905 ( .C (clk), .D (signal_10450), .Q (signal_10451) ) ;
    buf_clk cell_7921 ( .C (clk), .D (signal_10466), .Q (signal_10467) ) ;
    buf_clk cell_7937 ( .C (clk), .D (signal_10482), .Q (signal_10483) ) ;
    buf_clk cell_7953 ( .C (clk), .D (signal_10498), .Q (signal_10499) ) ;
    buf_clk cell_7969 ( .C (clk), .D (signal_10514), .Q (signal_10515) ) ;
    buf_clk cell_7985 ( .C (clk), .D (signal_10530), .Q (signal_10531) ) ;
    buf_clk cell_8001 ( .C (clk), .D (signal_10546), .Q (signal_10547) ) ;
    buf_clk cell_8017 ( .C (clk), .D (signal_10562), .Q (signal_10563) ) ;
    buf_clk cell_8033 ( .C (clk), .D (signal_10578), .Q (signal_10579) ) ;
    buf_clk cell_8049 ( .C (clk), .D (signal_10594), .Q (signal_10595) ) ;
    buf_clk cell_8065 ( .C (clk), .D (signal_10610), .Q (signal_10611) ) ;
    buf_clk cell_8081 ( .C (clk), .D (signal_10626), .Q (signal_10627) ) ;
    buf_clk cell_8097 ( .C (clk), .D (signal_10642), .Q (signal_10643) ) ;
    buf_clk cell_8113 ( .C (clk), .D (signal_10658), .Q (signal_10659) ) ;
    buf_clk cell_8129 ( .C (clk), .D (signal_10674), .Q (signal_10675) ) ;
    buf_clk cell_8145 ( .C (clk), .D (signal_10690), .Q (signal_10691) ) ;
    buf_clk cell_8161 ( .C (clk), .D (signal_10706), .Q (signal_10707) ) ;
    buf_clk cell_8177 ( .C (clk), .D (signal_10722), .Q (signal_10723) ) ;
    buf_clk cell_8193 ( .C (clk), .D (signal_10738), .Q (signal_10739) ) ;
    buf_clk cell_8209 ( .C (clk), .D (signal_10754), .Q (signal_10755) ) ;
    buf_clk cell_8225 ( .C (clk), .D (signal_10770), .Q (signal_10771) ) ;
    buf_clk cell_8241 ( .C (clk), .D (signal_10786), .Q (signal_10787) ) ;
    buf_clk cell_8257 ( .C (clk), .D (signal_10802), .Q (signal_10803) ) ;
    buf_clk cell_8273 ( .C (clk), .D (signal_10818), .Q (signal_10819) ) ;
    buf_clk cell_8289 ( .C (clk), .D (signal_10834), .Q (signal_10835) ) ;
    buf_clk cell_8305 ( .C (clk), .D (signal_10850), .Q (signal_10851) ) ;
    buf_clk cell_8321 ( .C (clk), .D (signal_10866), .Q (signal_10867) ) ;
    buf_clk cell_8337 ( .C (clk), .D (signal_10882), .Q (signal_10883) ) ;
    buf_clk cell_8353 ( .C (clk), .D (signal_10898), .Q (signal_10899) ) ;
    buf_clk cell_8369 ( .C (clk), .D (signal_10914), .Q (signal_10915) ) ;
    buf_clk cell_8385 ( .C (clk), .D (signal_10930), .Q (signal_10931) ) ;
    buf_clk cell_8401 ( .C (clk), .D (signal_10946), .Q (signal_10947) ) ;
    buf_clk cell_8417 ( .C (clk), .D (signal_10962), .Q (signal_10963) ) ;
    buf_clk cell_8433 ( .C (clk), .D (signal_10978), .Q (signal_10979) ) ;
    buf_clk cell_8449 ( .C (clk), .D (signal_10994), .Q (signal_10995) ) ;
    buf_clk cell_8465 ( .C (clk), .D (signal_11010), .Q (signal_11011) ) ;
    buf_clk cell_8481 ( .C (clk), .D (signal_11026), .Q (signal_11027) ) ;
    buf_clk cell_8497 ( .C (clk), .D (signal_11042), .Q (signal_11043) ) ;
    buf_clk cell_8513 ( .C (clk), .D (signal_11058), .Q (signal_11059) ) ;
    buf_clk cell_8529 ( .C (clk), .D (signal_11074), .Q (signal_11075) ) ;
    buf_clk cell_8545 ( .C (clk), .D (signal_11090), .Q (signal_11091) ) ;
    buf_clk cell_8561 ( .C (clk), .D (signal_11106), .Q (signal_11107) ) ;
    buf_clk cell_8577 ( .C (clk), .D (signal_11122), .Q (signal_11123) ) ;
    buf_clk cell_8593 ( .C (clk), .D (signal_11138), .Q (signal_11139) ) ;
    buf_clk cell_8609 ( .C (clk), .D (signal_11154), .Q (signal_11155) ) ;
    buf_clk cell_8625 ( .C (clk), .D (signal_11170), .Q (signal_11171) ) ;
    buf_clk cell_8641 ( .C (clk), .D (signal_11186), .Q (signal_11187) ) ;
    buf_clk cell_8657 ( .C (clk), .D (signal_11202), .Q (signal_11203) ) ;
    buf_clk cell_8673 ( .C (clk), .D (signal_11218), .Q (signal_11219) ) ;
    buf_clk cell_8689 ( .C (clk), .D (signal_11234), .Q (signal_11235) ) ;
    buf_clk cell_8705 ( .C (clk), .D (signal_11250), .Q (signal_11251) ) ;
    buf_clk cell_8721 ( .C (clk), .D (signal_11266), .Q (signal_11267) ) ;
    buf_clk cell_8737 ( .C (clk), .D (signal_11282), .Q (signal_11283) ) ;
    buf_clk cell_8753 ( .C (clk), .D (signal_11298), .Q (signal_11299) ) ;
    buf_clk cell_8769 ( .C (clk), .D (signal_11314), .Q (signal_11315) ) ;
    buf_clk cell_8785 ( .C (clk), .D (signal_11330), .Q (signal_11331) ) ;
    buf_clk cell_8801 ( .C (clk), .D (signal_11346), .Q (signal_11347) ) ;
    buf_clk cell_8817 ( .C (clk), .D (signal_11362), .Q (signal_11363) ) ;
    buf_clk cell_8833 ( .C (clk), .D (signal_11378), .Q (signal_11379) ) ;
    buf_clk cell_8849 ( .C (clk), .D (signal_11394), .Q (signal_11395) ) ;
    buf_clk cell_8865 ( .C (clk), .D (signal_11410), .Q (signal_11411) ) ;
    buf_clk cell_8881 ( .C (clk), .D (signal_11426), .Q (signal_11427) ) ;
    buf_clk cell_8897 ( .C (clk), .D (signal_11442), .Q (signal_11443) ) ;
    buf_clk cell_8913 ( .C (clk), .D (signal_11458), .Q (signal_11459) ) ;
    buf_clk cell_8929 ( .C (clk), .D (signal_11474), .Q (signal_11475) ) ;
    buf_clk cell_8945 ( .C (clk), .D (signal_11490), .Q (signal_11491) ) ;
    buf_clk cell_8961 ( .C (clk), .D (signal_11506), .Q (signal_11507) ) ;
    buf_clk cell_8977 ( .C (clk), .D (signal_11522), .Q (signal_11523) ) ;
    buf_clk cell_8993 ( .C (clk), .D (signal_11538), .Q (signal_11539) ) ;
    buf_clk cell_9009 ( .C (clk), .D (signal_11554), .Q (signal_11555) ) ;
    buf_clk cell_9025 ( .C (clk), .D (signal_11570), .Q (signal_11571) ) ;
    buf_clk cell_9041 ( .C (clk), .D (signal_11586), .Q (signal_11587) ) ;
    buf_clk cell_9057 ( .C (clk), .D (signal_11602), .Q (signal_11603) ) ;
    buf_clk cell_9073 ( .C (clk), .D (signal_11618), .Q (signal_11619) ) ;
    buf_clk cell_9089 ( .C (clk), .D (signal_11634), .Q (signal_11635) ) ;
    buf_clk cell_9105 ( .C (clk), .D (signal_11650), .Q (signal_11651) ) ;
    buf_clk cell_9121 ( .C (clk), .D (signal_11666), .Q (signal_11667) ) ;
    buf_clk cell_9137 ( .C (clk), .D (signal_11682), .Q (signal_11683) ) ;
    buf_clk cell_9153 ( .C (clk), .D (signal_11698), .Q (signal_11699) ) ;
    buf_clk cell_9169 ( .C (clk), .D (signal_11714), .Q (signal_11715) ) ;
    buf_clk cell_9185 ( .C (clk), .D (signal_11730), .Q (signal_11731) ) ;
    buf_clk cell_9201 ( .C (clk), .D (signal_11746), .Q (signal_11747) ) ;
    buf_clk cell_9217 ( .C (clk), .D (signal_11762), .Q (signal_11763) ) ;
    buf_clk cell_9233 ( .C (clk), .D (signal_11778), .Q (signal_11779) ) ;
    buf_clk cell_9249 ( .C (clk), .D (signal_11794), .Q (signal_11795) ) ;
    buf_clk cell_9265 ( .C (clk), .D (signal_11810), .Q (signal_11811) ) ;
    buf_clk cell_9281 ( .C (clk), .D (signal_11826), .Q (signal_11827) ) ;
    buf_clk cell_9297 ( .C (clk), .D (signal_11842), .Q (signal_11843) ) ;
    buf_clk cell_9313 ( .C (clk), .D (signal_11858), .Q (signal_11859) ) ;
    buf_clk cell_9329 ( .C (clk), .D (signal_11874), .Q (signal_11875) ) ;
    buf_clk cell_9345 ( .C (clk), .D (signal_11890), .Q (signal_11891) ) ;
    buf_clk cell_9361 ( .C (clk), .D (signal_11906), .Q (signal_11907) ) ;
    buf_clk cell_9377 ( .C (clk), .D (signal_11922), .Q (signal_11923) ) ;
    buf_clk cell_9393 ( .C (clk), .D (signal_11938), .Q (signal_11939) ) ;
    buf_clk cell_9409 ( .C (clk), .D (signal_11954), .Q (signal_11955) ) ;
    buf_clk cell_9425 ( .C (clk), .D (signal_11970), .Q (signal_11971) ) ;
    buf_clk cell_9441 ( .C (clk), .D (signal_11986), .Q (signal_11987) ) ;
    buf_clk cell_9457 ( .C (clk), .D (signal_12002), .Q (signal_12003) ) ;
    buf_clk cell_9473 ( .C (clk), .D (signal_12018), .Q (signal_12019) ) ;
    buf_clk cell_9489 ( .C (clk), .D (signal_12034), .Q (signal_12035) ) ;
    buf_clk cell_9505 ( .C (clk), .D (signal_12050), .Q (signal_12051) ) ;
    buf_clk cell_9521 ( .C (clk), .D (signal_12066), .Q (signal_12067) ) ;
    buf_clk cell_9537 ( .C (clk), .D (signal_12082), .Q (signal_12083) ) ;
    buf_clk cell_9553 ( .C (clk), .D (signal_12098), .Q (signal_12099) ) ;
    buf_clk cell_9569 ( .C (clk), .D (signal_12114), .Q (signal_12115) ) ;
    buf_clk cell_9585 ( .C (clk), .D (signal_12130), .Q (signal_12131) ) ;
    buf_clk cell_9601 ( .C (clk), .D (signal_12146), .Q (signal_12147) ) ;
    buf_clk cell_9617 ( .C (clk), .D (signal_12162), .Q (signal_12163) ) ;
    buf_clk cell_9633 ( .C (clk), .D (signal_12178), .Q (signal_12179) ) ;
    buf_clk cell_9649 ( .C (clk), .D (signal_12194), .Q (signal_12195) ) ;
    buf_clk cell_9665 ( .C (clk), .D (signal_12210), .Q (signal_12211) ) ;
    buf_clk cell_9681 ( .C (clk), .D (signal_12226), .Q (signal_12227) ) ;
    buf_clk cell_9697 ( .C (clk), .D (signal_12242), .Q (signal_12243) ) ;
    buf_clk cell_9713 ( .C (clk), .D (signal_12258), .Q (signal_12259) ) ;
    buf_clk cell_9729 ( .C (clk), .D (signal_12274), .Q (signal_12275) ) ;
    buf_clk cell_9745 ( .C (clk), .D (signal_12290), .Q (signal_12291) ) ;
    buf_clk cell_9761 ( .C (clk), .D (signal_12306), .Q (signal_12307) ) ;
    buf_clk cell_9777 ( .C (clk), .D (signal_12322), .Q (signal_12323) ) ;
    buf_clk cell_9793 ( .C (clk), .D (signal_12338), .Q (signal_12339) ) ;
    buf_clk cell_9809 ( .C (clk), .D (signal_12354), .Q (signal_12355) ) ;
    buf_clk cell_9825 ( .C (clk), .D (signal_12370), .Q (signal_12371) ) ;
    buf_clk cell_9841 ( .C (clk), .D (signal_12386), .Q (signal_12387) ) ;
    buf_clk cell_9857 ( .C (clk), .D (signal_12402), .Q (signal_12403) ) ;
    buf_clk cell_9873 ( .C (clk), .D (signal_12418), .Q (signal_12419) ) ;
    buf_clk cell_9889 ( .C (clk), .D (signal_12434), .Q (signal_12435) ) ;
    buf_clk cell_9905 ( .C (clk), .D (signal_12450), .Q (signal_12451) ) ;
    buf_clk cell_9921 ( .C (clk), .D (signal_12466), .Q (signal_12467) ) ;
    buf_clk cell_9937 ( .C (clk), .D (signal_12482), .Q (signal_12483) ) ;
    buf_clk cell_9953 ( .C (clk), .D (signal_12498), .Q (signal_12499) ) ;
    buf_clk cell_9969 ( .C (clk), .D (signal_12514), .Q (signal_12515) ) ;
    buf_clk cell_9985 ( .C (clk), .D (signal_12530), .Q (signal_12531) ) ;
    buf_clk cell_10001 ( .C (clk), .D (signal_12546), .Q (signal_12547) ) ;
    buf_clk cell_10017 ( .C (clk), .D (signal_12562), .Q (signal_12563) ) ;
    buf_clk cell_10033 ( .C (clk), .D (signal_12578), .Q (signal_12579) ) ;
    buf_clk cell_10049 ( .C (clk), .D (signal_12594), .Q (signal_12595) ) ;
    buf_clk cell_10065 ( .C (clk), .D (signal_12610), .Q (signal_12611) ) ;
    buf_clk cell_10081 ( .C (clk), .D (signal_12626), .Q (signal_12627) ) ;
    buf_clk cell_10097 ( .C (clk), .D (signal_12642), .Q (signal_12643) ) ;
    buf_clk cell_10113 ( .C (clk), .D (signal_12658), .Q (signal_12659) ) ;
    buf_clk cell_10129 ( .C (clk), .D (signal_12674), .Q (signal_12675) ) ;
    buf_clk cell_10145 ( .C (clk), .D (signal_12690), .Q (signal_12691) ) ;
    buf_clk cell_10161 ( .C (clk), .D (signal_12706), .Q (signal_12707) ) ;
    buf_clk cell_10177 ( .C (clk), .D (signal_12722), .Q (signal_12723) ) ;
    buf_clk cell_10193 ( .C (clk), .D (signal_12738), .Q (signal_12739) ) ;
    buf_clk cell_10209 ( .C (clk), .D (signal_12754), .Q (signal_12755) ) ;
    buf_clk cell_10225 ( .C (clk), .D (signal_12770), .Q (signal_12771) ) ;
    buf_clk cell_10241 ( .C (clk), .D (signal_12786), .Q (signal_12787) ) ;
    buf_clk cell_10257 ( .C (clk), .D (signal_12802), .Q (signal_12803) ) ;
    buf_clk cell_10273 ( .C (clk), .D (signal_12818), .Q (signal_12819) ) ;
    buf_clk cell_10289 ( .C (clk), .D (signal_12834), .Q (signal_12835) ) ;
    buf_clk cell_10305 ( .C (clk), .D (signal_12850), .Q (signal_12851) ) ;
    buf_clk cell_10321 ( .C (clk), .D (signal_12866), .Q (signal_12867) ) ;
    buf_clk cell_10337 ( .C (clk), .D (signal_12882), .Q (signal_12883) ) ;
    buf_clk cell_10353 ( .C (clk), .D (signal_12898), .Q (signal_12899) ) ;
    buf_clk cell_10369 ( .C (clk), .D (signal_12914), .Q (signal_12915) ) ;
    buf_clk cell_10385 ( .C (clk), .D (signal_12930), .Q (signal_12931) ) ;
    buf_clk cell_10401 ( .C (clk), .D (signal_12946), .Q (signal_12947) ) ;
    buf_clk cell_10417 ( .C (clk), .D (signal_12962), .Q (signal_12963) ) ;
    buf_clk cell_10433 ( .C (clk), .D (signal_12978), .Q (signal_12979) ) ;
    buf_clk cell_10449 ( .C (clk), .D (signal_12994), .Q (signal_12995) ) ;
    buf_clk cell_10465 ( .C (clk), .D (signal_13010), .Q (signal_13011) ) ;
    buf_clk cell_10481 ( .C (clk), .D (signal_13026), .Q (signal_13027) ) ;
    buf_clk cell_10497 ( .C (clk), .D (signal_13042), .Q (signal_13043) ) ;
    buf_clk cell_10513 ( .C (clk), .D (signal_13058), .Q (signal_13059) ) ;
    buf_clk cell_10529 ( .C (clk), .D (signal_13074), .Q (signal_13075) ) ;
    buf_clk cell_10545 ( .C (clk), .D (signal_13090), .Q (signal_13091) ) ;
    buf_clk cell_10561 ( .C (clk), .D (signal_13106), .Q (signal_13107) ) ;
    buf_clk cell_10577 ( .C (clk), .D (signal_13122), .Q (signal_13123) ) ;
    buf_clk cell_10593 ( .C (clk), .D (signal_13138), .Q (signal_13139) ) ;
    buf_clk cell_10609 ( .C (clk), .D (signal_13154), .Q (signal_13155) ) ;
    buf_clk cell_10625 ( .C (clk), .D (signal_13170), .Q (signal_13171) ) ;
    buf_clk cell_10641 ( .C (clk), .D (signal_13186), .Q (signal_13187) ) ;
    buf_clk cell_10657 ( .C (clk), .D (signal_13202), .Q (signal_13203) ) ;
    buf_clk cell_10673 ( .C (clk), .D (signal_13218), .Q (signal_13219) ) ;
    buf_clk cell_10689 ( .C (clk), .D (signal_13234), .Q (signal_13235) ) ;
    buf_clk cell_10705 ( .C (clk), .D (signal_13250), .Q (signal_13251) ) ;
    buf_clk cell_10721 ( .C (clk), .D (signal_13266), .Q (signal_13267) ) ;
    buf_clk cell_10737 ( .C (clk), .D (signal_13282), .Q (signal_13283) ) ;
    buf_clk cell_10753 ( .C (clk), .D (signal_13298), .Q (signal_13299) ) ;
    buf_clk cell_10769 ( .C (clk), .D (signal_13314), .Q (signal_13315) ) ;
    buf_clk cell_10785 ( .C (clk), .D (signal_13330), .Q (signal_13331) ) ;
    buf_clk cell_10801 ( .C (clk), .D (signal_13346), .Q (signal_13347) ) ;
    buf_clk cell_10817 ( .C (clk), .D (signal_13362), .Q (signal_13363) ) ;
    buf_clk cell_10833 ( .C (clk), .D (signal_13378), .Q (signal_13379) ) ;
    buf_clk cell_10849 ( .C (clk), .D (signal_13394), .Q (signal_13395) ) ;
    buf_clk cell_10865 ( .C (clk), .D (signal_13410), .Q (signal_13411) ) ;
    buf_clk cell_10881 ( .C (clk), .D (signal_13426), .Q (signal_13427) ) ;
    buf_clk cell_10897 ( .C (clk), .D (signal_13442), .Q (signal_13443) ) ;
    buf_clk cell_10913 ( .C (clk), .D (signal_13458), .Q (signal_13459) ) ;
    buf_clk cell_10929 ( .C (clk), .D (signal_13474), .Q (signal_13475) ) ;
    buf_clk cell_10945 ( .C (clk), .D (signal_13490), .Q (signal_13491) ) ;
    buf_clk cell_10961 ( .C (clk), .D (signal_13506), .Q (signal_13507) ) ;
    buf_clk cell_10977 ( .C (clk), .D (signal_13522), .Q (signal_13523) ) ;
    buf_clk cell_10993 ( .C (clk), .D (signal_13538), .Q (signal_13539) ) ;
    buf_clk cell_11009 ( .C (clk), .D (signal_13554), .Q (signal_13555) ) ;
    buf_clk cell_11025 ( .C (clk), .D (signal_13570), .Q (signal_13571) ) ;
    buf_clk cell_11041 ( .C (clk), .D (signal_13586), .Q (signal_13587) ) ;
    buf_clk cell_11057 ( .C (clk), .D (signal_13602), .Q (signal_13603) ) ;
    buf_clk cell_11073 ( .C (clk), .D (signal_13618), .Q (signal_13619) ) ;
    buf_clk cell_11089 ( .C (clk), .D (signal_13634), .Q (signal_13635) ) ;
    buf_clk cell_11105 ( .C (clk), .D (signal_13650), .Q (signal_13651) ) ;
    buf_clk cell_11121 ( .C (clk), .D (signal_13666), .Q (signal_13667) ) ;
    buf_clk cell_11137 ( .C (clk), .D (signal_13682), .Q (signal_13683) ) ;
    buf_clk cell_11153 ( .C (clk), .D (signal_13698), .Q (signal_13699) ) ;
    buf_clk cell_11169 ( .C (clk), .D (signal_13714), .Q (signal_13715) ) ;
    buf_clk cell_11185 ( .C (clk), .D (signal_13730), .Q (signal_13731) ) ;
    buf_clk cell_11201 ( .C (clk), .D (signal_13746), .Q (signal_13747) ) ;
    buf_clk cell_11217 ( .C (clk), .D (signal_13762), .Q (signal_13763) ) ;
    buf_clk cell_11233 ( .C (clk), .D (signal_13778), .Q (signal_13779) ) ;
    buf_clk cell_11249 ( .C (clk), .D (signal_13794), .Q (signal_13795) ) ;
    buf_clk cell_11265 ( .C (clk), .D (signal_13810), .Q (signal_13811) ) ;
    buf_clk cell_11281 ( .C (clk), .D (signal_13826), .Q (signal_13827) ) ;
    buf_clk cell_11297 ( .C (clk), .D (signal_13842), .Q (signal_13843) ) ;
    buf_clk cell_11313 ( .C (clk), .D (signal_13858), .Q (signal_13859) ) ;
    buf_clk cell_11329 ( .C (clk), .D (signal_13874), .Q (signal_13875) ) ;
    buf_clk cell_11345 ( .C (clk), .D (signal_13890), .Q (signal_13891) ) ;
    buf_clk cell_11361 ( .C (clk), .D (signal_13906), .Q (signal_13907) ) ;
    buf_clk cell_11377 ( .C (clk), .D (signal_13922), .Q (signal_13923) ) ;
    buf_clk cell_11393 ( .C (clk), .D (signal_13938), .Q (signal_13939) ) ;
    buf_clk cell_11409 ( .C (clk), .D (signal_13954), .Q (signal_13955) ) ;
    buf_clk cell_11425 ( .C (clk), .D (signal_13970), .Q (signal_13971) ) ;
    buf_clk cell_11441 ( .C (clk), .D (signal_13986), .Q (signal_13987) ) ;
    buf_clk cell_11457 ( .C (clk), .D (signal_14002), .Q (signal_14003) ) ;
    buf_clk cell_11473 ( .C (clk), .D (signal_14018), .Q (signal_14019) ) ;
    buf_clk cell_11489 ( .C (clk), .D (signal_14034), .Q (signal_14035) ) ;
    buf_clk cell_11505 ( .C (clk), .D (signal_14050), .Q (signal_14051) ) ;
    buf_clk cell_11521 ( .C (clk), .D (signal_14066), .Q (signal_14067) ) ;
    buf_clk cell_11537 ( .C (clk), .D (signal_14082), .Q (signal_14083) ) ;
    buf_clk cell_11553 ( .C (clk), .D (signal_14098), .Q (signal_14099) ) ;
    buf_clk cell_11569 ( .C (clk), .D (signal_14114), .Q (signal_14115) ) ;
    buf_clk cell_11585 ( .C (clk), .D (signal_14130), .Q (signal_14131) ) ;
    buf_clk cell_11601 ( .C (clk), .D (signal_14146), .Q (signal_14147) ) ;
    buf_clk cell_11617 ( .C (clk), .D (signal_14162), .Q (signal_14163) ) ;
    buf_clk cell_11633 ( .C (clk), .D (signal_14178), .Q (signal_14179) ) ;
    buf_clk cell_11649 ( .C (clk), .D (signal_14194), .Q (signal_14195) ) ;
    buf_clk cell_11665 ( .C (clk), .D (signal_14210), .Q (signal_14211) ) ;
    buf_clk cell_11681 ( .C (clk), .D (signal_14226), .Q (signal_14227) ) ;
    buf_clk cell_11697 ( .C (clk), .D (signal_14242), .Q (signal_14243) ) ;
    buf_clk cell_11713 ( .C (clk), .D (signal_14258), .Q (signal_14259) ) ;
    buf_clk cell_11729 ( .C (clk), .D (signal_14274), .Q (signal_14275) ) ;
    buf_clk cell_11745 ( .C (clk), .D (signal_14290), .Q (signal_14291) ) ;
    buf_clk cell_11761 ( .C (clk), .D (signal_14306), .Q (signal_14307) ) ;
    buf_clk cell_11777 ( .C (clk), .D (signal_14322), .Q (signal_14323) ) ;
    buf_clk cell_11793 ( .C (clk), .D (signal_14338), .Q (signal_14339) ) ;
    buf_clk cell_11809 ( .C (clk), .D (signal_14354), .Q (signal_14355) ) ;
    buf_clk cell_11825 ( .C (clk), .D (signal_14370), .Q (signal_14371) ) ;
    buf_clk cell_11841 ( .C (clk), .D (signal_14386), .Q (signal_14387) ) ;
    buf_clk cell_11857 ( .C (clk), .D (signal_14402), .Q (signal_14403) ) ;
    buf_clk cell_11873 ( .C (clk), .D (signal_14418), .Q (signal_14419) ) ;
    buf_clk cell_11889 ( .C (clk), .D (signal_14434), .Q (signal_14435) ) ;
    buf_clk cell_11905 ( .C (clk), .D (signal_14450), .Q (signal_14451) ) ;
    buf_clk cell_11921 ( .C (clk), .D (signal_14466), .Q (signal_14467) ) ;
    buf_clk cell_11937 ( .C (clk), .D (signal_14482), .Q (signal_14483) ) ;
    buf_clk cell_11953 ( .C (clk), .D (signal_14498), .Q (signal_14499) ) ;
    buf_clk cell_11969 ( .C (clk), .D (signal_14514), .Q (signal_14515) ) ;
    buf_clk cell_11985 ( .C (clk), .D (signal_14530), .Q (signal_14531) ) ;
    buf_clk cell_12001 ( .C (clk), .D (signal_14546), .Q (signal_14547) ) ;
    buf_clk cell_12017 ( .C (clk), .D (signal_14562), .Q (signal_14563) ) ;
    buf_clk cell_12033 ( .C (clk), .D (signal_14578), .Q (signal_14579) ) ;
    buf_clk cell_12049 ( .C (clk), .D (signal_14594), .Q (signal_14595) ) ;
    buf_clk cell_12065 ( .C (clk), .D (signal_14610), .Q (signal_14611) ) ;
    buf_clk cell_12081 ( .C (clk), .D (signal_14626), .Q (signal_14627) ) ;
    buf_clk cell_12097 ( .C (clk), .D (signal_14642), .Q (signal_14643) ) ;
    buf_clk cell_12113 ( .C (clk), .D (signal_14658), .Q (signal_14659) ) ;
    buf_clk cell_12129 ( .C (clk), .D (signal_14674), .Q (signal_14675) ) ;
    buf_clk cell_12145 ( .C (clk), .D (signal_14690), .Q (signal_14691) ) ;
    buf_clk cell_12161 ( .C (clk), .D (signal_14706), .Q (signal_14707) ) ;
    buf_clk cell_12177 ( .C (clk), .D (signal_14722), .Q (signal_14723) ) ;
    buf_clk cell_12193 ( .C (clk), .D (signal_14738), .Q (signal_14739) ) ;
    buf_clk cell_12209 ( .C (clk), .D (signal_14754), .Q (signal_14755) ) ;
    buf_clk cell_12225 ( .C (clk), .D (signal_14770), .Q (signal_14771) ) ;
    buf_clk cell_12241 ( .C (clk), .D (signal_14786), .Q (signal_14787) ) ;
    buf_clk cell_12257 ( .C (clk), .D (signal_14802), .Q (signal_14803) ) ;
    buf_clk cell_12273 ( .C (clk), .D (signal_14818), .Q (signal_14819) ) ;
    buf_clk cell_12289 ( .C (clk), .D (signal_14834), .Q (signal_14835) ) ;
    buf_clk cell_12305 ( .C (clk), .D (signal_14850), .Q (signal_14851) ) ;
    buf_clk cell_12321 ( .C (clk), .D (signal_14866), .Q (signal_14867) ) ;
    buf_clk cell_12337 ( .C (clk), .D (signal_14882), .Q (signal_14883) ) ;
    buf_clk cell_12353 ( .C (clk), .D (signal_14898), .Q (signal_14899) ) ;
    buf_clk cell_12369 ( .C (clk), .D (signal_14914), .Q (signal_14915) ) ;
    buf_clk cell_12385 ( .C (clk), .D (signal_14930), .Q (signal_14931) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1753 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[39]), .c ({signal_3476, signal_2021}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1754 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[40]), .c ({signal_3477, signal_2022}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1755 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[41]), .c ({signal_3478, signal_2023}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1756 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[42]), .c ({signal_3479, signal_2024}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1757 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[43]), .c ({signal_3480, signal_2025}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1758 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[44]), .c ({signal_3481, signal_2026}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1759 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[45]), .c ({signal_3482, signal_2027}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1760 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[46]), .c ({signal_3483, signal_2028}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1761 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[47]), .c ({signal_3484, signal_2029}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1762 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[48]), .c ({signal_3485, signal_2030}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1763 ( .s ({signal_4702, signal_4700}), .b ({signal_4710, signal_4708}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[49]), .c ({signal_3486, signal_2031}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1764 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[50]), .c ({signal_3487, signal_2032}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1765 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[51]), .c ({signal_3488, signal_2033}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1766 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[52]), .c ({signal_3489, signal_2034}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1767 ( .s ({signal_4722, signal_4718}), .b ({signal_3430, signal_1999}), .a ({signal_3429, signal_1998}), .clk (clk), .r (Fresh[53]), .c ({signal_3490, signal_2035}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1768 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[54]), .c ({signal_3491, signal_2036}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1769 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[55]), .c ({signal_3492, signal_2037}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1770 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[56]), .c ({signal_3493, signal_2038}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1771 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[57]), .c ({signal_3494, signal_2039}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1772 ( .s ({signal_4722, signal_4718}), .b ({signal_3432, signal_2001}), .a ({signal_3431, signal_2000}), .clk (clk), .r (Fresh[58]), .c ({signal_3495, signal_2040}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1773 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[59]), .c ({signal_3496, signal_2041}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1774 ( .s ({signal_4722, signal_4718}), .b ({signal_3435, signal_2004}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[60]), .c ({signal_3497, signal_2042}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1775 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[61]), .c ({signal_3498, signal_2043}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1776 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[62]), .c ({signal_3499, signal_2044}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1777 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[63]), .c ({signal_3500, signal_2045}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1778 ( .s ({signal_4702, signal_4700}), .b ({signal_4710, signal_4708}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[64]), .c ({signal_3501, signal_2046}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1779 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[65]), .c ({signal_3502, signal_2047}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1780 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[66]), .c ({signal_3503, signal_2048}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1781 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[67]), .c ({signal_3504, signal_2049}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1782 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[68]), .c ({signal_3505, signal_2050}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1783 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[69]), .c ({signal_3506, signal_2051}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1784 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[70]), .c ({signal_3507, signal_2052}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1785 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[71]), .c ({signal_3508, signal_2053}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1786 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[72]), .c ({signal_3509, signal_2054}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1787 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[73]), .c ({signal_3510, signal_2055}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1788 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[74]), .c ({signal_3511, signal_2056}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1789 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[75]), .c ({signal_3512, signal_2057}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1790 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[76]), .c ({signal_3513, signal_2058}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1791 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[77]), .c ({signal_3514, signal_2059}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1792 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[78]), .c ({signal_3515, signal_2060}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1793 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[79]), .c ({signal_3516, signal_2061}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1794 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[80]), .c ({signal_3517, signal_2062}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1795 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[81]), .c ({signal_3518, signal_2063}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1796 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[82]), .c ({signal_3519, signal_2064}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1797 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[83]), .c ({signal_3520, signal_2065}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1798 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[84]), .c ({signal_3521, signal_2066}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1799 ( .s ({signal_4702, signal_4700}), .b ({signal_4710, signal_4708}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[85]), .c ({signal_3522, signal_2067}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1800 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[86]), .c ({signal_3523, signal_2068}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1801 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[87]), .c ({signal_3524, signal_2069}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1802 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[88]), .c ({signal_3525, signal_2070}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1803 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[89]), .c ({signal_3526, signal_2071}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1804 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[90]), .c ({signal_3527, signal_2072}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1805 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[91]), .c ({signal_3528, signal_2073}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1806 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[92]), .c ({signal_3529, signal_2074}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1807 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[93]), .c ({signal_3530, signal_2075}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1808 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[94]), .c ({signal_3531, signal_2076}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1809 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[95]), .c ({signal_3532, signal_2077}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1810 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[96]), .c ({signal_3533, signal_2078}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1811 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[97]), .c ({signal_3534, signal_2079}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1812 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[98]), .c ({signal_3535, signal_2080}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1813 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[99]), .c ({signal_3536, signal_2081}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1814 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[100]), .c ({signal_3537, signal_2082}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1815 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[101]), .c ({signal_3538, signal_2083}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1816 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[102]), .c ({signal_3539, signal_2084}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1817 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[103]), .c ({signal_3540, signal_2085}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1818 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[104]), .c ({signal_3541, signal_2086}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1819 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[105]), .c ({signal_3542, signal_2087}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1820 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b0}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[106]), .c ({signal_3543, signal_2088}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1821 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[107]), .c ({signal_3544, signal_2089}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1822 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[108]), .c ({signal_3545, signal_2090}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1823 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[109]), .c ({signal_3546, signal_2091}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1824 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[110]), .c ({signal_3547, signal_2092}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1825 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[111]), .c ({signal_3548, signal_2093}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1826 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[112]), .c ({signal_3549, signal_2094}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1827 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[113]), .c ({signal_3550, signal_2095}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1828 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[114]), .c ({signal_3551, signal_2096}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1829 ( .s ({signal_4722, signal_4718}), .b ({signal_3443, signal_2012}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[115]), .c ({signal_3552, signal_2097}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1830 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[116]), .c ({signal_3553, signal_2098}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1831 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[117]), .c ({signal_3554, signal_2099}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1832 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[118]), .c ({signal_3555, signal_2100}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1833 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[119]), .c ({signal_3556, signal_2101}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1834 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b0}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[120]), .c ({signal_3557, signal_2102}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1835 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[121]), .c ({signal_3558, signal_2103}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1836 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[122]), .c ({signal_3559, signal_2104}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1837 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[123]), .c ({signal_3560, signal_2105}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1838 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[124]), .c ({signal_3561, signal_2106}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1839 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[125]), .c ({signal_3562, signal_2107}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1840 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[126]), .c ({signal_3563, signal_2108}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1841 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[127]), .c ({signal_3564, signal_2109}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1842 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[128]), .c ({signal_3565, signal_2110}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1843 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[129]), .c ({signal_3566, signal_2111}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1844 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[130]), .c ({signal_3567, signal_2112}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1845 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[131]), .c ({signal_3568, signal_2113}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1846 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[132]), .c ({signal_3569, signal_2114}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1847 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[133]), .c ({signal_3570, signal_2115}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1848 ( .s ({signal_4722, signal_4718}), .b ({signal_3446, signal_2015}), .a ({signal_3445, signal_2014}), .clk (clk), .r (Fresh[134]), .c ({signal_3571, signal_2116}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1849 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[135]), .c ({signal_3572, signal_2117}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1850 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[136]), .c ({signal_3573, signal_2118}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1851 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[137]), .c ({signal_3574, signal_2119}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1852 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[138]), .c ({signal_3575, signal_2120}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1853 ( .s ({signal_4702, signal_4700}), .b ({signal_4710, signal_4708}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[139]), .c ({signal_3576, signal_2121}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1854 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[140]), .c ({signal_3577, signal_2122}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1855 ( .s ({signal_4702, signal_4700}), .b ({signal_3434, signal_2003}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[141]), .c ({signal_3578, signal_2123}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1856 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[142]), .c ({signal_3579, signal_2124}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1857 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[143]), .c ({signal_3580, signal_2125}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1858 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[144]), .c ({signal_3581, signal_2126}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1859 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b0}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[145]), .c ({signal_3582, signal_2127}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1860 ( .s ({signal_4702, signal_4700}), .b ({signal_4710, signal_4708}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[146]), .c ({signal_3583, signal_2128}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1861 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b0}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[147]), .c ({signal_3584, signal_2129}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1862 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[148]), .c ({signal_3585, signal_2130}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1863 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[149]), .c ({signal_3586, signal_2131}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1864 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[150]), .c ({signal_3587, signal_2132}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1865 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[151]), .c ({signal_3588, signal_2133}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1866 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[152]), .c ({signal_3589, signal_2134}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1867 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[153]), .c ({signal_3590, signal_2135}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1868 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_3418, signal_1987}), .clk (clk), .r (Fresh[154]), .c ({signal_3591, signal_2136}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1869 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_4714, signal_4712}), .clk (clk), .r (Fresh[155]), .c ({signal_3592, signal_2137}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1870 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_4710, signal_4708}), .clk (clk), .r (Fresh[156]), .c ({signal_3593, signal_2138}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1871 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[157]), .c ({signal_3594, signal_2139}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1872 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[158]), .c ({signal_3595, signal_2140}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1873 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[159]), .c ({signal_3596, signal_2141}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1874 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[160]), .c ({signal_3597, signal_2142}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1875 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[161]), .c ({signal_3598, signal_2143}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1876 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[162]), .c ({signal_3599, signal_2144}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1877 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[163]), .c ({signal_3600, signal_2145}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1878 ( .s ({signal_4722, signal_4718}), .b ({signal_4730, signal_4728}), .a ({signal_3431, signal_2000}), .clk (clk), .r (Fresh[164]), .c ({signal_3601, signal_2146}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1879 ( .s ({signal_4722, signal_4718}), .b ({signal_3446, signal_2015}), .a ({signal_3450, signal_2019}), .clk (clk), .r (Fresh[165]), .c ({signal_3602, signal_2147}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1880 ( .s ({signal_4702, signal_4700}), .b ({signal_3428, signal_1997}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[166]), .c ({signal_3603, signal_2148}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1881 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_3419, signal_1988}), .clk (clk), .r (Fresh[167]), .c ({signal_3604, signal_2149}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1882 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[168]), .c ({signal_3605, signal_2150}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1883 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[169]), .c ({signal_3606, signal_2151}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1884 ( .s ({signal_4702, signal_4700}), .b ({signal_4714, signal_4712}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[170]), .c ({signal_3607, signal_2152}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1885 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b0}), .a ({signal_3421, signal_1990}), .clk (clk), .r (Fresh[171]), .c ({signal_3608, signal_2153}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1886 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[172]), .c ({signal_3609, signal_2154}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1887 ( .s ({signal_4702, signal_4700}), .b ({signal_3419, signal_1988}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[173]), .c ({signal_3610, signal_2155}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1888 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[174]), .c ({signal_3611, signal_2156}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1889 ( .s ({signal_4702, signal_4700}), .b ({signal_4706, signal_4704}), .a ({signal_3434, signal_2003}), .clk (clk), .r (Fresh[175]), .c ({signal_3612, signal_2157}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1890 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b1}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[176]), .c ({signal_3613, signal_2158}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1891 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[177]), .c ({signal_3614, signal_2159}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1892 ( .s ({signal_4702, signal_4700}), .b ({signal_3421, signal_1990}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[178]), .c ({signal_3615, signal_2160}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1893 ( .s ({signal_4702, signal_4700}), .b ({signal_3427, signal_1996}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[179]), .c ({signal_3616, signal_2161}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1894 ( .s ({signal_4702, signal_4700}), .b ({signal_3423, signal_1992}), .a ({signal_4706, signal_4704}), .clk (clk), .r (Fresh[180]), .c ({signal_3617, signal_2162}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1895 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3425, signal_1994}), .clk (clk), .r (Fresh[181]), .c ({signal_3618, signal_2163}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1896 ( .s ({signal_4702, signal_4700}), .b ({signal_4726, signal_4724}), .a ({signal_3428, signal_1997}), .clk (clk), .r (Fresh[182]), .c ({signal_3619, signal_2164}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1897 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[183]), .c ({signal_3620, signal_2165}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1898 ( .s ({signal_4702, signal_4700}), .b ({signal_3425, signal_1994}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[184]), .c ({signal_3621, signal_2166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1899 ( .s ({signal_4702, signal_4700}), .b ({signal_3422, signal_1991}), .a ({signal_3420, signal_1989}), .clk (clk), .r (Fresh[185]), .c ({signal_3622, signal_2167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1900 ( .s ({signal_4702, signal_4700}), .b ({1'b0, 1'b0}), .a ({signal_3423, signal_1992}), .clk (clk), .r (Fresh[186]), .c ({signal_3623, signal_2168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1901 ( .s ({signal_4702, signal_4700}), .b ({signal_3420, signal_1989}), .a ({signal_3427, signal_1996}), .clk (clk), .r (Fresh[187]), .c ({signal_3624, signal_2169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1902 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_4726, signal_4724}), .clk (clk), .r (Fresh[188]), .c ({signal_3625, signal_2170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1903 ( .s ({signal_4702, signal_4700}), .b ({signal_3418, signal_1987}), .a ({signal_3422, signal_1991}), .clk (clk), .r (Fresh[189]), .c ({signal_3626, signal_2171}) ) ;
    buf_clk cell_2186 ( .C (clk), .D (signal_4731), .Q (signal_4732) ) ;
    buf_clk cell_2188 ( .C (clk), .D (signal_4733), .Q (signal_4734) ) ;
    buf_clk cell_2190 ( .C (clk), .D (signal_4735), .Q (signal_4736) ) ;
    buf_clk cell_2192 ( .C (clk), .D (signal_4737), .Q (signal_4738) ) ;
    buf_clk cell_2194 ( .C (clk), .D (signal_4739), .Q (signal_4740) ) ;
    buf_clk cell_2196 ( .C (clk), .D (signal_4741), .Q (signal_4742) ) ;
    buf_clk cell_2198 ( .C (clk), .D (signal_4743), .Q (signal_4744) ) ;
    buf_clk cell_2200 ( .C (clk), .D (signal_4745), .Q (signal_4746) ) ;
    buf_clk cell_2202 ( .C (clk), .D (signal_4747), .Q (signal_4748) ) ;
    buf_clk cell_2204 ( .C (clk), .D (signal_4749), .Q (signal_4750) ) ;
    buf_clk cell_2206 ( .C (clk), .D (signal_4751), .Q (signal_4752) ) ;
    buf_clk cell_2208 ( .C (clk), .D (signal_4753), .Q (signal_4754) ) ;
    buf_clk cell_2210 ( .C (clk), .D (signal_4755), .Q (signal_4756) ) ;
    buf_clk cell_2212 ( .C (clk), .D (signal_4757), .Q (signal_4758) ) ;
    buf_clk cell_2214 ( .C (clk), .D (signal_4759), .Q (signal_4760) ) ;
    buf_clk cell_2216 ( .C (clk), .D (signal_4761), .Q (signal_4762) ) ;
    buf_clk cell_2218 ( .C (clk), .D (signal_4763), .Q (signal_4764) ) ;
    buf_clk cell_2220 ( .C (clk), .D (signal_4765), .Q (signal_4766) ) ;
    buf_clk cell_2222 ( .C (clk), .D (signal_4767), .Q (signal_4768) ) ;
    buf_clk cell_2224 ( .C (clk), .D (signal_4769), .Q (signal_4770) ) ;
    buf_clk cell_2226 ( .C (clk), .D (signal_4771), .Q (signal_4772) ) ;
    buf_clk cell_2228 ( .C (clk), .D (signal_4773), .Q (signal_4774) ) ;
    buf_clk cell_2230 ( .C (clk), .D (signal_4775), .Q (signal_4776) ) ;
    buf_clk cell_2232 ( .C (clk), .D (signal_4777), .Q (signal_4778) ) ;
    buf_clk cell_2234 ( .C (clk), .D (signal_4779), .Q (signal_4780) ) ;
    buf_clk cell_2236 ( .C (clk), .D (signal_4781), .Q (signal_4782) ) ;
    buf_clk cell_2238 ( .C (clk), .D (signal_4783), .Q (signal_4784) ) ;
    buf_clk cell_2240 ( .C (clk), .D (signal_4785), .Q (signal_4786) ) ;
    buf_clk cell_2242 ( .C (clk), .D (signal_4787), .Q (signal_4788) ) ;
    buf_clk cell_2244 ( .C (clk), .D (signal_4789), .Q (signal_4790) ) ;
    buf_clk cell_2246 ( .C (clk), .D (signal_4791), .Q (signal_4792) ) ;
    buf_clk cell_2248 ( .C (clk), .D (signal_4793), .Q (signal_4794) ) ;
    buf_clk cell_2250 ( .C (clk), .D (signal_4795), .Q (signal_4796) ) ;
    buf_clk cell_2252 ( .C (clk), .D (signal_4797), .Q (signal_4798) ) ;
    buf_clk cell_2254 ( .C (clk), .D (signal_4799), .Q (signal_4800) ) ;
    buf_clk cell_2256 ( .C (clk), .D (signal_4801), .Q (signal_4802) ) ;
    buf_clk cell_2258 ( .C (clk), .D (signal_4803), .Q (signal_4804) ) ;
    buf_clk cell_2260 ( .C (clk), .D (signal_4805), .Q (signal_4806) ) ;
    buf_clk cell_2262 ( .C (clk), .D (signal_4807), .Q (signal_4808) ) ;
    buf_clk cell_2264 ( .C (clk), .D (signal_4809), .Q (signal_4810) ) ;
    buf_clk cell_2266 ( .C (clk), .D (signal_4811), .Q (signal_4812) ) ;
    buf_clk cell_2268 ( .C (clk), .D (signal_4813), .Q (signal_4814) ) ;
    buf_clk cell_2270 ( .C (clk), .D (signal_4815), .Q (signal_4816) ) ;
    buf_clk cell_2272 ( .C (clk), .D (signal_4817), .Q (signal_4818) ) ;
    buf_clk cell_2274 ( .C (clk), .D (signal_4819), .Q (signal_4820) ) ;
    buf_clk cell_2276 ( .C (clk), .D (signal_4821), .Q (signal_4822) ) ;
    buf_clk cell_2278 ( .C (clk), .D (signal_4823), .Q (signal_4824) ) ;
    buf_clk cell_2280 ( .C (clk), .D (signal_4825), .Q (signal_4826) ) ;
    buf_clk cell_2282 ( .C (clk), .D (signal_4827), .Q (signal_4828) ) ;
    buf_clk cell_2284 ( .C (clk), .D (signal_4829), .Q (signal_4830) ) ;
    buf_clk cell_2286 ( .C (clk), .D (signal_4831), .Q (signal_4832) ) ;
    buf_clk cell_2288 ( .C (clk), .D (signal_4833), .Q (signal_4834) ) ;
    buf_clk cell_2290 ( .C (clk), .D (signal_4835), .Q (signal_4836) ) ;
    buf_clk cell_2292 ( .C (clk), .D (signal_4837), .Q (signal_4838) ) ;
    buf_clk cell_2294 ( .C (clk), .D (signal_4839), .Q (signal_4840) ) ;
    buf_clk cell_2296 ( .C (clk), .D (signal_4841), .Q (signal_4842) ) ;
    buf_clk cell_2302 ( .C (clk), .D (signal_4847), .Q (signal_4848) ) ;
    buf_clk cell_2310 ( .C (clk), .D (signal_4855), .Q (signal_4856) ) ;
    buf_clk cell_2346 ( .C (clk), .D (signal_4891), .Q (signal_4892) ) ;
    buf_clk cell_2356 ( .C (clk), .D (signal_4901), .Q (signal_4902) ) ;
    buf_clk cell_2366 ( .C (clk), .D (signal_4911), .Q (signal_4912) ) ;
    buf_clk cell_2378 ( .C (clk), .D (signal_4923), .Q (signal_4924) ) ;
    buf_clk cell_2390 ( .C (clk), .D (signal_4935), .Q (signal_4936) ) ;
    buf_clk cell_2406 ( .C (clk), .D (signal_4951), .Q (signal_4952) ) ;
    buf_clk cell_2422 ( .C (clk), .D (signal_4967), .Q (signal_4968) ) ;
    buf_clk cell_2438 ( .C (clk), .D (signal_4983), .Q (signal_4984) ) ;
    buf_clk cell_2454 ( .C (clk), .D (signal_4999), .Q (signal_5000) ) ;
    buf_clk cell_2470 ( .C (clk), .D (signal_5015), .Q (signal_5016) ) ;
    buf_clk cell_2486 ( .C (clk), .D (signal_5031), .Q (signal_5032) ) ;
    buf_clk cell_2502 ( .C (clk), .D (signal_5047), .Q (signal_5048) ) ;
    buf_clk cell_2518 ( .C (clk), .D (signal_5063), .Q (signal_5064) ) ;
    buf_clk cell_2534 ( .C (clk), .D (signal_5079), .Q (signal_5080) ) ;
    buf_clk cell_2550 ( .C (clk), .D (signal_5095), .Q (signal_5096) ) ;
    buf_clk cell_2566 ( .C (clk), .D (signal_5111), .Q (signal_5112) ) ;
    buf_clk cell_2582 ( .C (clk), .D (signal_5127), .Q (signal_5128) ) ;
    buf_clk cell_2598 ( .C (clk), .D (signal_5143), .Q (signal_5144) ) ;
    buf_clk cell_2614 ( .C (clk), .D (signal_5159), .Q (signal_5160) ) ;
    buf_clk cell_2630 ( .C (clk), .D (signal_5175), .Q (signal_5176) ) ;
    buf_clk cell_2646 ( .C (clk), .D (signal_5191), .Q (signal_5192) ) ;
    buf_clk cell_2662 ( .C (clk), .D (signal_5207), .Q (signal_5208) ) ;
    buf_clk cell_2678 ( .C (clk), .D (signal_5223), .Q (signal_5224) ) ;
    buf_clk cell_2694 ( .C (clk), .D (signal_5239), .Q (signal_5240) ) ;
    buf_clk cell_2710 ( .C (clk), .D (signal_5255), .Q (signal_5256) ) ;
    buf_clk cell_2726 ( .C (clk), .D (signal_5271), .Q (signal_5272) ) ;
    buf_clk cell_2742 ( .C (clk), .D (signal_5287), .Q (signal_5288) ) ;
    buf_clk cell_2758 ( .C (clk), .D (signal_5303), .Q (signal_5304) ) ;
    buf_clk cell_2774 ( .C (clk), .D (signal_5319), .Q (signal_5320) ) ;
    buf_clk cell_2790 ( .C (clk), .D (signal_5335), .Q (signal_5336) ) ;
    buf_clk cell_2806 ( .C (clk), .D (signal_5351), .Q (signal_5352) ) ;
    buf_clk cell_2822 ( .C (clk), .D (signal_5367), .Q (signal_5368) ) ;
    buf_clk cell_2838 ( .C (clk), .D (signal_5383), .Q (signal_5384) ) ;
    buf_clk cell_2854 ( .C (clk), .D (signal_5399), .Q (signal_5400) ) ;
    buf_clk cell_2870 ( .C (clk), .D (signal_5415), .Q (signal_5416) ) ;
    buf_clk cell_2886 ( .C (clk), .D (signal_5431), .Q (signal_5432) ) ;
    buf_clk cell_2902 ( .C (clk), .D (signal_5447), .Q (signal_5448) ) ;
    buf_clk cell_2918 ( .C (clk), .D (signal_5463), .Q (signal_5464) ) ;
    buf_clk cell_2934 ( .C (clk), .D (signal_5479), .Q (signal_5480) ) ;
    buf_clk cell_2950 ( .C (clk), .D (signal_5495), .Q (signal_5496) ) ;
    buf_clk cell_2966 ( .C (clk), .D (signal_5511), .Q (signal_5512) ) ;
    buf_clk cell_2982 ( .C (clk), .D (signal_5527), .Q (signal_5528) ) ;
    buf_clk cell_2998 ( .C (clk), .D (signal_5543), .Q (signal_5544) ) ;
    buf_clk cell_3014 ( .C (clk), .D (signal_5559), .Q (signal_5560) ) ;
    buf_clk cell_3030 ( .C (clk), .D (signal_5575), .Q (signal_5576) ) ;
    buf_clk cell_3046 ( .C (clk), .D (signal_5591), .Q (signal_5592) ) ;
    buf_clk cell_3062 ( .C (clk), .D (signal_5607), .Q (signal_5608) ) ;
    buf_clk cell_3078 ( .C (clk), .D (signal_5623), .Q (signal_5624) ) ;
    buf_clk cell_3094 ( .C (clk), .D (signal_5639), .Q (signal_5640) ) ;
    buf_clk cell_3110 ( .C (clk), .D (signal_5655), .Q (signal_5656) ) ;
    buf_clk cell_3126 ( .C (clk), .D (signal_5671), .Q (signal_5672) ) ;
    buf_clk cell_3142 ( .C (clk), .D (signal_5687), .Q (signal_5688) ) ;
    buf_clk cell_3158 ( .C (clk), .D (signal_5703), .Q (signal_5704) ) ;
    buf_clk cell_3174 ( .C (clk), .D (signal_5719), .Q (signal_5720) ) ;
    buf_clk cell_3190 ( .C (clk), .D (signal_5735), .Q (signal_5736) ) ;
    buf_clk cell_3206 ( .C (clk), .D (signal_5751), .Q (signal_5752) ) ;
    buf_clk cell_3222 ( .C (clk), .D (signal_5767), .Q (signal_5768) ) ;
    buf_clk cell_3238 ( .C (clk), .D (signal_5783), .Q (signal_5784) ) ;
    buf_clk cell_3254 ( .C (clk), .D (signal_5799), .Q (signal_5800) ) ;
    buf_clk cell_3270 ( .C (clk), .D (signal_5815), .Q (signal_5816) ) ;
    buf_clk cell_3286 ( .C (clk), .D (signal_5831), .Q (signal_5832) ) ;
    buf_clk cell_3302 ( .C (clk), .D (signal_5847), .Q (signal_5848) ) ;
    buf_clk cell_3318 ( .C (clk), .D (signal_5863), .Q (signal_5864) ) ;
    buf_clk cell_3334 ( .C (clk), .D (signal_5879), .Q (signal_5880) ) ;
    buf_clk cell_3350 ( .C (clk), .D (signal_5895), .Q (signal_5896) ) ;
    buf_clk cell_3366 ( .C (clk), .D (signal_5911), .Q (signal_5912) ) ;
    buf_clk cell_3382 ( .C (clk), .D (signal_5927), .Q (signal_5928) ) ;
    buf_clk cell_3398 ( .C (clk), .D (signal_5943), .Q (signal_5944) ) ;
    buf_clk cell_3414 ( .C (clk), .D (signal_5959), .Q (signal_5960) ) ;
    buf_clk cell_3430 ( .C (clk), .D (signal_5975), .Q (signal_5976) ) ;
    buf_clk cell_3446 ( .C (clk), .D (signal_5991), .Q (signal_5992) ) ;
    buf_clk cell_3462 ( .C (clk), .D (signal_6007), .Q (signal_6008) ) ;
    buf_clk cell_3478 ( .C (clk), .D (signal_6023), .Q (signal_6024) ) ;
    buf_clk cell_3494 ( .C (clk), .D (signal_6039), .Q (signal_6040) ) ;
    buf_clk cell_3510 ( .C (clk), .D (signal_6055), .Q (signal_6056) ) ;
    buf_clk cell_3526 ( .C (clk), .D (signal_6071), .Q (signal_6072) ) ;
    buf_clk cell_3542 ( .C (clk), .D (signal_6087), .Q (signal_6088) ) ;
    buf_clk cell_3558 ( .C (clk), .D (signal_6103), .Q (signal_6104) ) ;
    buf_clk cell_3574 ( .C (clk), .D (signal_6119), .Q (signal_6120) ) ;
    buf_clk cell_3590 ( .C (clk), .D (signal_6135), .Q (signal_6136) ) ;
    buf_clk cell_3606 ( .C (clk), .D (signal_6151), .Q (signal_6152) ) ;
    buf_clk cell_3622 ( .C (clk), .D (signal_6167), .Q (signal_6168) ) ;
    buf_clk cell_3638 ( .C (clk), .D (signal_6183), .Q (signal_6184) ) ;
    buf_clk cell_3654 ( .C (clk), .D (signal_6199), .Q (signal_6200) ) ;
    buf_clk cell_3670 ( .C (clk), .D (signal_6215), .Q (signal_6216) ) ;
    buf_clk cell_3686 ( .C (clk), .D (signal_6231), .Q (signal_6232) ) ;
    buf_clk cell_3702 ( .C (clk), .D (signal_6247), .Q (signal_6248) ) ;
    buf_clk cell_3718 ( .C (clk), .D (signal_6263), .Q (signal_6264) ) ;
    buf_clk cell_3734 ( .C (clk), .D (signal_6279), .Q (signal_6280) ) ;
    buf_clk cell_3750 ( .C (clk), .D (signal_6295), .Q (signal_6296) ) ;
    buf_clk cell_3766 ( .C (clk), .D (signal_6311), .Q (signal_6312) ) ;
    buf_clk cell_3782 ( .C (clk), .D (signal_6327), .Q (signal_6328) ) ;
    buf_clk cell_3798 ( .C (clk), .D (signal_6343), .Q (signal_6344) ) ;
    buf_clk cell_3814 ( .C (clk), .D (signal_6359), .Q (signal_6360) ) ;
    buf_clk cell_3830 ( .C (clk), .D (signal_6375), .Q (signal_6376) ) ;
    buf_clk cell_3846 ( .C (clk), .D (signal_6391), .Q (signal_6392) ) ;
    buf_clk cell_3862 ( .C (clk), .D (signal_6407), .Q (signal_6408) ) ;
    buf_clk cell_3878 ( .C (clk), .D (signal_6423), .Q (signal_6424) ) ;
    buf_clk cell_3894 ( .C (clk), .D (signal_6439), .Q (signal_6440) ) ;
    buf_clk cell_3910 ( .C (clk), .D (signal_6455), .Q (signal_6456) ) ;
    buf_clk cell_3926 ( .C (clk), .D (signal_6471), .Q (signal_6472) ) ;
    buf_clk cell_3942 ( .C (clk), .D (signal_6487), .Q (signal_6488) ) ;
    buf_clk cell_3958 ( .C (clk), .D (signal_6503), .Q (signal_6504) ) ;
    buf_clk cell_3974 ( .C (clk), .D (signal_6519), .Q (signal_6520) ) ;
    buf_clk cell_3990 ( .C (clk), .D (signal_6535), .Q (signal_6536) ) ;
    buf_clk cell_4006 ( .C (clk), .D (signal_6551), .Q (signal_6552) ) ;
    buf_clk cell_4022 ( .C (clk), .D (signal_6567), .Q (signal_6568) ) ;
    buf_clk cell_4038 ( .C (clk), .D (signal_6583), .Q (signal_6584) ) ;
    buf_clk cell_4054 ( .C (clk), .D (signal_6599), .Q (signal_6600) ) ;
    buf_clk cell_4070 ( .C (clk), .D (signal_6615), .Q (signal_6616) ) ;
    buf_clk cell_4086 ( .C (clk), .D (signal_6631), .Q (signal_6632) ) ;
    buf_clk cell_4102 ( .C (clk), .D (signal_6647), .Q (signal_6648) ) ;
    buf_clk cell_4118 ( .C (clk), .D (signal_6663), .Q (signal_6664) ) ;
    buf_clk cell_4134 ( .C (clk), .D (signal_6679), .Q (signal_6680) ) ;
    buf_clk cell_4150 ( .C (clk), .D (signal_6695), .Q (signal_6696) ) ;
    buf_clk cell_4166 ( .C (clk), .D (signal_6711), .Q (signal_6712) ) ;
    buf_clk cell_4182 ( .C (clk), .D (signal_6727), .Q (signal_6728) ) ;
    buf_clk cell_4198 ( .C (clk), .D (signal_6743), .Q (signal_6744) ) ;
    buf_clk cell_4214 ( .C (clk), .D (signal_6759), .Q (signal_6760) ) ;
    buf_clk cell_4230 ( .C (clk), .D (signal_6775), .Q (signal_6776) ) ;
    buf_clk cell_4246 ( .C (clk), .D (signal_6791), .Q (signal_6792) ) ;
    buf_clk cell_4262 ( .C (clk), .D (signal_6807), .Q (signal_6808) ) ;
    buf_clk cell_4278 ( .C (clk), .D (signal_6823), .Q (signal_6824) ) ;
    buf_clk cell_4294 ( .C (clk), .D (signal_6839), .Q (signal_6840) ) ;
    buf_clk cell_4310 ( .C (clk), .D (signal_6855), .Q (signal_6856) ) ;
    buf_clk cell_4326 ( .C (clk), .D (signal_6871), .Q (signal_6872) ) ;
    buf_clk cell_4342 ( .C (clk), .D (signal_6887), .Q (signal_6888) ) ;
    buf_clk cell_4358 ( .C (clk), .D (signal_6903), .Q (signal_6904) ) ;
    buf_clk cell_4374 ( .C (clk), .D (signal_6919), .Q (signal_6920) ) ;
    buf_clk cell_4390 ( .C (clk), .D (signal_6935), .Q (signal_6936) ) ;
    buf_clk cell_4406 ( .C (clk), .D (signal_6951), .Q (signal_6952) ) ;
    buf_clk cell_4420 ( .C (clk), .D (signal_6965), .Q (signal_6966) ) ;
    buf_clk cell_4434 ( .C (clk), .D (signal_6979), .Q (signal_6980) ) ;
    buf_clk cell_4450 ( .C (clk), .D (signal_6995), .Q (signal_6996) ) ;
    buf_clk cell_4466 ( .C (clk), .D (signal_7011), .Q (signal_7012) ) ;
    buf_clk cell_4482 ( .C (clk), .D (signal_7027), .Q (signal_7028) ) ;
    buf_clk cell_4498 ( .C (clk), .D (signal_7043), .Q (signal_7044) ) ;
    buf_clk cell_4514 ( .C (clk), .D (signal_7059), .Q (signal_7060) ) ;
    buf_clk cell_4530 ( .C (clk), .D (signal_7075), .Q (signal_7076) ) ;
    buf_clk cell_4546 ( .C (clk), .D (signal_7091), .Q (signal_7092) ) ;
    buf_clk cell_4562 ( .C (clk), .D (signal_7107), .Q (signal_7108) ) ;
    buf_clk cell_4578 ( .C (clk), .D (signal_7123), .Q (signal_7124) ) ;
    buf_clk cell_4594 ( .C (clk), .D (signal_7139), .Q (signal_7140) ) ;
    buf_clk cell_4610 ( .C (clk), .D (signal_7155), .Q (signal_7156) ) ;
    buf_clk cell_4626 ( .C (clk), .D (signal_7171), .Q (signal_7172) ) ;
    buf_clk cell_4642 ( .C (clk), .D (signal_7187), .Q (signal_7188) ) ;
    buf_clk cell_4658 ( .C (clk), .D (signal_7203), .Q (signal_7204) ) ;
    buf_clk cell_4674 ( .C (clk), .D (signal_7219), .Q (signal_7220) ) ;
    buf_clk cell_4690 ( .C (clk), .D (signal_7235), .Q (signal_7236) ) ;
    buf_clk cell_4706 ( .C (clk), .D (signal_7251), .Q (signal_7252) ) ;
    buf_clk cell_4722 ( .C (clk), .D (signal_7267), .Q (signal_7268) ) ;
    buf_clk cell_4738 ( .C (clk), .D (signal_7283), .Q (signal_7284) ) ;
    buf_clk cell_4754 ( .C (clk), .D (signal_7299), .Q (signal_7300) ) ;
    buf_clk cell_4770 ( .C (clk), .D (signal_7315), .Q (signal_7316) ) ;
    buf_clk cell_4786 ( .C (clk), .D (signal_7331), .Q (signal_7332) ) ;
    buf_clk cell_4802 ( .C (clk), .D (signal_7347), .Q (signal_7348) ) ;
    buf_clk cell_4818 ( .C (clk), .D (signal_7363), .Q (signal_7364) ) ;
    buf_clk cell_4834 ( .C (clk), .D (signal_7379), .Q (signal_7380) ) ;
    buf_clk cell_4850 ( .C (clk), .D (signal_7395), .Q (signal_7396) ) ;
    buf_clk cell_4866 ( .C (clk), .D (signal_7411), .Q (signal_7412) ) ;
    buf_clk cell_4882 ( .C (clk), .D (signal_7427), .Q (signal_7428) ) ;
    buf_clk cell_4898 ( .C (clk), .D (signal_7443), .Q (signal_7444) ) ;
    buf_clk cell_4914 ( .C (clk), .D (signal_7459), .Q (signal_7460) ) ;
    buf_clk cell_4930 ( .C (clk), .D (signal_7475), .Q (signal_7476) ) ;
    buf_clk cell_4946 ( .C (clk), .D (signal_7491), .Q (signal_7492) ) ;
    buf_clk cell_4962 ( .C (clk), .D (signal_7507), .Q (signal_7508) ) ;
    buf_clk cell_4978 ( .C (clk), .D (signal_7523), .Q (signal_7524) ) ;
    buf_clk cell_4994 ( .C (clk), .D (signal_7539), .Q (signal_7540) ) ;
    buf_clk cell_5010 ( .C (clk), .D (signal_7555), .Q (signal_7556) ) ;
    buf_clk cell_5026 ( .C (clk), .D (signal_7571), .Q (signal_7572) ) ;
    buf_clk cell_5042 ( .C (clk), .D (signal_7587), .Q (signal_7588) ) ;
    buf_clk cell_5058 ( .C (clk), .D (signal_7603), .Q (signal_7604) ) ;
    buf_clk cell_5074 ( .C (clk), .D (signal_7619), .Q (signal_7620) ) ;
    buf_clk cell_5090 ( .C (clk), .D (signal_7635), .Q (signal_7636) ) ;
    buf_clk cell_5106 ( .C (clk), .D (signal_7651), .Q (signal_7652) ) ;
    buf_clk cell_5122 ( .C (clk), .D (signal_7667), .Q (signal_7668) ) ;
    buf_clk cell_5138 ( .C (clk), .D (signal_7683), .Q (signal_7684) ) ;
    buf_clk cell_5154 ( .C (clk), .D (signal_7699), .Q (signal_7700) ) ;
    buf_clk cell_5170 ( .C (clk), .D (signal_7715), .Q (signal_7716) ) ;
    buf_clk cell_5186 ( .C (clk), .D (signal_7731), .Q (signal_7732) ) ;
    buf_clk cell_5202 ( .C (clk), .D (signal_7747), .Q (signal_7748) ) ;
    buf_clk cell_5218 ( .C (clk), .D (signal_7763), .Q (signal_7764) ) ;
    buf_clk cell_5234 ( .C (clk), .D (signal_7779), .Q (signal_7780) ) ;
    buf_clk cell_5250 ( .C (clk), .D (signal_7795), .Q (signal_7796) ) ;
    buf_clk cell_5266 ( .C (clk), .D (signal_7811), .Q (signal_7812) ) ;
    buf_clk cell_5282 ( .C (clk), .D (signal_7827), .Q (signal_7828) ) ;
    buf_clk cell_5298 ( .C (clk), .D (signal_7843), .Q (signal_7844) ) ;
    buf_clk cell_5314 ( .C (clk), .D (signal_7859), .Q (signal_7860) ) ;
    buf_clk cell_5330 ( .C (clk), .D (signal_7875), .Q (signal_7876) ) ;
    buf_clk cell_5346 ( .C (clk), .D (signal_7891), .Q (signal_7892) ) ;
    buf_clk cell_5362 ( .C (clk), .D (signal_7907), .Q (signal_7908) ) ;
    buf_clk cell_5378 ( .C (clk), .D (signal_7923), .Q (signal_7924) ) ;
    buf_clk cell_5394 ( .C (clk), .D (signal_7939), .Q (signal_7940) ) ;
    buf_clk cell_5410 ( .C (clk), .D (signal_7955), .Q (signal_7956) ) ;
    buf_clk cell_5426 ( .C (clk), .D (signal_7971), .Q (signal_7972) ) ;
    buf_clk cell_5442 ( .C (clk), .D (signal_7987), .Q (signal_7988) ) ;
    buf_clk cell_5458 ( .C (clk), .D (signal_8003), .Q (signal_8004) ) ;
    buf_clk cell_5474 ( .C (clk), .D (signal_8019), .Q (signal_8020) ) ;
    buf_clk cell_5490 ( .C (clk), .D (signal_8035), .Q (signal_8036) ) ;
    buf_clk cell_5506 ( .C (clk), .D (signal_8051), .Q (signal_8052) ) ;
    buf_clk cell_5522 ( .C (clk), .D (signal_8067), .Q (signal_8068) ) ;
    buf_clk cell_5538 ( .C (clk), .D (signal_8083), .Q (signal_8084) ) ;
    buf_clk cell_5554 ( .C (clk), .D (signal_8099), .Q (signal_8100) ) ;
    buf_clk cell_5570 ( .C (clk), .D (signal_8115), .Q (signal_8116) ) ;
    buf_clk cell_5586 ( .C (clk), .D (signal_8131), .Q (signal_8132) ) ;
    buf_clk cell_5602 ( .C (clk), .D (signal_8147), .Q (signal_8148) ) ;
    buf_clk cell_5618 ( .C (clk), .D (signal_8163), .Q (signal_8164) ) ;
    buf_clk cell_5634 ( .C (clk), .D (signal_8179), .Q (signal_8180) ) ;
    buf_clk cell_5650 ( .C (clk), .D (signal_8195), .Q (signal_8196) ) ;
    buf_clk cell_5666 ( .C (clk), .D (signal_8211), .Q (signal_8212) ) ;
    buf_clk cell_5682 ( .C (clk), .D (signal_8227), .Q (signal_8228) ) ;
    buf_clk cell_5698 ( .C (clk), .D (signal_8243), .Q (signal_8244) ) ;
    buf_clk cell_5714 ( .C (clk), .D (signal_8259), .Q (signal_8260) ) ;
    buf_clk cell_5730 ( .C (clk), .D (signal_8275), .Q (signal_8276) ) ;
    buf_clk cell_5746 ( .C (clk), .D (signal_8291), .Q (signal_8292) ) ;
    buf_clk cell_5762 ( .C (clk), .D (signal_8307), .Q (signal_8308) ) ;
    buf_clk cell_5778 ( .C (clk), .D (signal_8323), .Q (signal_8324) ) ;
    buf_clk cell_5794 ( .C (clk), .D (signal_8339), .Q (signal_8340) ) ;
    buf_clk cell_5810 ( .C (clk), .D (signal_8355), .Q (signal_8356) ) ;
    buf_clk cell_5826 ( .C (clk), .D (signal_8371), .Q (signal_8372) ) ;
    buf_clk cell_5842 ( .C (clk), .D (signal_8387), .Q (signal_8388) ) ;
    buf_clk cell_5858 ( .C (clk), .D (signal_8403), .Q (signal_8404) ) ;
    buf_clk cell_5874 ( .C (clk), .D (signal_8419), .Q (signal_8420) ) ;
    buf_clk cell_5890 ( .C (clk), .D (signal_8435), .Q (signal_8436) ) ;
    buf_clk cell_5906 ( .C (clk), .D (signal_8451), .Q (signal_8452) ) ;
    buf_clk cell_5922 ( .C (clk), .D (signal_8467), .Q (signal_8468) ) ;
    buf_clk cell_5938 ( .C (clk), .D (signal_8483), .Q (signal_8484) ) ;
    buf_clk cell_5954 ( .C (clk), .D (signal_8499), .Q (signal_8500) ) ;
    buf_clk cell_5970 ( .C (clk), .D (signal_8515), .Q (signal_8516) ) ;
    buf_clk cell_5986 ( .C (clk), .D (signal_8531), .Q (signal_8532) ) ;
    buf_clk cell_6002 ( .C (clk), .D (signal_8547), .Q (signal_8548) ) ;
    buf_clk cell_6018 ( .C (clk), .D (signal_8563), .Q (signal_8564) ) ;
    buf_clk cell_6034 ( .C (clk), .D (signal_8579), .Q (signal_8580) ) ;
    buf_clk cell_6050 ( .C (clk), .D (signal_8595), .Q (signal_8596) ) ;
    buf_clk cell_6066 ( .C (clk), .D (signal_8611), .Q (signal_8612) ) ;
    buf_clk cell_6082 ( .C (clk), .D (signal_8627), .Q (signal_8628) ) ;
    buf_clk cell_6098 ( .C (clk), .D (signal_8643), .Q (signal_8644) ) ;
    buf_clk cell_6114 ( .C (clk), .D (signal_8659), .Q (signal_8660) ) ;
    buf_clk cell_6130 ( .C (clk), .D (signal_8675), .Q (signal_8676) ) ;
    buf_clk cell_6146 ( .C (clk), .D (signal_8691), .Q (signal_8692) ) ;
    buf_clk cell_6162 ( .C (clk), .D (signal_8707), .Q (signal_8708) ) ;
    buf_clk cell_6178 ( .C (clk), .D (signal_8723), .Q (signal_8724) ) ;
    buf_clk cell_6194 ( .C (clk), .D (signal_8739), .Q (signal_8740) ) ;
    buf_clk cell_6210 ( .C (clk), .D (signal_8755), .Q (signal_8756) ) ;
    buf_clk cell_6226 ( .C (clk), .D (signal_8771), .Q (signal_8772) ) ;
    buf_clk cell_6242 ( .C (clk), .D (signal_8787), .Q (signal_8788) ) ;
    buf_clk cell_6258 ( .C (clk), .D (signal_8803), .Q (signal_8804) ) ;
    buf_clk cell_6274 ( .C (clk), .D (signal_8819), .Q (signal_8820) ) ;
    buf_clk cell_6290 ( .C (clk), .D (signal_8835), .Q (signal_8836) ) ;
    buf_clk cell_6306 ( .C (clk), .D (signal_8851), .Q (signal_8852) ) ;
    buf_clk cell_6322 ( .C (clk), .D (signal_8867), .Q (signal_8868) ) ;
    buf_clk cell_6338 ( .C (clk), .D (signal_8883), .Q (signal_8884) ) ;
    buf_clk cell_6354 ( .C (clk), .D (signal_8899), .Q (signal_8900) ) ;
    buf_clk cell_6370 ( .C (clk), .D (signal_8915), .Q (signal_8916) ) ;
    buf_clk cell_6386 ( .C (clk), .D (signal_8931), .Q (signal_8932) ) ;
    buf_clk cell_6402 ( .C (clk), .D (signal_8947), .Q (signal_8948) ) ;
    buf_clk cell_6418 ( .C (clk), .D (signal_8963), .Q (signal_8964) ) ;
    buf_clk cell_6434 ( .C (clk), .D (signal_8979), .Q (signal_8980) ) ;
    buf_clk cell_6450 ( .C (clk), .D (signal_8995), .Q (signal_8996) ) ;
    buf_clk cell_6466 ( .C (clk), .D (signal_9011), .Q (signal_9012) ) ;
    buf_clk cell_6482 ( .C (clk), .D (signal_9027), .Q (signal_9028) ) ;
    buf_clk cell_6498 ( .C (clk), .D (signal_9043), .Q (signal_9044) ) ;
    buf_clk cell_6514 ( .C (clk), .D (signal_9059), .Q (signal_9060) ) ;
    buf_clk cell_6530 ( .C (clk), .D (signal_9075), .Q (signal_9076) ) ;
    buf_clk cell_6546 ( .C (clk), .D (signal_9091), .Q (signal_9092) ) ;
    buf_clk cell_6562 ( .C (clk), .D (signal_9107), .Q (signal_9108) ) ;
    buf_clk cell_6578 ( .C (clk), .D (signal_9123), .Q (signal_9124) ) ;
    buf_clk cell_6594 ( .C (clk), .D (signal_9139), .Q (signal_9140) ) ;
    buf_clk cell_6610 ( .C (clk), .D (signal_9155), .Q (signal_9156) ) ;
    buf_clk cell_6626 ( .C (clk), .D (signal_9171), .Q (signal_9172) ) ;
    buf_clk cell_6642 ( .C (clk), .D (signal_9187), .Q (signal_9188) ) ;
    buf_clk cell_6658 ( .C (clk), .D (signal_9203), .Q (signal_9204) ) ;
    buf_clk cell_6674 ( .C (clk), .D (signal_9219), .Q (signal_9220) ) ;
    buf_clk cell_6690 ( .C (clk), .D (signal_9235), .Q (signal_9236) ) ;
    buf_clk cell_6706 ( .C (clk), .D (signal_9251), .Q (signal_9252) ) ;
    buf_clk cell_6722 ( .C (clk), .D (signal_9267), .Q (signal_9268) ) ;
    buf_clk cell_6738 ( .C (clk), .D (signal_9283), .Q (signal_9284) ) ;
    buf_clk cell_6754 ( .C (clk), .D (signal_9299), .Q (signal_9300) ) ;
    buf_clk cell_6770 ( .C (clk), .D (signal_9315), .Q (signal_9316) ) ;
    buf_clk cell_6786 ( .C (clk), .D (signal_9331), .Q (signal_9332) ) ;
    buf_clk cell_6802 ( .C (clk), .D (signal_9347), .Q (signal_9348) ) ;
    buf_clk cell_6818 ( .C (clk), .D (signal_9363), .Q (signal_9364) ) ;
    buf_clk cell_6834 ( .C (clk), .D (signal_9379), .Q (signal_9380) ) ;
    buf_clk cell_6850 ( .C (clk), .D (signal_9395), .Q (signal_9396) ) ;
    buf_clk cell_6866 ( .C (clk), .D (signal_9411), .Q (signal_9412) ) ;
    buf_clk cell_6882 ( .C (clk), .D (signal_9427), .Q (signal_9428) ) ;
    buf_clk cell_6898 ( .C (clk), .D (signal_9443), .Q (signal_9444) ) ;
    buf_clk cell_6914 ( .C (clk), .D (signal_9459), .Q (signal_9460) ) ;
    buf_clk cell_6930 ( .C (clk), .D (signal_9475), .Q (signal_9476) ) ;
    buf_clk cell_6946 ( .C (clk), .D (signal_9491), .Q (signal_9492) ) ;
    buf_clk cell_6962 ( .C (clk), .D (signal_9507), .Q (signal_9508) ) ;
    buf_clk cell_6978 ( .C (clk), .D (signal_9523), .Q (signal_9524) ) ;
    buf_clk cell_6994 ( .C (clk), .D (signal_9539), .Q (signal_9540) ) ;
    buf_clk cell_7010 ( .C (clk), .D (signal_9555), .Q (signal_9556) ) ;
    buf_clk cell_7026 ( .C (clk), .D (signal_9571), .Q (signal_9572) ) ;
    buf_clk cell_7042 ( .C (clk), .D (signal_9587), .Q (signal_9588) ) ;
    buf_clk cell_7058 ( .C (clk), .D (signal_9603), .Q (signal_9604) ) ;
    buf_clk cell_7074 ( .C (clk), .D (signal_9619), .Q (signal_9620) ) ;
    buf_clk cell_7090 ( .C (clk), .D (signal_9635), .Q (signal_9636) ) ;
    buf_clk cell_7106 ( .C (clk), .D (signal_9651), .Q (signal_9652) ) ;
    buf_clk cell_7122 ( .C (clk), .D (signal_9667), .Q (signal_9668) ) ;
    buf_clk cell_7138 ( .C (clk), .D (signal_9683), .Q (signal_9684) ) ;
    buf_clk cell_7154 ( .C (clk), .D (signal_9699), .Q (signal_9700) ) ;
    buf_clk cell_7170 ( .C (clk), .D (signal_9715), .Q (signal_9716) ) ;
    buf_clk cell_7186 ( .C (clk), .D (signal_9731), .Q (signal_9732) ) ;
    buf_clk cell_7202 ( .C (clk), .D (signal_9747), .Q (signal_9748) ) ;
    buf_clk cell_7218 ( .C (clk), .D (signal_9763), .Q (signal_9764) ) ;
    buf_clk cell_7234 ( .C (clk), .D (signal_9779), .Q (signal_9780) ) ;
    buf_clk cell_7250 ( .C (clk), .D (signal_9795), .Q (signal_9796) ) ;
    buf_clk cell_7266 ( .C (clk), .D (signal_9811), .Q (signal_9812) ) ;
    buf_clk cell_7282 ( .C (clk), .D (signal_9827), .Q (signal_9828) ) ;
    buf_clk cell_7298 ( .C (clk), .D (signal_9843), .Q (signal_9844) ) ;
    buf_clk cell_7314 ( .C (clk), .D (signal_9859), .Q (signal_9860) ) ;
    buf_clk cell_7330 ( .C (clk), .D (signal_9875), .Q (signal_9876) ) ;
    buf_clk cell_7346 ( .C (clk), .D (signal_9891), .Q (signal_9892) ) ;
    buf_clk cell_7362 ( .C (clk), .D (signal_9907), .Q (signal_9908) ) ;
    buf_clk cell_7378 ( .C (clk), .D (signal_9923), .Q (signal_9924) ) ;
    buf_clk cell_7394 ( .C (clk), .D (signal_9939), .Q (signal_9940) ) ;
    buf_clk cell_7410 ( .C (clk), .D (signal_9955), .Q (signal_9956) ) ;
    buf_clk cell_7426 ( .C (clk), .D (signal_9971), .Q (signal_9972) ) ;
    buf_clk cell_7442 ( .C (clk), .D (signal_9987), .Q (signal_9988) ) ;
    buf_clk cell_7458 ( .C (clk), .D (signal_10003), .Q (signal_10004) ) ;
    buf_clk cell_7474 ( .C (clk), .D (signal_10019), .Q (signal_10020) ) ;
    buf_clk cell_7490 ( .C (clk), .D (signal_10035), .Q (signal_10036) ) ;
    buf_clk cell_7506 ( .C (clk), .D (signal_10051), .Q (signal_10052) ) ;
    buf_clk cell_7522 ( .C (clk), .D (signal_10067), .Q (signal_10068) ) ;
    buf_clk cell_7538 ( .C (clk), .D (signal_10083), .Q (signal_10084) ) ;
    buf_clk cell_7554 ( .C (clk), .D (signal_10099), .Q (signal_10100) ) ;
    buf_clk cell_7570 ( .C (clk), .D (signal_10115), .Q (signal_10116) ) ;
    buf_clk cell_7586 ( .C (clk), .D (signal_10131), .Q (signal_10132) ) ;
    buf_clk cell_7602 ( .C (clk), .D (signal_10147), .Q (signal_10148) ) ;
    buf_clk cell_7618 ( .C (clk), .D (signal_10163), .Q (signal_10164) ) ;
    buf_clk cell_7634 ( .C (clk), .D (signal_10179), .Q (signal_10180) ) ;
    buf_clk cell_7650 ( .C (clk), .D (signal_10195), .Q (signal_10196) ) ;
    buf_clk cell_7666 ( .C (clk), .D (signal_10211), .Q (signal_10212) ) ;
    buf_clk cell_7682 ( .C (clk), .D (signal_10227), .Q (signal_10228) ) ;
    buf_clk cell_7698 ( .C (clk), .D (signal_10243), .Q (signal_10244) ) ;
    buf_clk cell_7714 ( .C (clk), .D (signal_10259), .Q (signal_10260) ) ;
    buf_clk cell_7730 ( .C (clk), .D (signal_10275), .Q (signal_10276) ) ;
    buf_clk cell_7746 ( .C (clk), .D (signal_10291), .Q (signal_10292) ) ;
    buf_clk cell_7762 ( .C (clk), .D (signal_10307), .Q (signal_10308) ) ;
    buf_clk cell_7778 ( .C (clk), .D (signal_10323), .Q (signal_10324) ) ;
    buf_clk cell_7794 ( .C (clk), .D (signal_10339), .Q (signal_10340) ) ;
    buf_clk cell_7810 ( .C (clk), .D (signal_10355), .Q (signal_10356) ) ;
    buf_clk cell_7826 ( .C (clk), .D (signal_10371), .Q (signal_10372) ) ;
    buf_clk cell_7842 ( .C (clk), .D (signal_10387), .Q (signal_10388) ) ;
    buf_clk cell_7858 ( .C (clk), .D (signal_10403), .Q (signal_10404) ) ;
    buf_clk cell_7874 ( .C (clk), .D (signal_10419), .Q (signal_10420) ) ;
    buf_clk cell_7890 ( .C (clk), .D (signal_10435), .Q (signal_10436) ) ;
    buf_clk cell_7906 ( .C (clk), .D (signal_10451), .Q (signal_10452) ) ;
    buf_clk cell_7922 ( .C (clk), .D (signal_10467), .Q (signal_10468) ) ;
    buf_clk cell_7938 ( .C (clk), .D (signal_10483), .Q (signal_10484) ) ;
    buf_clk cell_7954 ( .C (clk), .D (signal_10499), .Q (signal_10500) ) ;
    buf_clk cell_7970 ( .C (clk), .D (signal_10515), .Q (signal_10516) ) ;
    buf_clk cell_7986 ( .C (clk), .D (signal_10531), .Q (signal_10532) ) ;
    buf_clk cell_8002 ( .C (clk), .D (signal_10547), .Q (signal_10548) ) ;
    buf_clk cell_8018 ( .C (clk), .D (signal_10563), .Q (signal_10564) ) ;
    buf_clk cell_8034 ( .C (clk), .D (signal_10579), .Q (signal_10580) ) ;
    buf_clk cell_8050 ( .C (clk), .D (signal_10595), .Q (signal_10596) ) ;
    buf_clk cell_8066 ( .C (clk), .D (signal_10611), .Q (signal_10612) ) ;
    buf_clk cell_8082 ( .C (clk), .D (signal_10627), .Q (signal_10628) ) ;
    buf_clk cell_8098 ( .C (clk), .D (signal_10643), .Q (signal_10644) ) ;
    buf_clk cell_8114 ( .C (clk), .D (signal_10659), .Q (signal_10660) ) ;
    buf_clk cell_8130 ( .C (clk), .D (signal_10675), .Q (signal_10676) ) ;
    buf_clk cell_8146 ( .C (clk), .D (signal_10691), .Q (signal_10692) ) ;
    buf_clk cell_8162 ( .C (clk), .D (signal_10707), .Q (signal_10708) ) ;
    buf_clk cell_8178 ( .C (clk), .D (signal_10723), .Q (signal_10724) ) ;
    buf_clk cell_8194 ( .C (clk), .D (signal_10739), .Q (signal_10740) ) ;
    buf_clk cell_8210 ( .C (clk), .D (signal_10755), .Q (signal_10756) ) ;
    buf_clk cell_8226 ( .C (clk), .D (signal_10771), .Q (signal_10772) ) ;
    buf_clk cell_8242 ( .C (clk), .D (signal_10787), .Q (signal_10788) ) ;
    buf_clk cell_8258 ( .C (clk), .D (signal_10803), .Q (signal_10804) ) ;
    buf_clk cell_8274 ( .C (clk), .D (signal_10819), .Q (signal_10820) ) ;
    buf_clk cell_8290 ( .C (clk), .D (signal_10835), .Q (signal_10836) ) ;
    buf_clk cell_8306 ( .C (clk), .D (signal_10851), .Q (signal_10852) ) ;
    buf_clk cell_8322 ( .C (clk), .D (signal_10867), .Q (signal_10868) ) ;
    buf_clk cell_8338 ( .C (clk), .D (signal_10883), .Q (signal_10884) ) ;
    buf_clk cell_8354 ( .C (clk), .D (signal_10899), .Q (signal_10900) ) ;
    buf_clk cell_8370 ( .C (clk), .D (signal_10915), .Q (signal_10916) ) ;
    buf_clk cell_8386 ( .C (clk), .D (signal_10931), .Q (signal_10932) ) ;
    buf_clk cell_8402 ( .C (clk), .D (signal_10947), .Q (signal_10948) ) ;
    buf_clk cell_8418 ( .C (clk), .D (signal_10963), .Q (signal_10964) ) ;
    buf_clk cell_8434 ( .C (clk), .D (signal_10979), .Q (signal_10980) ) ;
    buf_clk cell_8450 ( .C (clk), .D (signal_10995), .Q (signal_10996) ) ;
    buf_clk cell_8466 ( .C (clk), .D (signal_11011), .Q (signal_11012) ) ;
    buf_clk cell_8482 ( .C (clk), .D (signal_11027), .Q (signal_11028) ) ;
    buf_clk cell_8498 ( .C (clk), .D (signal_11043), .Q (signal_11044) ) ;
    buf_clk cell_8514 ( .C (clk), .D (signal_11059), .Q (signal_11060) ) ;
    buf_clk cell_8530 ( .C (clk), .D (signal_11075), .Q (signal_11076) ) ;
    buf_clk cell_8546 ( .C (clk), .D (signal_11091), .Q (signal_11092) ) ;
    buf_clk cell_8562 ( .C (clk), .D (signal_11107), .Q (signal_11108) ) ;
    buf_clk cell_8578 ( .C (clk), .D (signal_11123), .Q (signal_11124) ) ;
    buf_clk cell_8594 ( .C (clk), .D (signal_11139), .Q (signal_11140) ) ;
    buf_clk cell_8610 ( .C (clk), .D (signal_11155), .Q (signal_11156) ) ;
    buf_clk cell_8626 ( .C (clk), .D (signal_11171), .Q (signal_11172) ) ;
    buf_clk cell_8642 ( .C (clk), .D (signal_11187), .Q (signal_11188) ) ;
    buf_clk cell_8658 ( .C (clk), .D (signal_11203), .Q (signal_11204) ) ;
    buf_clk cell_8674 ( .C (clk), .D (signal_11219), .Q (signal_11220) ) ;
    buf_clk cell_8690 ( .C (clk), .D (signal_11235), .Q (signal_11236) ) ;
    buf_clk cell_8706 ( .C (clk), .D (signal_11251), .Q (signal_11252) ) ;
    buf_clk cell_8722 ( .C (clk), .D (signal_11267), .Q (signal_11268) ) ;
    buf_clk cell_8738 ( .C (clk), .D (signal_11283), .Q (signal_11284) ) ;
    buf_clk cell_8754 ( .C (clk), .D (signal_11299), .Q (signal_11300) ) ;
    buf_clk cell_8770 ( .C (clk), .D (signal_11315), .Q (signal_11316) ) ;
    buf_clk cell_8786 ( .C (clk), .D (signal_11331), .Q (signal_11332) ) ;
    buf_clk cell_8802 ( .C (clk), .D (signal_11347), .Q (signal_11348) ) ;
    buf_clk cell_8818 ( .C (clk), .D (signal_11363), .Q (signal_11364) ) ;
    buf_clk cell_8834 ( .C (clk), .D (signal_11379), .Q (signal_11380) ) ;
    buf_clk cell_8850 ( .C (clk), .D (signal_11395), .Q (signal_11396) ) ;
    buf_clk cell_8866 ( .C (clk), .D (signal_11411), .Q (signal_11412) ) ;
    buf_clk cell_8882 ( .C (clk), .D (signal_11427), .Q (signal_11428) ) ;
    buf_clk cell_8898 ( .C (clk), .D (signal_11443), .Q (signal_11444) ) ;
    buf_clk cell_8914 ( .C (clk), .D (signal_11459), .Q (signal_11460) ) ;
    buf_clk cell_8930 ( .C (clk), .D (signal_11475), .Q (signal_11476) ) ;
    buf_clk cell_8946 ( .C (clk), .D (signal_11491), .Q (signal_11492) ) ;
    buf_clk cell_8962 ( .C (clk), .D (signal_11507), .Q (signal_11508) ) ;
    buf_clk cell_8978 ( .C (clk), .D (signal_11523), .Q (signal_11524) ) ;
    buf_clk cell_8994 ( .C (clk), .D (signal_11539), .Q (signal_11540) ) ;
    buf_clk cell_9010 ( .C (clk), .D (signal_11555), .Q (signal_11556) ) ;
    buf_clk cell_9026 ( .C (clk), .D (signal_11571), .Q (signal_11572) ) ;
    buf_clk cell_9042 ( .C (clk), .D (signal_11587), .Q (signal_11588) ) ;
    buf_clk cell_9058 ( .C (clk), .D (signal_11603), .Q (signal_11604) ) ;
    buf_clk cell_9074 ( .C (clk), .D (signal_11619), .Q (signal_11620) ) ;
    buf_clk cell_9090 ( .C (clk), .D (signal_11635), .Q (signal_11636) ) ;
    buf_clk cell_9106 ( .C (clk), .D (signal_11651), .Q (signal_11652) ) ;
    buf_clk cell_9122 ( .C (clk), .D (signal_11667), .Q (signal_11668) ) ;
    buf_clk cell_9138 ( .C (clk), .D (signal_11683), .Q (signal_11684) ) ;
    buf_clk cell_9154 ( .C (clk), .D (signal_11699), .Q (signal_11700) ) ;
    buf_clk cell_9170 ( .C (clk), .D (signal_11715), .Q (signal_11716) ) ;
    buf_clk cell_9186 ( .C (clk), .D (signal_11731), .Q (signal_11732) ) ;
    buf_clk cell_9202 ( .C (clk), .D (signal_11747), .Q (signal_11748) ) ;
    buf_clk cell_9218 ( .C (clk), .D (signal_11763), .Q (signal_11764) ) ;
    buf_clk cell_9234 ( .C (clk), .D (signal_11779), .Q (signal_11780) ) ;
    buf_clk cell_9250 ( .C (clk), .D (signal_11795), .Q (signal_11796) ) ;
    buf_clk cell_9266 ( .C (clk), .D (signal_11811), .Q (signal_11812) ) ;
    buf_clk cell_9282 ( .C (clk), .D (signal_11827), .Q (signal_11828) ) ;
    buf_clk cell_9298 ( .C (clk), .D (signal_11843), .Q (signal_11844) ) ;
    buf_clk cell_9314 ( .C (clk), .D (signal_11859), .Q (signal_11860) ) ;
    buf_clk cell_9330 ( .C (clk), .D (signal_11875), .Q (signal_11876) ) ;
    buf_clk cell_9346 ( .C (clk), .D (signal_11891), .Q (signal_11892) ) ;
    buf_clk cell_9362 ( .C (clk), .D (signal_11907), .Q (signal_11908) ) ;
    buf_clk cell_9378 ( .C (clk), .D (signal_11923), .Q (signal_11924) ) ;
    buf_clk cell_9394 ( .C (clk), .D (signal_11939), .Q (signal_11940) ) ;
    buf_clk cell_9410 ( .C (clk), .D (signal_11955), .Q (signal_11956) ) ;
    buf_clk cell_9426 ( .C (clk), .D (signal_11971), .Q (signal_11972) ) ;
    buf_clk cell_9442 ( .C (clk), .D (signal_11987), .Q (signal_11988) ) ;
    buf_clk cell_9458 ( .C (clk), .D (signal_12003), .Q (signal_12004) ) ;
    buf_clk cell_9474 ( .C (clk), .D (signal_12019), .Q (signal_12020) ) ;
    buf_clk cell_9490 ( .C (clk), .D (signal_12035), .Q (signal_12036) ) ;
    buf_clk cell_9506 ( .C (clk), .D (signal_12051), .Q (signal_12052) ) ;
    buf_clk cell_9522 ( .C (clk), .D (signal_12067), .Q (signal_12068) ) ;
    buf_clk cell_9538 ( .C (clk), .D (signal_12083), .Q (signal_12084) ) ;
    buf_clk cell_9554 ( .C (clk), .D (signal_12099), .Q (signal_12100) ) ;
    buf_clk cell_9570 ( .C (clk), .D (signal_12115), .Q (signal_12116) ) ;
    buf_clk cell_9586 ( .C (clk), .D (signal_12131), .Q (signal_12132) ) ;
    buf_clk cell_9602 ( .C (clk), .D (signal_12147), .Q (signal_12148) ) ;
    buf_clk cell_9618 ( .C (clk), .D (signal_12163), .Q (signal_12164) ) ;
    buf_clk cell_9634 ( .C (clk), .D (signal_12179), .Q (signal_12180) ) ;
    buf_clk cell_9650 ( .C (clk), .D (signal_12195), .Q (signal_12196) ) ;
    buf_clk cell_9666 ( .C (clk), .D (signal_12211), .Q (signal_12212) ) ;
    buf_clk cell_9682 ( .C (clk), .D (signal_12227), .Q (signal_12228) ) ;
    buf_clk cell_9698 ( .C (clk), .D (signal_12243), .Q (signal_12244) ) ;
    buf_clk cell_9714 ( .C (clk), .D (signal_12259), .Q (signal_12260) ) ;
    buf_clk cell_9730 ( .C (clk), .D (signal_12275), .Q (signal_12276) ) ;
    buf_clk cell_9746 ( .C (clk), .D (signal_12291), .Q (signal_12292) ) ;
    buf_clk cell_9762 ( .C (clk), .D (signal_12307), .Q (signal_12308) ) ;
    buf_clk cell_9778 ( .C (clk), .D (signal_12323), .Q (signal_12324) ) ;
    buf_clk cell_9794 ( .C (clk), .D (signal_12339), .Q (signal_12340) ) ;
    buf_clk cell_9810 ( .C (clk), .D (signal_12355), .Q (signal_12356) ) ;
    buf_clk cell_9826 ( .C (clk), .D (signal_12371), .Q (signal_12372) ) ;
    buf_clk cell_9842 ( .C (clk), .D (signal_12387), .Q (signal_12388) ) ;
    buf_clk cell_9858 ( .C (clk), .D (signal_12403), .Q (signal_12404) ) ;
    buf_clk cell_9874 ( .C (clk), .D (signal_12419), .Q (signal_12420) ) ;
    buf_clk cell_9890 ( .C (clk), .D (signal_12435), .Q (signal_12436) ) ;
    buf_clk cell_9906 ( .C (clk), .D (signal_12451), .Q (signal_12452) ) ;
    buf_clk cell_9922 ( .C (clk), .D (signal_12467), .Q (signal_12468) ) ;
    buf_clk cell_9938 ( .C (clk), .D (signal_12483), .Q (signal_12484) ) ;
    buf_clk cell_9954 ( .C (clk), .D (signal_12499), .Q (signal_12500) ) ;
    buf_clk cell_9970 ( .C (clk), .D (signal_12515), .Q (signal_12516) ) ;
    buf_clk cell_9986 ( .C (clk), .D (signal_12531), .Q (signal_12532) ) ;
    buf_clk cell_10002 ( .C (clk), .D (signal_12547), .Q (signal_12548) ) ;
    buf_clk cell_10018 ( .C (clk), .D (signal_12563), .Q (signal_12564) ) ;
    buf_clk cell_10034 ( .C (clk), .D (signal_12579), .Q (signal_12580) ) ;
    buf_clk cell_10050 ( .C (clk), .D (signal_12595), .Q (signal_12596) ) ;
    buf_clk cell_10066 ( .C (clk), .D (signal_12611), .Q (signal_12612) ) ;
    buf_clk cell_10082 ( .C (clk), .D (signal_12627), .Q (signal_12628) ) ;
    buf_clk cell_10098 ( .C (clk), .D (signal_12643), .Q (signal_12644) ) ;
    buf_clk cell_10114 ( .C (clk), .D (signal_12659), .Q (signal_12660) ) ;
    buf_clk cell_10130 ( .C (clk), .D (signal_12675), .Q (signal_12676) ) ;
    buf_clk cell_10146 ( .C (clk), .D (signal_12691), .Q (signal_12692) ) ;
    buf_clk cell_10162 ( .C (clk), .D (signal_12707), .Q (signal_12708) ) ;
    buf_clk cell_10178 ( .C (clk), .D (signal_12723), .Q (signal_12724) ) ;
    buf_clk cell_10194 ( .C (clk), .D (signal_12739), .Q (signal_12740) ) ;
    buf_clk cell_10210 ( .C (clk), .D (signal_12755), .Q (signal_12756) ) ;
    buf_clk cell_10226 ( .C (clk), .D (signal_12771), .Q (signal_12772) ) ;
    buf_clk cell_10242 ( .C (clk), .D (signal_12787), .Q (signal_12788) ) ;
    buf_clk cell_10258 ( .C (clk), .D (signal_12803), .Q (signal_12804) ) ;
    buf_clk cell_10274 ( .C (clk), .D (signal_12819), .Q (signal_12820) ) ;
    buf_clk cell_10290 ( .C (clk), .D (signal_12835), .Q (signal_12836) ) ;
    buf_clk cell_10306 ( .C (clk), .D (signal_12851), .Q (signal_12852) ) ;
    buf_clk cell_10322 ( .C (clk), .D (signal_12867), .Q (signal_12868) ) ;
    buf_clk cell_10338 ( .C (clk), .D (signal_12883), .Q (signal_12884) ) ;
    buf_clk cell_10354 ( .C (clk), .D (signal_12899), .Q (signal_12900) ) ;
    buf_clk cell_10370 ( .C (clk), .D (signal_12915), .Q (signal_12916) ) ;
    buf_clk cell_10386 ( .C (clk), .D (signal_12931), .Q (signal_12932) ) ;
    buf_clk cell_10402 ( .C (clk), .D (signal_12947), .Q (signal_12948) ) ;
    buf_clk cell_10418 ( .C (clk), .D (signal_12963), .Q (signal_12964) ) ;
    buf_clk cell_10434 ( .C (clk), .D (signal_12979), .Q (signal_12980) ) ;
    buf_clk cell_10450 ( .C (clk), .D (signal_12995), .Q (signal_12996) ) ;
    buf_clk cell_10466 ( .C (clk), .D (signal_13011), .Q (signal_13012) ) ;
    buf_clk cell_10482 ( .C (clk), .D (signal_13027), .Q (signal_13028) ) ;
    buf_clk cell_10498 ( .C (clk), .D (signal_13043), .Q (signal_13044) ) ;
    buf_clk cell_10514 ( .C (clk), .D (signal_13059), .Q (signal_13060) ) ;
    buf_clk cell_10530 ( .C (clk), .D (signal_13075), .Q (signal_13076) ) ;
    buf_clk cell_10546 ( .C (clk), .D (signal_13091), .Q (signal_13092) ) ;
    buf_clk cell_10562 ( .C (clk), .D (signal_13107), .Q (signal_13108) ) ;
    buf_clk cell_10578 ( .C (clk), .D (signal_13123), .Q (signal_13124) ) ;
    buf_clk cell_10594 ( .C (clk), .D (signal_13139), .Q (signal_13140) ) ;
    buf_clk cell_10610 ( .C (clk), .D (signal_13155), .Q (signal_13156) ) ;
    buf_clk cell_10626 ( .C (clk), .D (signal_13171), .Q (signal_13172) ) ;
    buf_clk cell_10642 ( .C (clk), .D (signal_13187), .Q (signal_13188) ) ;
    buf_clk cell_10658 ( .C (clk), .D (signal_13203), .Q (signal_13204) ) ;
    buf_clk cell_10674 ( .C (clk), .D (signal_13219), .Q (signal_13220) ) ;
    buf_clk cell_10690 ( .C (clk), .D (signal_13235), .Q (signal_13236) ) ;
    buf_clk cell_10706 ( .C (clk), .D (signal_13251), .Q (signal_13252) ) ;
    buf_clk cell_10722 ( .C (clk), .D (signal_13267), .Q (signal_13268) ) ;
    buf_clk cell_10738 ( .C (clk), .D (signal_13283), .Q (signal_13284) ) ;
    buf_clk cell_10754 ( .C (clk), .D (signal_13299), .Q (signal_13300) ) ;
    buf_clk cell_10770 ( .C (clk), .D (signal_13315), .Q (signal_13316) ) ;
    buf_clk cell_10786 ( .C (clk), .D (signal_13331), .Q (signal_13332) ) ;
    buf_clk cell_10802 ( .C (clk), .D (signal_13347), .Q (signal_13348) ) ;
    buf_clk cell_10818 ( .C (clk), .D (signal_13363), .Q (signal_13364) ) ;
    buf_clk cell_10834 ( .C (clk), .D (signal_13379), .Q (signal_13380) ) ;
    buf_clk cell_10850 ( .C (clk), .D (signal_13395), .Q (signal_13396) ) ;
    buf_clk cell_10866 ( .C (clk), .D (signal_13411), .Q (signal_13412) ) ;
    buf_clk cell_10882 ( .C (clk), .D (signal_13427), .Q (signal_13428) ) ;
    buf_clk cell_10898 ( .C (clk), .D (signal_13443), .Q (signal_13444) ) ;
    buf_clk cell_10914 ( .C (clk), .D (signal_13459), .Q (signal_13460) ) ;
    buf_clk cell_10930 ( .C (clk), .D (signal_13475), .Q (signal_13476) ) ;
    buf_clk cell_10946 ( .C (clk), .D (signal_13491), .Q (signal_13492) ) ;
    buf_clk cell_10962 ( .C (clk), .D (signal_13507), .Q (signal_13508) ) ;
    buf_clk cell_10978 ( .C (clk), .D (signal_13523), .Q (signal_13524) ) ;
    buf_clk cell_10994 ( .C (clk), .D (signal_13539), .Q (signal_13540) ) ;
    buf_clk cell_11010 ( .C (clk), .D (signal_13555), .Q (signal_13556) ) ;
    buf_clk cell_11026 ( .C (clk), .D (signal_13571), .Q (signal_13572) ) ;
    buf_clk cell_11042 ( .C (clk), .D (signal_13587), .Q (signal_13588) ) ;
    buf_clk cell_11058 ( .C (clk), .D (signal_13603), .Q (signal_13604) ) ;
    buf_clk cell_11074 ( .C (clk), .D (signal_13619), .Q (signal_13620) ) ;
    buf_clk cell_11090 ( .C (clk), .D (signal_13635), .Q (signal_13636) ) ;
    buf_clk cell_11106 ( .C (clk), .D (signal_13651), .Q (signal_13652) ) ;
    buf_clk cell_11122 ( .C (clk), .D (signal_13667), .Q (signal_13668) ) ;
    buf_clk cell_11138 ( .C (clk), .D (signal_13683), .Q (signal_13684) ) ;
    buf_clk cell_11154 ( .C (clk), .D (signal_13699), .Q (signal_13700) ) ;
    buf_clk cell_11170 ( .C (clk), .D (signal_13715), .Q (signal_13716) ) ;
    buf_clk cell_11186 ( .C (clk), .D (signal_13731), .Q (signal_13732) ) ;
    buf_clk cell_11202 ( .C (clk), .D (signal_13747), .Q (signal_13748) ) ;
    buf_clk cell_11218 ( .C (clk), .D (signal_13763), .Q (signal_13764) ) ;
    buf_clk cell_11234 ( .C (clk), .D (signal_13779), .Q (signal_13780) ) ;
    buf_clk cell_11250 ( .C (clk), .D (signal_13795), .Q (signal_13796) ) ;
    buf_clk cell_11266 ( .C (clk), .D (signal_13811), .Q (signal_13812) ) ;
    buf_clk cell_11282 ( .C (clk), .D (signal_13827), .Q (signal_13828) ) ;
    buf_clk cell_11298 ( .C (clk), .D (signal_13843), .Q (signal_13844) ) ;
    buf_clk cell_11314 ( .C (clk), .D (signal_13859), .Q (signal_13860) ) ;
    buf_clk cell_11330 ( .C (clk), .D (signal_13875), .Q (signal_13876) ) ;
    buf_clk cell_11346 ( .C (clk), .D (signal_13891), .Q (signal_13892) ) ;
    buf_clk cell_11362 ( .C (clk), .D (signal_13907), .Q (signal_13908) ) ;
    buf_clk cell_11378 ( .C (clk), .D (signal_13923), .Q (signal_13924) ) ;
    buf_clk cell_11394 ( .C (clk), .D (signal_13939), .Q (signal_13940) ) ;
    buf_clk cell_11410 ( .C (clk), .D (signal_13955), .Q (signal_13956) ) ;
    buf_clk cell_11426 ( .C (clk), .D (signal_13971), .Q (signal_13972) ) ;
    buf_clk cell_11442 ( .C (clk), .D (signal_13987), .Q (signal_13988) ) ;
    buf_clk cell_11458 ( .C (clk), .D (signal_14003), .Q (signal_14004) ) ;
    buf_clk cell_11474 ( .C (clk), .D (signal_14019), .Q (signal_14020) ) ;
    buf_clk cell_11490 ( .C (clk), .D (signal_14035), .Q (signal_14036) ) ;
    buf_clk cell_11506 ( .C (clk), .D (signal_14051), .Q (signal_14052) ) ;
    buf_clk cell_11522 ( .C (clk), .D (signal_14067), .Q (signal_14068) ) ;
    buf_clk cell_11538 ( .C (clk), .D (signal_14083), .Q (signal_14084) ) ;
    buf_clk cell_11554 ( .C (clk), .D (signal_14099), .Q (signal_14100) ) ;
    buf_clk cell_11570 ( .C (clk), .D (signal_14115), .Q (signal_14116) ) ;
    buf_clk cell_11586 ( .C (clk), .D (signal_14131), .Q (signal_14132) ) ;
    buf_clk cell_11602 ( .C (clk), .D (signal_14147), .Q (signal_14148) ) ;
    buf_clk cell_11618 ( .C (clk), .D (signal_14163), .Q (signal_14164) ) ;
    buf_clk cell_11634 ( .C (clk), .D (signal_14179), .Q (signal_14180) ) ;
    buf_clk cell_11650 ( .C (clk), .D (signal_14195), .Q (signal_14196) ) ;
    buf_clk cell_11666 ( .C (clk), .D (signal_14211), .Q (signal_14212) ) ;
    buf_clk cell_11682 ( .C (clk), .D (signal_14227), .Q (signal_14228) ) ;
    buf_clk cell_11698 ( .C (clk), .D (signal_14243), .Q (signal_14244) ) ;
    buf_clk cell_11714 ( .C (clk), .D (signal_14259), .Q (signal_14260) ) ;
    buf_clk cell_11730 ( .C (clk), .D (signal_14275), .Q (signal_14276) ) ;
    buf_clk cell_11746 ( .C (clk), .D (signal_14291), .Q (signal_14292) ) ;
    buf_clk cell_11762 ( .C (clk), .D (signal_14307), .Q (signal_14308) ) ;
    buf_clk cell_11778 ( .C (clk), .D (signal_14323), .Q (signal_14324) ) ;
    buf_clk cell_11794 ( .C (clk), .D (signal_14339), .Q (signal_14340) ) ;
    buf_clk cell_11810 ( .C (clk), .D (signal_14355), .Q (signal_14356) ) ;
    buf_clk cell_11826 ( .C (clk), .D (signal_14371), .Q (signal_14372) ) ;
    buf_clk cell_11842 ( .C (clk), .D (signal_14387), .Q (signal_14388) ) ;
    buf_clk cell_11858 ( .C (clk), .D (signal_14403), .Q (signal_14404) ) ;
    buf_clk cell_11874 ( .C (clk), .D (signal_14419), .Q (signal_14420) ) ;
    buf_clk cell_11890 ( .C (clk), .D (signal_14435), .Q (signal_14436) ) ;
    buf_clk cell_11906 ( .C (clk), .D (signal_14451), .Q (signal_14452) ) ;
    buf_clk cell_11922 ( .C (clk), .D (signal_14467), .Q (signal_14468) ) ;
    buf_clk cell_11938 ( .C (clk), .D (signal_14483), .Q (signal_14484) ) ;
    buf_clk cell_11954 ( .C (clk), .D (signal_14499), .Q (signal_14500) ) ;
    buf_clk cell_11970 ( .C (clk), .D (signal_14515), .Q (signal_14516) ) ;
    buf_clk cell_11986 ( .C (clk), .D (signal_14531), .Q (signal_14532) ) ;
    buf_clk cell_12002 ( .C (clk), .D (signal_14547), .Q (signal_14548) ) ;
    buf_clk cell_12018 ( .C (clk), .D (signal_14563), .Q (signal_14564) ) ;
    buf_clk cell_12034 ( .C (clk), .D (signal_14579), .Q (signal_14580) ) ;
    buf_clk cell_12050 ( .C (clk), .D (signal_14595), .Q (signal_14596) ) ;
    buf_clk cell_12066 ( .C (clk), .D (signal_14611), .Q (signal_14612) ) ;
    buf_clk cell_12082 ( .C (clk), .D (signal_14627), .Q (signal_14628) ) ;
    buf_clk cell_12098 ( .C (clk), .D (signal_14643), .Q (signal_14644) ) ;
    buf_clk cell_12114 ( .C (clk), .D (signal_14659), .Q (signal_14660) ) ;
    buf_clk cell_12130 ( .C (clk), .D (signal_14675), .Q (signal_14676) ) ;
    buf_clk cell_12146 ( .C (clk), .D (signal_14691), .Q (signal_14692) ) ;
    buf_clk cell_12162 ( .C (clk), .D (signal_14707), .Q (signal_14708) ) ;
    buf_clk cell_12178 ( .C (clk), .D (signal_14723), .Q (signal_14724) ) ;
    buf_clk cell_12194 ( .C (clk), .D (signal_14739), .Q (signal_14740) ) ;
    buf_clk cell_12210 ( .C (clk), .D (signal_14755), .Q (signal_14756) ) ;
    buf_clk cell_12226 ( .C (clk), .D (signal_14771), .Q (signal_14772) ) ;
    buf_clk cell_12242 ( .C (clk), .D (signal_14787), .Q (signal_14788) ) ;
    buf_clk cell_12258 ( .C (clk), .D (signal_14803), .Q (signal_14804) ) ;
    buf_clk cell_12274 ( .C (clk), .D (signal_14819), .Q (signal_14820) ) ;
    buf_clk cell_12290 ( .C (clk), .D (signal_14835), .Q (signal_14836) ) ;
    buf_clk cell_12306 ( .C (clk), .D (signal_14851), .Q (signal_14852) ) ;
    buf_clk cell_12322 ( .C (clk), .D (signal_14867), .Q (signal_14868) ) ;
    buf_clk cell_12338 ( .C (clk), .D (signal_14883), .Q (signal_14884) ) ;
    buf_clk cell_12354 ( .C (clk), .D (signal_14899), .Q (signal_14900) ) ;
    buf_clk cell_12370 ( .C (clk), .D (signal_14915), .Q (signal_14916) ) ;
    buf_clk cell_12386 ( .C (clk), .D (signal_14931), .Q (signal_14932) ) ;

    /* cells in depth 7 */
    buf_clk cell_2303 ( .C (clk), .D (signal_4848), .Q (signal_4849) ) ;
    buf_clk cell_2311 ( .C (clk), .D (signal_4856), .Q (signal_4857) ) ;
    buf_clk cell_2313 ( .C (clk), .D (signal_2035), .Q (signal_4859) ) ;
    buf_clk cell_2315 ( .C (clk), .D (signal_3490), .Q (signal_4861) ) ;
    buf_clk cell_2317 ( .C (clk), .D (signal_2040), .Q (signal_4863) ) ;
    buf_clk cell_2319 ( .C (clk), .D (signal_3495), .Q (signal_4865) ) ;
    buf_clk cell_2321 ( .C (clk), .D (signal_2042), .Q (signal_4867) ) ;
    buf_clk cell_2323 ( .C (clk), .D (signal_3497), .Q (signal_4869) ) ;
    buf_clk cell_2325 ( .C (clk), .D (signal_2097), .Q (signal_4871) ) ;
    buf_clk cell_2327 ( .C (clk), .D (signal_3552), .Q (signal_4873) ) ;
    buf_clk cell_2329 ( .C (clk), .D (signal_2116), .Q (signal_4875) ) ;
    buf_clk cell_2331 ( .C (clk), .D (signal_3571), .Q (signal_4877) ) ;
    buf_clk cell_2333 ( .C (clk), .D (signal_2146), .Q (signal_4879) ) ;
    buf_clk cell_2335 ( .C (clk), .D (signal_3601), .Q (signal_4881) ) ;
    buf_clk cell_2337 ( .C (clk), .D (signal_2147), .Q (signal_4883) ) ;
    buf_clk cell_2339 ( .C (clk), .D (signal_3602), .Q (signal_4885) ) ;
    buf_clk cell_2347 ( .C (clk), .D (signal_4892), .Q (signal_4893) ) ;
    buf_clk cell_2357 ( .C (clk), .D (signal_4902), .Q (signal_4903) ) ;
    buf_clk cell_2367 ( .C (clk), .D (signal_4912), .Q (signal_4913) ) ;
    buf_clk cell_2379 ( .C (clk), .D (signal_4924), .Q (signal_4925) ) ;
    buf_clk cell_2391 ( .C (clk), .D (signal_4936), .Q (signal_4937) ) ;
    buf_clk cell_2407 ( .C (clk), .D (signal_4952), .Q (signal_4953) ) ;
    buf_clk cell_2423 ( .C (clk), .D (signal_4968), .Q (signal_4969) ) ;
    buf_clk cell_2439 ( .C (clk), .D (signal_4984), .Q (signal_4985) ) ;
    buf_clk cell_2455 ( .C (clk), .D (signal_5000), .Q (signal_5001) ) ;
    buf_clk cell_2471 ( .C (clk), .D (signal_5016), .Q (signal_5017) ) ;
    buf_clk cell_2487 ( .C (clk), .D (signal_5032), .Q (signal_5033) ) ;
    buf_clk cell_2503 ( .C (clk), .D (signal_5048), .Q (signal_5049) ) ;
    buf_clk cell_2519 ( .C (clk), .D (signal_5064), .Q (signal_5065) ) ;
    buf_clk cell_2535 ( .C (clk), .D (signal_5080), .Q (signal_5081) ) ;
    buf_clk cell_2551 ( .C (clk), .D (signal_5096), .Q (signal_5097) ) ;
    buf_clk cell_2567 ( .C (clk), .D (signal_5112), .Q (signal_5113) ) ;
    buf_clk cell_2583 ( .C (clk), .D (signal_5128), .Q (signal_5129) ) ;
    buf_clk cell_2599 ( .C (clk), .D (signal_5144), .Q (signal_5145) ) ;
    buf_clk cell_2615 ( .C (clk), .D (signal_5160), .Q (signal_5161) ) ;
    buf_clk cell_2631 ( .C (clk), .D (signal_5176), .Q (signal_5177) ) ;
    buf_clk cell_2647 ( .C (clk), .D (signal_5192), .Q (signal_5193) ) ;
    buf_clk cell_2663 ( .C (clk), .D (signal_5208), .Q (signal_5209) ) ;
    buf_clk cell_2679 ( .C (clk), .D (signal_5224), .Q (signal_5225) ) ;
    buf_clk cell_2695 ( .C (clk), .D (signal_5240), .Q (signal_5241) ) ;
    buf_clk cell_2711 ( .C (clk), .D (signal_5256), .Q (signal_5257) ) ;
    buf_clk cell_2727 ( .C (clk), .D (signal_5272), .Q (signal_5273) ) ;
    buf_clk cell_2743 ( .C (clk), .D (signal_5288), .Q (signal_5289) ) ;
    buf_clk cell_2759 ( .C (clk), .D (signal_5304), .Q (signal_5305) ) ;
    buf_clk cell_2775 ( .C (clk), .D (signal_5320), .Q (signal_5321) ) ;
    buf_clk cell_2791 ( .C (clk), .D (signal_5336), .Q (signal_5337) ) ;
    buf_clk cell_2807 ( .C (clk), .D (signal_5352), .Q (signal_5353) ) ;
    buf_clk cell_2823 ( .C (clk), .D (signal_5368), .Q (signal_5369) ) ;
    buf_clk cell_2839 ( .C (clk), .D (signal_5384), .Q (signal_5385) ) ;
    buf_clk cell_2855 ( .C (clk), .D (signal_5400), .Q (signal_5401) ) ;
    buf_clk cell_2871 ( .C (clk), .D (signal_5416), .Q (signal_5417) ) ;
    buf_clk cell_2887 ( .C (clk), .D (signal_5432), .Q (signal_5433) ) ;
    buf_clk cell_2903 ( .C (clk), .D (signal_5448), .Q (signal_5449) ) ;
    buf_clk cell_2919 ( .C (clk), .D (signal_5464), .Q (signal_5465) ) ;
    buf_clk cell_2935 ( .C (clk), .D (signal_5480), .Q (signal_5481) ) ;
    buf_clk cell_2951 ( .C (clk), .D (signal_5496), .Q (signal_5497) ) ;
    buf_clk cell_2967 ( .C (clk), .D (signal_5512), .Q (signal_5513) ) ;
    buf_clk cell_2983 ( .C (clk), .D (signal_5528), .Q (signal_5529) ) ;
    buf_clk cell_2999 ( .C (clk), .D (signal_5544), .Q (signal_5545) ) ;
    buf_clk cell_3015 ( .C (clk), .D (signal_5560), .Q (signal_5561) ) ;
    buf_clk cell_3031 ( .C (clk), .D (signal_5576), .Q (signal_5577) ) ;
    buf_clk cell_3047 ( .C (clk), .D (signal_5592), .Q (signal_5593) ) ;
    buf_clk cell_3063 ( .C (clk), .D (signal_5608), .Q (signal_5609) ) ;
    buf_clk cell_3079 ( .C (clk), .D (signal_5624), .Q (signal_5625) ) ;
    buf_clk cell_3095 ( .C (clk), .D (signal_5640), .Q (signal_5641) ) ;
    buf_clk cell_3111 ( .C (clk), .D (signal_5656), .Q (signal_5657) ) ;
    buf_clk cell_3127 ( .C (clk), .D (signal_5672), .Q (signal_5673) ) ;
    buf_clk cell_3143 ( .C (clk), .D (signal_5688), .Q (signal_5689) ) ;
    buf_clk cell_3159 ( .C (clk), .D (signal_5704), .Q (signal_5705) ) ;
    buf_clk cell_3175 ( .C (clk), .D (signal_5720), .Q (signal_5721) ) ;
    buf_clk cell_3191 ( .C (clk), .D (signal_5736), .Q (signal_5737) ) ;
    buf_clk cell_3207 ( .C (clk), .D (signal_5752), .Q (signal_5753) ) ;
    buf_clk cell_3223 ( .C (clk), .D (signal_5768), .Q (signal_5769) ) ;
    buf_clk cell_3239 ( .C (clk), .D (signal_5784), .Q (signal_5785) ) ;
    buf_clk cell_3255 ( .C (clk), .D (signal_5800), .Q (signal_5801) ) ;
    buf_clk cell_3271 ( .C (clk), .D (signal_5816), .Q (signal_5817) ) ;
    buf_clk cell_3287 ( .C (clk), .D (signal_5832), .Q (signal_5833) ) ;
    buf_clk cell_3303 ( .C (clk), .D (signal_5848), .Q (signal_5849) ) ;
    buf_clk cell_3319 ( .C (clk), .D (signal_5864), .Q (signal_5865) ) ;
    buf_clk cell_3335 ( .C (clk), .D (signal_5880), .Q (signal_5881) ) ;
    buf_clk cell_3351 ( .C (clk), .D (signal_5896), .Q (signal_5897) ) ;
    buf_clk cell_3367 ( .C (clk), .D (signal_5912), .Q (signal_5913) ) ;
    buf_clk cell_3383 ( .C (clk), .D (signal_5928), .Q (signal_5929) ) ;
    buf_clk cell_3399 ( .C (clk), .D (signal_5944), .Q (signal_5945) ) ;
    buf_clk cell_3415 ( .C (clk), .D (signal_5960), .Q (signal_5961) ) ;
    buf_clk cell_3431 ( .C (clk), .D (signal_5976), .Q (signal_5977) ) ;
    buf_clk cell_3447 ( .C (clk), .D (signal_5992), .Q (signal_5993) ) ;
    buf_clk cell_3463 ( .C (clk), .D (signal_6008), .Q (signal_6009) ) ;
    buf_clk cell_3479 ( .C (clk), .D (signal_6024), .Q (signal_6025) ) ;
    buf_clk cell_3495 ( .C (clk), .D (signal_6040), .Q (signal_6041) ) ;
    buf_clk cell_3511 ( .C (clk), .D (signal_6056), .Q (signal_6057) ) ;
    buf_clk cell_3527 ( .C (clk), .D (signal_6072), .Q (signal_6073) ) ;
    buf_clk cell_3543 ( .C (clk), .D (signal_6088), .Q (signal_6089) ) ;
    buf_clk cell_3559 ( .C (clk), .D (signal_6104), .Q (signal_6105) ) ;
    buf_clk cell_3575 ( .C (clk), .D (signal_6120), .Q (signal_6121) ) ;
    buf_clk cell_3591 ( .C (clk), .D (signal_6136), .Q (signal_6137) ) ;
    buf_clk cell_3607 ( .C (clk), .D (signal_6152), .Q (signal_6153) ) ;
    buf_clk cell_3623 ( .C (clk), .D (signal_6168), .Q (signal_6169) ) ;
    buf_clk cell_3639 ( .C (clk), .D (signal_6184), .Q (signal_6185) ) ;
    buf_clk cell_3655 ( .C (clk), .D (signal_6200), .Q (signal_6201) ) ;
    buf_clk cell_3671 ( .C (clk), .D (signal_6216), .Q (signal_6217) ) ;
    buf_clk cell_3687 ( .C (clk), .D (signal_6232), .Q (signal_6233) ) ;
    buf_clk cell_3703 ( .C (clk), .D (signal_6248), .Q (signal_6249) ) ;
    buf_clk cell_3719 ( .C (clk), .D (signal_6264), .Q (signal_6265) ) ;
    buf_clk cell_3735 ( .C (clk), .D (signal_6280), .Q (signal_6281) ) ;
    buf_clk cell_3751 ( .C (clk), .D (signal_6296), .Q (signal_6297) ) ;
    buf_clk cell_3767 ( .C (clk), .D (signal_6312), .Q (signal_6313) ) ;
    buf_clk cell_3783 ( .C (clk), .D (signal_6328), .Q (signal_6329) ) ;
    buf_clk cell_3799 ( .C (clk), .D (signal_6344), .Q (signal_6345) ) ;
    buf_clk cell_3815 ( .C (clk), .D (signal_6360), .Q (signal_6361) ) ;
    buf_clk cell_3831 ( .C (clk), .D (signal_6376), .Q (signal_6377) ) ;
    buf_clk cell_3847 ( .C (clk), .D (signal_6392), .Q (signal_6393) ) ;
    buf_clk cell_3863 ( .C (clk), .D (signal_6408), .Q (signal_6409) ) ;
    buf_clk cell_3879 ( .C (clk), .D (signal_6424), .Q (signal_6425) ) ;
    buf_clk cell_3895 ( .C (clk), .D (signal_6440), .Q (signal_6441) ) ;
    buf_clk cell_3911 ( .C (clk), .D (signal_6456), .Q (signal_6457) ) ;
    buf_clk cell_3927 ( .C (clk), .D (signal_6472), .Q (signal_6473) ) ;
    buf_clk cell_3943 ( .C (clk), .D (signal_6488), .Q (signal_6489) ) ;
    buf_clk cell_3959 ( .C (clk), .D (signal_6504), .Q (signal_6505) ) ;
    buf_clk cell_3975 ( .C (clk), .D (signal_6520), .Q (signal_6521) ) ;
    buf_clk cell_3991 ( .C (clk), .D (signal_6536), .Q (signal_6537) ) ;
    buf_clk cell_4007 ( .C (clk), .D (signal_6552), .Q (signal_6553) ) ;
    buf_clk cell_4023 ( .C (clk), .D (signal_6568), .Q (signal_6569) ) ;
    buf_clk cell_4039 ( .C (clk), .D (signal_6584), .Q (signal_6585) ) ;
    buf_clk cell_4055 ( .C (clk), .D (signal_6600), .Q (signal_6601) ) ;
    buf_clk cell_4071 ( .C (clk), .D (signal_6616), .Q (signal_6617) ) ;
    buf_clk cell_4087 ( .C (clk), .D (signal_6632), .Q (signal_6633) ) ;
    buf_clk cell_4103 ( .C (clk), .D (signal_6648), .Q (signal_6649) ) ;
    buf_clk cell_4119 ( .C (clk), .D (signal_6664), .Q (signal_6665) ) ;
    buf_clk cell_4135 ( .C (clk), .D (signal_6680), .Q (signal_6681) ) ;
    buf_clk cell_4151 ( .C (clk), .D (signal_6696), .Q (signal_6697) ) ;
    buf_clk cell_4167 ( .C (clk), .D (signal_6712), .Q (signal_6713) ) ;
    buf_clk cell_4183 ( .C (clk), .D (signal_6728), .Q (signal_6729) ) ;
    buf_clk cell_4199 ( .C (clk), .D (signal_6744), .Q (signal_6745) ) ;
    buf_clk cell_4215 ( .C (clk), .D (signal_6760), .Q (signal_6761) ) ;
    buf_clk cell_4231 ( .C (clk), .D (signal_6776), .Q (signal_6777) ) ;
    buf_clk cell_4247 ( .C (clk), .D (signal_6792), .Q (signal_6793) ) ;
    buf_clk cell_4263 ( .C (clk), .D (signal_6808), .Q (signal_6809) ) ;
    buf_clk cell_4279 ( .C (clk), .D (signal_6824), .Q (signal_6825) ) ;
    buf_clk cell_4295 ( .C (clk), .D (signal_6840), .Q (signal_6841) ) ;
    buf_clk cell_4311 ( .C (clk), .D (signal_6856), .Q (signal_6857) ) ;
    buf_clk cell_4327 ( .C (clk), .D (signal_6872), .Q (signal_6873) ) ;
    buf_clk cell_4343 ( .C (clk), .D (signal_6888), .Q (signal_6889) ) ;
    buf_clk cell_4359 ( .C (clk), .D (signal_6904), .Q (signal_6905) ) ;
    buf_clk cell_4375 ( .C (clk), .D (signal_6920), .Q (signal_6921) ) ;
    buf_clk cell_4391 ( .C (clk), .D (signal_6936), .Q (signal_6937) ) ;
    buf_clk cell_4407 ( .C (clk), .D (signal_6952), .Q (signal_6953) ) ;
    buf_clk cell_4421 ( .C (clk), .D (signal_6966), .Q (signal_6967) ) ;
    buf_clk cell_4435 ( .C (clk), .D (signal_6980), .Q (signal_6981) ) ;
    buf_clk cell_4451 ( .C (clk), .D (signal_6996), .Q (signal_6997) ) ;
    buf_clk cell_4467 ( .C (clk), .D (signal_7012), .Q (signal_7013) ) ;
    buf_clk cell_4483 ( .C (clk), .D (signal_7028), .Q (signal_7029) ) ;
    buf_clk cell_4499 ( .C (clk), .D (signal_7044), .Q (signal_7045) ) ;
    buf_clk cell_4515 ( .C (clk), .D (signal_7060), .Q (signal_7061) ) ;
    buf_clk cell_4531 ( .C (clk), .D (signal_7076), .Q (signal_7077) ) ;
    buf_clk cell_4547 ( .C (clk), .D (signal_7092), .Q (signal_7093) ) ;
    buf_clk cell_4563 ( .C (clk), .D (signal_7108), .Q (signal_7109) ) ;
    buf_clk cell_4579 ( .C (clk), .D (signal_7124), .Q (signal_7125) ) ;
    buf_clk cell_4595 ( .C (clk), .D (signal_7140), .Q (signal_7141) ) ;
    buf_clk cell_4611 ( .C (clk), .D (signal_7156), .Q (signal_7157) ) ;
    buf_clk cell_4627 ( .C (clk), .D (signal_7172), .Q (signal_7173) ) ;
    buf_clk cell_4643 ( .C (clk), .D (signal_7188), .Q (signal_7189) ) ;
    buf_clk cell_4659 ( .C (clk), .D (signal_7204), .Q (signal_7205) ) ;
    buf_clk cell_4675 ( .C (clk), .D (signal_7220), .Q (signal_7221) ) ;
    buf_clk cell_4691 ( .C (clk), .D (signal_7236), .Q (signal_7237) ) ;
    buf_clk cell_4707 ( .C (clk), .D (signal_7252), .Q (signal_7253) ) ;
    buf_clk cell_4723 ( .C (clk), .D (signal_7268), .Q (signal_7269) ) ;
    buf_clk cell_4739 ( .C (clk), .D (signal_7284), .Q (signal_7285) ) ;
    buf_clk cell_4755 ( .C (clk), .D (signal_7300), .Q (signal_7301) ) ;
    buf_clk cell_4771 ( .C (clk), .D (signal_7316), .Q (signal_7317) ) ;
    buf_clk cell_4787 ( .C (clk), .D (signal_7332), .Q (signal_7333) ) ;
    buf_clk cell_4803 ( .C (clk), .D (signal_7348), .Q (signal_7349) ) ;
    buf_clk cell_4819 ( .C (clk), .D (signal_7364), .Q (signal_7365) ) ;
    buf_clk cell_4835 ( .C (clk), .D (signal_7380), .Q (signal_7381) ) ;
    buf_clk cell_4851 ( .C (clk), .D (signal_7396), .Q (signal_7397) ) ;
    buf_clk cell_4867 ( .C (clk), .D (signal_7412), .Q (signal_7413) ) ;
    buf_clk cell_4883 ( .C (clk), .D (signal_7428), .Q (signal_7429) ) ;
    buf_clk cell_4899 ( .C (clk), .D (signal_7444), .Q (signal_7445) ) ;
    buf_clk cell_4915 ( .C (clk), .D (signal_7460), .Q (signal_7461) ) ;
    buf_clk cell_4931 ( .C (clk), .D (signal_7476), .Q (signal_7477) ) ;
    buf_clk cell_4947 ( .C (clk), .D (signal_7492), .Q (signal_7493) ) ;
    buf_clk cell_4963 ( .C (clk), .D (signal_7508), .Q (signal_7509) ) ;
    buf_clk cell_4979 ( .C (clk), .D (signal_7524), .Q (signal_7525) ) ;
    buf_clk cell_4995 ( .C (clk), .D (signal_7540), .Q (signal_7541) ) ;
    buf_clk cell_5011 ( .C (clk), .D (signal_7556), .Q (signal_7557) ) ;
    buf_clk cell_5027 ( .C (clk), .D (signal_7572), .Q (signal_7573) ) ;
    buf_clk cell_5043 ( .C (clk), .D (signal_7588), .Q (signal_7589) ) ;
    buf_clk cell_5059 ( .C (clk), .D (signal_7604), .Q (signal_7605) ) ;
    buf_clk cell_5075 ( .C (clk), .D (signal_7620), .Q (signal_7621) ) ;
    buf_clk cell_5091 ( .C (clk), .D (signal_7636), .Q (signal_7637) ) ;
    buf_clk cell_5107 ( .C (clk), .D (signal_7652), .Q (signal_7653) ) ;
    buf_clk cell_5123 ( .C (clk), .D (signal_7668), .Q (signal_7669) ) ;
    buf_clk cell_5139 ( .C (clk), .D (signal_7684), .Q (signal_7685) ) ;
    buf_clk cell_5155 ( .C (clk), .D (signal_7700), .Q (signal_7701) ) ;
    buf_clk cell_5171 ( .C (clk), .D (signal_7716), .Q (signal_7717) ) ;
    buf_clk cell_5187 ( .C (clk), .D (signal_7732), .Q (signal_7733) ) ;
    buf_clk cell_5203 ( .C (clk), .D (signal_7748), .Q (signal_7749) ) ;
    buf_clk cell_5219 ( .C (clk), .D (signal_7764), .Q (signal_7765) ) ;
    buf_clk cell_5235 ( .C (clk), .D (signal_7780), .Q (signal_7781) ) ;
    buf_clk cell_5251 ( .C (clk), .D (signal_7796), .Q (signal_7797) ) ;
    buf_clk cell_5267 ( .C (clk), .D (signal_7812), .Q (signal_7813) ) ;
    buf_clk cell_5283 ( .C (clk), .D (signal_7828), .Q (signal_7829) ) ;
    buf_clk cell_5299 ( .C (clk), .D (signal_7844), .Q (signal_7845) ) ;
    buf_clk cell_5315 ( .C (clk), .D (signal_7860), .Q (signal_7861) ) ;
    buf_clk cell_5331 ( .C (clk), .D (signal_7876), .Q (signal_7877) ) ;
    buf_clk cell_5347 ( .C (clk), .D (signal_7892), .Q (signal_7893) ) ;
    buf_clk cell_5363 ( .C (clk), .D (signal_7908), .Q (signal_7909) ) ;
    buf_clk cell_5379 ( .C (clk), .D (signal_7924), .Q (signal_7925) ) ;
    buf_clk cell_5395 ( .C (clk), .D (signal_7940), .Q (signal_7941) ) ;
    buf_clk cell_5411 ( .C (clk), .D (signal_7956), .Q (signal_7957) ) ;
    buf_clk cell_5427 ( .C (clk), .D (signal_7972), .Q (signal_7973) ) ;
    buf_clk cell_5443 ( .C (clk), .D (signal_7988), .Q (signal_7989) ) ;
    buf_clk cell_5459 ( .C (clk), .D (signal_8004), .Q (signal_8005) ) ;
    buf_clk cell_5475 ( .C (clk), .D (signal_8020), .Q (signal_8021) ) ;
    buf_clk cell_5491 ( .C (clk), .D (signal_8036), .Q (signal_8037) ) ;
    buf_clk cell_5507 ( .C (clk), .D (signal_8052), .Q (signal_8053) ) ;
    buf_clk cell_5523 ( .C (clk), .D (signal_8068), .Q (signal_8069) ) ;
    buf_clk cell_5539 ( .C (clk), .D (signal_8084), .Q (signal_8085) ) ;
    buf_clk cell_5555 ( .C (clk), .D (signal_8100), .Q (signal_8101) ) ;
    buf_clk cell_5571 ( .C (clk), .D (signal_8116), .Q (signal_8117) ) ;
    buf_clk cell_5587 ( .C (clk), .D (signal_8132), .Q (signal_8133) ) ;
    buf_clk cell_5603 ( .C (clk), .D (signal_8148), .Q (signal_8149) ) ;
    buf_clk cell_5619 ( .C (clk), .D (signal_8164), .Q (signal_8165) ) ;
    buf_clk cell_5635 ( .C (clk), .D (signal_8180), .Q (signal_8181) ) ;
    buf_clk cell_5651 ( .C (clk), .D (signal_8196), .Q (signal_8197) ) ;
    buf_clk cell_5667 ( .C (clk), .D (signal_8212), .Q (signal_8213) ) ;
    buf_clk cell_5683 ( .C (clk), .D (signal_8228), .Q (signal_8229) ) ;
    buf_clk cell_5699 ( .C (clk), .D (signal_8244), .Q (signal_8245) ) ;
    buf_clk cell_5715 ( .C (clk), .D (signal_8260), .Q (signal_8261) ) ;
    buf_clk cell_5731 ( .C (clk), .D (signal_8276), .Q (signal_8277) ) ;
    buf_clk cell_5747 ( .C (clk), .D (signal_8292), .Q (signal_8293) ) ;
    buf_clk cell_5763 ( .C (clk), .D (signal_8308), .Q (signal_8309) ) ;
    buf_clk cell_5779 ( .C (clk), .D (signal_8324), .Q (signal_8325) ) ;
    buf_clk cell_5795 ( .C (clk), .D (signal_8340), .Q (signal_8341) ) ;
    buf_clk cell_5811 ( .C (clk), .D (signal_8356), .Q (signal_8357) ) ;
    buf_clk cell_5827 ( .C (clk), .D (signal_8372), .Q (signal_8373) ) ;
    buf_clk cell_5843 ( .C (clk), .D (signal_8388), .Q (signal_8389) ) ;
    buf_clk cell_5859 ( .C (clk), .D (signal_8404), .Q (signal_8405) ) ;
    buf_clk cell_5875 ( .C (clk), .D (signal_8420), .Q (signal_8421) ) ;
    buf_clk cell_5891 ( .C (clk), .D (signal_8436), .Q (signal_8437) ) ;
    buf_clk cell_5907 ( .C (clk), .D (signal_8452), .Q (signal_8453) ) ;
    buf_clk cell_5923 ( .C (clk), .D (signal_8468), .Q (signal_8469) ) ;
    buf_clk cell_5939 ( .C (clk), .D (signal_8484), .Q (signal_8485) ) ;
    buf_clk cell_5955 ( .C (clk), .D (signal_8500), .Q (signal_8501) ) ;
    buf_clk cell_5971 ( .C (clk), .D (signal_8516), .Q (signal_8517) ) ;
    buf_clk cell_5987 ( .C (clk), .D (signal_8532), .Q (signal_8533) ) ;
    buf_clk cell_6003 ( .C (clk), .D (signal_8548), .Q (signal_8549) ) ;
    buf_clk cell_6019 ( .C (clk), .D (signal_8564), .Q (signal_8565) ) ;
    buf_clk cell_6035 ( .C (clk), .D (signal_8580), .Q (signal_8581) ) ;
    buf_clk cell_6051 ( .C (clk), .D (signal_8596), .Q (signal_8597) ) ;
    buf_clk cell_6067 ( .C (clk), .D (signal_8612), .Q (signal_8613) ) ;
    buf_clk cell_6083 ( .C (clk), .D (signal_8628), .Q (signal_8629) ) ;
    buf_clk cell_6099 ( .C (clk), .D (signal_8644), .Q (signal_8645) ) ;
    buf_clk cell_6115 ( .C (clk), .D (signal_8660), .Q (signal_8661) ) ;
    buf_clk cell_6131 ( .C (clk), .D (signal_8676), .Q (signal_8677) ) ;
    buf_clk cell_6147 ( .C (clk), .D (signal_8692), .Q (signal_8693) ) ;
    buf_clk cell_6163 ( .C (clk), .D (signal_8708), .Q (signal_8709) ) ;
    buf_clk cell_6179 ( .C (clk), .D (signal_8724), .Q (signal_8725) ) ;
    buf_clk cell_6195 ( .C (clk), .D (signal_8740), .Q (signal_8741) ) ;
    buf_clk cell_6211 ( .C (clk), .D (signal_8756), .Q (signal_8757) ) ;
    buf_clk cell_6227 ( .C (clk), .D (signal_8772), .Q (signal_8773) ) ;
    buf_clk cell_6243 ( .C (clk), .D (signal_8788), .Q (signal_8789) ) ;
    buf_clk cell_6259 ( .C (clk), .D (signal_8804), .Q (signal_8805) ) ;
    buf_clk cell_6275 ( .C (clk), .D (signal_8820), .Q (signal_8821) ) ;
    buf_clk cell_6291 ( .C (clk), .D (signal_8836), .Q (signal_8837) ) ;
    buf_clk cell_6307 ( .C (clk), .D (signal_8852), .Q (signal_8853) ) ;
    buf_clk cell_6323 ( .C (clk), .D (signal_8868), .Q (signal_8869) ) ;
    buf_clk cell_6339 ( .C (clk), .D (signal_8884), .Q (signal_8885) ) ;
    buf_clk cell_6355 ( .C (clk), .D (signal_8900), .Q (signal_8901) ) ;
    buf_clk cell_6371 ( .C (clk), .D (signal_8916), .Q (signal_8917) ) ;
    buf_clk cell_6387 ( .C (clk), .D (signal_8932), .Q (signal_8933) ) ;
    buf_clk cell_6403 ( .C (clk), .D (signal_8948), .Q (signal_8949) ) ;
    buf_clk cell_6419 ( .C (clk), .D (signal_8964), .Q (signal_8965) ) ;
    buf_clk cell_6435 ( .C (clk), .D (signal_8980), .Q (signal_8981) ) ;
    buf_clk cell_6451 ( .C (clk), .D (signal_8996), .Q (signal_8997) ) ;
    buf_clk cell_6467 ( .C (clk), .D (signal_9012), .Q (signal_9013) ) ;
    buf_clk cell_6483 ( .C (clk), .D (signal_9028), .Q (signal_9029) ) ;
    buf_clk cell_6499 ( .C (clk), .D (signal_9044), .Q (signal_9045) ) ;
    buf_clk cell_6515 ( .C (clk), .D (signal_9060), .Q (signal_9061) ) ;
    buf_clk cell_6531 ( .C (clk), .D (signal_9076), .Q (signal_9077) ) ;
    buf_clk cell_6547 ( .C (clk), .D (signal_9092), .Q (signal_9093) ) ;
    buf_clk cell_6563 ( .C (clk), .D (signal_9108), .Q (signal_9109) ) ;
    buf_clk cell_6579 ( .C (clk), .D (signal_9124), .Q (signal_9125) ) ;
    buf_clk cell_6595 ( .C (clk), .D (signal_9140), .Q (signal_9141) ) ;
    buf_clk cell_6611 ( .C (clk), .D (signal_9156), .Q (signal_9157) ) ;
    buf_clk cell_6627 ( .C (clk), .D (signal_9172), .Q (signal_9173) ) ;
    buf_clk cell_6643 ( .C (clk), .D (signal_9188), .Q (signal_9189) ) ;
    buf_clk cell_6659 ( .C (clk), .D (signal_9204), .Q (signal_9205) ) ;
    buf_clk cell_6675 ( .C (clk), .D (signal_9220), .Q (signal_9221) ) ;
    buf_clk cell_6691 ( .C (clk), .D (signal_9236), .Q (signal_9237) ) ;
    buf_clk cell_6707 ( .C (clk), .D (signal_9252), .Q (signal_9253) ) ;
    buf_clk cell_6723 ( .C (clk), .D (signal_9268), .Q (signal_9269) ) ;
    buf_clk cell_6739 ( .C (clk), .D (signal_9284), .Q (signal_9285) ) ;
    buf_clk cell_6755 ( .C (clk), .D (signal_9300), .Q (signal_9301) ) ;
    buf_clk cell_6771 ( .C (clk), .D (signal_9316), .Q (signal_9317) ) ;
    buf_clk cell_6787 ( .C (clk), .D (signal_9332), .Q (signal_9333) ) ;
    buf_clk cell_6803 ( .C (clk), .D (signal_9348), .Q (signal_9349) ) ;
    buf_clk cell_6819 ( .C (clk), .D (signal_9364), .Q (signal_9365) ) ;
    buf_clk cell_6835 ( .C (clk), .D (signal_9380), .Q (signal_9381) ) ;
    buf_clk cell_6851 ( .C (clk), .D (signal_9396), .Q (signal_9397) ) ;
    buf_clk cell_6867 ( .C (clk), .D (signal_9412), .Q (signal_9413) ) ;
    buf_clk cell_6883 ( .C (clk), .D (signal_9428), .Q (signal_9429) ) ;
    buf_clk cell_6899 ( .C (clk), .D (signal_9444), .Q (signal_9445) ) ;
    buf_clk cell_6915 ( .C (clk), .D (signal_9460), .Q (signal_9461) ) ;
    buf_clk cell_6931 ( .C (clk), .D (signal_9476), .Q (signal_9477) ) ;
    buf_clk cell_6947 ( .C (clk), .D (signal_9492), .Q (signal_9493) ) ;
    buf_clk cell_6963 ( .C (clk), .D (signal_9508), .Q (signal_9509) ) ;
    buf_clk cell_6979 ( .C (clk), .D (signal_9524), .Q (signal_9525) ) ;
    buf_clk cell_6995 ( .C (clk), .D (signal_9540), .Q (signal_9541) ) ;
    buf_clk cell_7011 ( .C (clk), .D (signal_9556), .Q (signal_9557) ) ;
    buf_clk cell_7027 ( .C (clk), .D (signal_9572), .Q (signal_9573) ) ;
    buf_clk cell_7043 ( .C (clk), .D (signal_9588), .Q (signal_9589) ) ;
    buf_clk cell_7059 ( .C (clk), .D (signal_9604), .Q (signal_9605) ) ;
    buf_clk cell_7075 ( .C (clk), .D (signal_9620), .Q (signal_9621) ) ;
    buf_clk cell_7091 ( .C (clk), .D (signal_9636), .Q (signal_9637) ) ;
    buf_clk cell_7107 ( .C (clk), .D (signal_9652), .Q (signal_9653) ) ;
    buf_clk cell_7123 ( .C (clk), .D (signal_9668), .Q (signal_9669) ) ;
    buf_clk cell_7139 ( .C (clk), .D (signal_9684), .Q (signal_9685) ) ;
    buf_clk cell_7155 ( .C (clk), .D (signal_9700), .Q (signal_9701) ) ;
    buf_clk cell_7171 ( .C (clk), .D (signal_9716), .Q (signal_9717) ) ;
    buf_clk cell_7187 ( .C (clk), .D (signal_9732), .Q (signal_9733) ) ;
    buf_clk cell_7203 ( .C (clk), .D (signal_9748), .Q (signal_9749) ) ;
    buf_clk cell_7219 ( .C (clk), .D (signal_9764), .Q (signal_9765) ) ;
    buf_clk cell_7235 ( .C (clk), .D (signal_9780), .Q (signal_9781) ) ;
    buf_clk cell_7251 ( .C (clk), .D (signal_9796), .Q (signal_9797) ) ;
    buf_clk cell_7267 ( .C (clk), .D (signal_9812), .Q (signal_9813) ) ;
    buf_clk cell_7283 ( .C (clk), .D (signal_9828), .Q (signal_9829) ) ;
    buf_clk cell_7299 ( .C (clk), .D (signal_9844), .Q (signal_9845) ) ;
    buf_clk cell_7315 ( .C (clk), .D (signal_9860), .Q (signal_9861) ) ;
    buf_clk cell_7331 ( .C (clk), .D (signal_9876), .Q (signal_9877) ) ;
    buf_clk cell_7347 ( .C (clk), .D (signal_9892), .Q (signal_9893) ) ;
    buf_clk cell_7363 ( .C (clk), .D (signal_9908), .Q (signal_9909) ) ;
    buf_clk cell_7379 ( .C (clk), .D (signal_9924), .Q (signal_9925) ) ;
    buf_clk cell_7395 ( .C (clk), .D (signal_9940), .Q (signal_9941) ) ;
    buf_clk cell_7411 ( .C (clk), .D (signal_9956), .Q (signal_9957) ) ;
    buf_clk cell_7427 ( .C (clk), .D (signal_9972), .Q (signal_9973) ) ;
    buf_clk cell_7443 ( .C (clk), .D (signal_9988), .Q (signal_9989) ) ;
    buf_clk cell_7459 ( .C (clk), .D (signal_10004), .Q (signal_10005) ) ;
    buf_clk cell_7475 ( .C (clk), .D (signal_10020), .Q (signal_10021) ) ;
    buf_clk cell_7491 ( .C (clk), .D (signal_10036), .Q (signal_10037) ) ;
    buf_clk cell_7507 ( .C (clk), .D (signal_10052), .Q (signal_10053) ) ;
    buf_clk cell_7523 ( .C (clk), .D (signal_10068), .Q (signal_10069) ) ;
    buf_clk cell_7539 ( .C (clk), .D (signal_10084), .Q (signal_10085) ) ;
    buf_clk cell_7555 ( .C (clk), .D (signal_10100), .Q (signal_10101) ) ;
    buf_clk cell_7571 ( .C (clk), .D (signal_10116), .Q (signal_10117) ) ;
    buf_clk cell_7587 ( .C (clk), .D (signal_10132), .Q (signal_10133) ) ;
    buf_clk cell_7603 ( .C (clk), .D (signal_10148), .Q (signal_10149) ) ;
    buf_clk cell_7619 ( .C (clk), .D (signal_10164), .Q (signal_10165) ) ;
    buf_clk cell_7635 ( .C (clk), .D (signal_10180), .Q (signal_10181) ) ;
    buf_clk cell_7651 ( .C (clk), .D (signal_10196), .Q (signal_10197) ) ;
    buf_clk cell_7667 ( .C (clk), .D (signal_10212), .Q (signal_10213) ) ;
    buf_clk cell_7683 ( .C (clk), .D (signal_10228), .Q (signal_10229) ) ;
    buf_clk cell_7699 ( .C (clk), .D (signal_10244), .Q (signal_10245) ) ;
    buf_clk cell_7715 ( .C (clk), .D (signal_10260), .Q (signal_10261) ) ;
    buf_clk cell_7731 ( .C (clk), .D (signal_10276), .Q (signal_10277) ) ;
    buf_clk cell_7747 ( .C (clk), .D (signal_10292), .Q (signal_10293) ) ;
    buf_clk cell_7763 ( .C (clk), .D (signal_10308), .Q (signal_10309) ) ;
    buf_clk cell_7779 ( .C (clk), .D (signal_10324), .Q (signal_10325) ) ;
    buf_clk cell_7795 ( .C (clk), .D (signal_10340), .Q (signal_10341) ) ;
    buf_clk cell_7811 ( .C (clk), .D (signal_10356), .Q (signal_10357) ) ;
    buf_clk cell_7827 ( .C (clk), .D (signal_10372), .Q (signal_10373) ) ;
    buf_clk cell_7843 ( .C (clk), .D (signal_10388), .Q (signal_10389) ) ;
    buf_clk cell_7859 ( .C (clk), .D (signal_10404), .Q (signal_10405) ) ;
    buf_clk cell_7875 ( .C (clk), .D (signal_10420), .Q (signal_10421) ) ;
    buf_clk cell_7891 ( .C (clk), .D (signal_10436), .Q (signal_10437) ) ;
    buf_clk cell_7907 ( .C (clk), .D (signal_10452), .Q (signal_10453) ) ;
    buf_clk cell_7923 ( .C (clk), .D (signal_10468), .Q (signal_10469) ) ;
    buf_clk cell_7939 ( .C (clk), .D (signal_10484), .Q (signal_10485) ) ;
    buf_clk cell_7955 ( .C (clk), .D (signal_10500), .Q (signal_10501) ) ;
    buf_clk cell_7971 ( .C (clk), .D (signal_10516), .Q (signal_10517) ) ;
    buf_clk cell_7987 ( .C (clk), .D (signal_10532), .Q (signal_10533) ) ;
    buf_clk cell_8003 ( .C (clk), .D (signal_10548), .Q (signal_10549) ) ;
    buf_clk cell_8019 ( .C (clk), .D (signal_10564), .Q (signal_10565) ) ;
    buf_clk cell_8035 ( .C (clk), .D (signal_10580), .Q (signal_10581) ) ;
    buf_clk cell_8051 ( .C (clk), .D (signal_10596), .Q (signal_10597) ) ;
    buf_clk cell_8067 ( .C (clk), .D (signal_10612), .Q (signal_10613) ) ;
    buf_clk cell_8083 ( .C (clk), .D (signal_10628), .Q (signal_10629) ) ;
    buf_clk cell_8099 ( .C (clk), .D (signal_10644), .Q (signal_10645) ) ;
    buf_clk cell_8115 ( .C (clk), .D (signal_10660), .Q (signal_10661) ) ;
    buf_clk cell_8131 ( .C (clk), .D (signal_10676), .Q (signal_10677) ) ;
    buf_clk cell_8147 ( .C (clk), .D (signal_10692), .Q (signal_10693) ) ;
    buf_clk cell_8163 ( .C (clk), .D (signal_10708), .Q (signal_10709) ) ;
    buf_clk cell_8179 ( .C (clk), .D (signal_10724), .Q (signal_10725) ) ;
    buf_clk cell_8195 ( .C (clk), .D (signal_10740), .Q (signal_10741) ) ;
    buf_clk cell_8211 ( .C (clk), .D (signal_10756), .Q (signal_10757) ) ;
    buf_clk cell_8227 ( .C (clk), .D (signal_10772), .Q (signal_10773) ) ;
    buf_clk cell_8243 ( .C (clk), .D (signal_10788), .Q (signal_10789) ) ;
    buf_clk cell_8259 ( .C (clk), .D (signal_10804), .Q (signal_10805) ) ;
    buf_clk cell_8275 ( .C (clk), .D (signal_10820), .Q (signal_10821) ) ;
    buf_clk cell_8291 ( .C (clk), .D (signal_10836), .Q (signal_10837) ) ;
    buf_clk cell_8307 ( .C (clk), .D (signal_10852), .Q (signal_10853) ) ;
    buf_clk cell_8323 ( .C (clk), .D (signal_10868), .Q (signal_10869) ) ;
    buf_clk cell_8339 ( .C (clk), .D (signal_10884), .Q (signal_10885) ) ;
    buf_clk cell_8355 ( .C (clk), .D (signal_10900), .Q (signal_10901) ) ;
    buf_clk cell_8371 ( .C (clk), .D (signal_10916), .Q (signal_10917) ) ;
    buf_clk cell_8387 ( .C (clk), .D (signal_10932), .Q (signal_10933) ) ;
    buf_clk cell_8403 ( .C (clk), .D (signal_10948), .Q (signal_10949) ) ;
    buf_clk cell_8419 ( .C (clk), .D (signal_10964), .Q (signal_10965) ) ;
    buf_clk cell_8435 ( .C (clk), .D (signal_10980), .Q (signal_10981) ) ;
    buf_clk cell_8451 ( .C (clk), .D (signal_10996), .Q (signal_10997) ) ;
    buf_clk cell_8467 ( .C (clk), .D (signal_11012), .Q (signal_11013) ) ;
    buf_clk cell_8483 ( .C (clk), .D (signal_11028), .Q (signal_11029) ) ;
    buf_clk cell_8499 ( .C (clk), .D (signal_11044), .Q (signal_11045) ) ;
    buf_clk cell_8515 ( .C (clk), .D (signal_11060), .Q (signal_11061) ) ;
    buf_clk cell_8531 ( .C (clk), .D (signal_11076), .Q (signal_11077) ) ;
    buf_clk cell_8547 ( .C (clk), .D (signal_11092), .Q (signal_11093) ) ;
    buf_clk cell_8563 ( .C (clk), .D (signal_11108), .Q (signal_11109) ) ;
    buf_clk cell_8579 ( .C (clk), .D (signal_11124), .Q (signal_11125) ) ;
    buf_clk cell_8595 ( .C (clk), .D (signal_11140), .Q (signal_11141) ) ;
    buf_clk cell_8611 ( .C (clk), .D (signal_11156), .Q (signal_11157) ) ;
    buf_clk cell_8627 ( .C (clk), .D (signal_11172), .Q (signal_11173) ) ;
    buf_clk cell_8643 ( .C (clk), .D (signal_11188), .Q (signal_11189) ) ;
    buf_clk cell_8659 ( .C (clk), .D (signal_11204), .Q (signal_11205) ) ;
    buf_clk cell_8675 ( .C (clk), .D (signal_11220), .Q (signal_11221) ) ;
    buf_clk cell_8691 ( .C (clk), .D (signal_11236), .Q (signal_11237) ) ;
    buf_clk cell_8707 ( .C (clk), .D (signal_11252), .Q (signal_11253) ) ;
    buf_clk cell_8723 ( .C (clk), .D (signal_11268), .Q (signal_11269) ) ;
    buf_clk cell_8739 ( .C (clk), .D (signal_11284), .Q (signal_11285) ) ;
    buf_clk cell_8755 ( .C (clk), .D (signal_11300), .Q (signal_11301) ) ;
    buf_clk cell_8771 ( .C (clk), .D (signal_11316), .Q (signal_11317) ) ;
    buf_clk cell_8787 ( .C (clk), .D (signal_11332), .Q (signal_11333) ) ;
    buf_clk cell_8803 ( .C (clk), .D (signal_11348), .Q (signal_11349) ) ;
    buf_clk cell_8819 ( .C (clk), .D (signal_11364), .Q (signal_11365) ) ;
    buf_clk cell_8835 ( .C (clk), .D (signal_11380), .Q (signal_11381) ) ;
    buf_clk cell_8851 ( .C (clk), .D (signal_11396), .Q (signal_11397) ) ;
    buf_clk cell_8867 ( .C (clk), .D (signal_11412), .Q (signal_11413) ) ;
    buf_clk cell_8883 ( .C (clk), .D (signal_11428), .Q (signal_11429) ) ;
    buf_clk cell_8899 ( .C (clk), .D (signal_11444), .Q (signal_11445) ) ;
    buf_clk cell_8915 ( .C (clk), .D (signal_11460), .Q (signal_11461) ) ;
    buf_clk cell_8931 ( .C (clk), .D (signal_11476), .Q (signal_11477) ) ;
    buf_clk cell_8947 ( .C (clk), .D (signal_11492), .Q (signal_11493) ) ;
    buf_clk cell_8963 ( .C (clk), .D (signal_11508), .Q (signal_11509) ) ;
    buf_clk cell_8979 ( .C (clk), .D (signal_11524), .Q (signal_11525) ) ;
    buf_clk cell_8995 ( .C (clk), .D (signal_11540), .Q (signal_11541) ) ;
    buf_clk cell_9011 ( .C (clk), .D (signal_11556), .Q (signal_11557) ) ;
    buf_clk cell_9027 ( .C (clk), .D (signal_11572), .Q (signal_11573) ) ;
    buf_clk cell_9043 ( .C (clk), .D (signal_11588), .Q (signal_11589) ) ;
    buf_clk cell_9059 ( .C (clk), .D (signal_11604), .Q (signal_11605) ) ;
    buf_clk cell_9075 ( .C (clk), .D (signal_11620), .Q (signal_11621) ) ;
    buf_clk cell_9091 ( .C (clk), .D (signal_11636), .Q (signal_11637) ) ;
    buf_clk cell_9107 ( .C (clk), .D (signal_11652), .Q (signal_11653) ) ;
    buf_clk cell_9123 ( .C (clk), .D (signal_11668), .Q (signal_11669) ) ;
    buf_clk cell_9139 ( .C (clk), .D (signal_11684), .Q (signal_11685) ) ;
    buf_clk cell_9155 ( .C (clk), .D (signal_11700), .Q (signal_11701) ) ;
    buf_clk cell_9171 ( .C (clk), .D (signal_11716), .Q (signal_11717) ) ;
    buf_clk cell_9187 ( .C (clk), .D (signal_11732), .Q (signal_11733) ) ;
    buf_clk cell_9203 ( .C (clk), .D (signal_11748), .Q (signal_11749) ) ;
    buf_clk cell_9219 ( .C (clk), .D (signal_11764), .Q (signal_11765) ) ;
    buf_clk cell_9235 ( .C (clk), .D (signal_11780), .Q (signal_11781) ) ;
    buf_clk cell_9251 ( .C (clk), .D (signal_11796), .Q (signal_11797) ) ;
    buf_clk cell_9267 ( .C (clk), .D (signal_11812), .Q (signal_11813) ) ;
    buf_clk cell_9283 ( .C (clk), .D (signal_11828), .Q (signal_11829) ) ;
    buf_clk cell_9299 ( .C (clk), .D (signal_11844), .Q (signal_11845) ) ;
    buf_clk cell_9315 ( .C (clk), .D (signal_11860), .Q (signal_11861) ) ;
    buf_clk cell_9331 ( .C (clk), .D (signal_11876), .Q (signal_11877) ) ;
    buf_clk cell_9347 ( .C (clk), .D (signal_11892), .Q (signal_11893) ) ;
    buf_clk cell_9363 ( .C (clk), .D (signal_11908), .Q (signal_11909) ) ;
    buf_clk cell_9379 ( .C (clk), .D (signal_11924), .Q (signal_11925) ) ;
    buf_clk cell_9395 ( .C (clk), .D (signal_11940), .Q (signal_11941) ) ;
    buf_clk cell_9411 ( .C (clk), .D (signal_11956), .Q (signal_11957) ) ;
    buf_clk cell_9427 ( .C (clk), .D (signal_11972), .Q (signal_11973) ) ;
    buf_clk cell_9443 ( .C (clk), .D (signal_11988), .Q (signal_11989) ) ;
    buf_clk cell_9459 ( .C (clk), .D (signal_12004), .Q (signal_12005) ) ;
    buf_clk cell_9475 ( .C (clk), .D (signal_12020), .Q (signal_12021) ) ;
    buf_clk cell_9491 ( .C (clk), .D (signal_12036), .Q (signal_12037) ) ;
    buf_clk cell_9507 ( .C (clk), .D (signal_12052), .Q (signal_12053) ) ;
    buf_clk cell_9523 ( .C (clk), .D (signal_12068), .Q (signal_12069) ) ;
    buf_clk cell_9539 ( .C (clk), .D (signal_12084), .Q (signal_12085) ) ;
    buf_clk cell_9555 ( .C (clk), .D (signal_12100), .Q (signal_12101) ) ;
    buf_clk cell_9571 ( .C (clk), .D (signal_12116), .Q (signal_12117) ) ;
    buf_clk cell_9587 ( .C (clk), .D (signal_12132), .Q (signal_12133) ) ;
    buf_clk cell_9603 ( .C (clk), .D (signal_12148), .Q (signal_12149) ) ;
    buf_clk cell_9619 ( .C (clk), .D (signal_12164), .Q (signal_12165) ) ;
    buf_clk cell_9635 ( .C (clk), .D (signal_12180), .Q (signal_12181) ) ;
    buf_clk cell_9651 ( .C (clk), .D (signal_12196), .Q (signal_12197) ) ;
    buf_clk cell_9667 ( .C (clk), .D (signal_12212), .Q (signal_12213) ) ;
    buf_clk cell_9683 ( .C (clk), .D (signal_12228), .Q (signal_12229) ) ;
    buf_clk cell_9699 ( .C (clk), .D (signal_12244), .Q (signal_12245) ) ;
    buf_clk cell_9715 ( .C (clk), .D (signal_12260), .Q (signal_12261) ) ;
    buf_clk cell_9731 ( .C (clk), .D (signal_12276), .Q (signal_12277) ) ;
    buf_clk cell_9747 ( .C (clk), .D (signal_12292), .Q (signal_12293) ) ;
    buf_clk cell_9763 ( .C (clk), .D (signal_12308), .Q (signal_12309) ) ;
    buf_clk cell_9779 ( .C (clk), .D (signal_12324), .Q (signal_12325) ) ;
    buf_clk cell_9795 ( .C (clk), .D (signal_12340), .Q (signal_12341) ) ;
    buf_clk cell_9811 ( .C (clk), .D (signal_12356), .Q (signal_12357) ) ;
    buf_clk cell_9827 ( .C (clk), .D (signal_12372), .Q (signal_12373) ) ;
    buf_clk cell_9843 ( .C (clk), .D (signal_12388), .Q (signal_12389) ) ;
    buf_clk cell_9859 ( .C (clk), .D (signal_12404), .Q (signal_12405) ) ;
    buf_clk cell_9875 ( .C (clk), .D (signal_12420), .Q (signal_12421) ) ;
    buf_clk cell_9891 ( .C (clk), .D (signal_12436), .Q (signal_12437) ) ;
    buf_clk cell_9907 ( .C (clk), .D (signal_12452), .Q (signal_12453) ) ;
    buf_clk cell_9923 ( .C (clk), .D (signal_12468), .Q (signal_12469) ) ;
    buf_clk cell_9939 ( .C (clk), .D (signal_12484), .Q (signal_12485) ) ;
    buf_clk cell_9955 ( .C (clk), .D (signal_12500), .Q (signal_12501) ) ;
    buf_clk cell_9971 ( .C (clk), .D (signal_12516), .Q (signal_12517) ) ;
    buf_clk cell_9987 ( .C (clk), .D (signal_12532), .Q (signal_12533) ) ;
    buf_clk cell_10003 ( .C (clk), .D (signal_12548), .Q (signal_12549) ) ;
    buf_clk cell_10019 ( .C (clk), .D (signal_12564), .Q (signal_12565) ) ;
    buf_clk cell_10035 ( .C (clk), .D (signal_12580), .Q (signal_12581) ) ;
    buf_clk cell_10051 ( .C (clk), .D (signal_12596), .Q (signal_12597) ) ;
    buf_clk cell_10067 ( .C (clk), .D (signal_12612), .Q (signal_12613) ) ;
    buf_clk cell_10083 ( .C (clk), .D (signal_12628), .Q (signal_12629) ) ;
    buf_clk cell_10099 ( .C (clk), .D (signal_12644), .Q (signal_12645) ) ;
    buf_clk cell_10115 ( .C (clk), .D (signal_12660), .Q (signal_12661) ) ;
    buf_clk cell_10131 ( .C (clk), .D (signal_12676), .Q (signal_12677) ) ;
    buf_clk cell_10147 ( .C (clk), .D (signal_12692), .Q (signal_12693) ) ;
    buf_clk cell_10163 ( .C (clk), .D (signal_12708), .Q (signal_12709) ) ;
    buf_clk cell_10179 ( .C (clk), .D (signal_12724), .Q (signal_12725) ) ;
    buf_clk cell_10195 ( .C (clk), .D (signal_12740), .Q (signal_12741) ) ;
    buf_clk cell_10211 ( .C (clk), .D (signal_12756), .Q (signal_12757) ) ;
    buf_clk cell_10227 ( .C (clk), .D (signal_12772), .Q (signal_12773) ) ;
    buf_clk cell_10243 ( .C (clk), .D (signal_12788), .Q (signal_12789) ) ;
    buf_clk cell_10259 ( .C (clk), .D (signal_12804), .Q (signal_12805) ) ;
    buf_clk cell_10275 ( .C (clk), .D (signal_12820), .Q (signal_12821) ) ;
    buf_clk cell_10291 ( .C (clk), .D (signal_12836), .Q (signal_12837) ) ;
    buf_clk cell_10307 ( .C (clk), .D (signal_12852), .Q (signal_12853) ) ;
    buf_clk cell_10323 ( .C (clk), .D (signal_12868), .Q (signal_12869) ) ;
    buf_clk cell_10339 ( .C (clk), .D (signal_12884), .Q (signal_12885) ) ;
    buf_clk cell_10355 ( .C (clk), .D (signal_12900), .Q (signal_12901) ) ;
    buf_clk cell_10371 ( .C (clk), .D (signal_12916), .Q (signal_12917) ) ;
    buf_clk cell_10387 ( .C (clk), .D (signal_12932), .Q (signal_12933) ) ;
    buf_clk cell_10403 ( .C (clk), .D (signal_12948), .Q (signal_12949) ) ;
    buf_clk cell_10419 ( .C (clk), .D (signal_12964), .Q (signal_12965) ) ;
    buf_clk cell_10435 ( .C (clk), .D (signal_12980), .Q (signal_12981) ) ;
    buf_clk cell_10451 ( .C (clk), .D (signal_12996), .Q (signal_12997) ) ;
    buf_clk cell_10467 ( .C (clk), .D (signal_13012), .Q (signal_13013) ) ;
    buf_clk cell_10483 ( .C (clk), .D (signal_13028), .Q (signal_13029) ) ;
    buf_clk cell_10499 ( .C (clk), .D (signal_13044), .Q (signal_13045) ) ;
    buf_clk cell_10515 ( .C (clk), .D (signal_13060), .Q (signal_13061) ) ;
    buf_clk cell_10531 ( .C (clk), .D (signal_13076), .Q (signal_13077) ) ;
    buf_clk cell_10547 ( .C (clk), .D (signal_13092), .Q (signal_13093) ) ;
    buf_clk cell_10563 ( .C (clk), .D (signal_13108), .Q (signal_13109) ) ;
    buf_clk cell_10579 ( .C (clk), .D (signal_13124), .Q (signal_13125) ) ;
    buf_clk cell_10595 ( .C (clk), .D (signal_13140), .Q (signal_13141) ) ;
    buf_clk cell_10611 ( .C (clk), .D (signal_13156), .Q (signal_13157) ) ;
    buf_clk cell_10627 ( .C (clk), .D (signal_13172), .Q (signal_13173) ) ;
    buf_clk cell_10643 ( .C (clk), .D (signal_13188), .Q (signal_13189) ) ;
    buf_clk cell_10659 ( .C (clk), .D (signal_13204), .Q (signal_13205) ) ;
    buf_clk cell_10675 ( .C (clk), .D (signal_13220), .Q (signal_13221) ) ;
    buf_clk cell_10691 ( .C (clk), .D (signal_13236), .Q (signal_13237) ) ;
    buf_clk cell_10707 ( .C (clk), .D (signal_13252), .Q (signal_13253) ) ;
    buf_clk cell_10723 ( .C (clk), .D (signal_13268), .Q (signal_13269) ) ;
    buf_clk cell_10739 ( .C (clk), .D (signal_13284), .Q (signal_13285) ) ;
    buf_clk cell_10755 ( .C (clk), .D (signal_13300), .Q (signal_13301) ) ;
    buf_clk cell_10771 ( .C (clk), .D (signal_13316), .Q (signal_13317) ) ;
    buf_clk cell_10787 ( .C (clk), .D (signal_13332), .Q (signal_13333) ) ;
    buf_clk cell_10803 ( .C (clk), .D (signal_13348), .Q (signal_13349) ) ;
    buf_clk cell_10819 ( .C (clk), .D (signal_13364), .Q (signal_13365) ) ;
    buf_clk cell_10835 ( .C (clk), .D (signal_13380), .Q (signal_13381) ) ;
    buf_clk cell_10851 ( .C (clk), .D (signal_13396), .Q (signal_13397) ) ;
    buf_clk cell_10867 ( .C (clk), .D (signal_13412), .Q (signal_13413) ) ;
    buf_clk cell_10883 ( .C (clk), .D (signal_13428), .Q (signal_13429) ) ;
    buf_clk cell_10899 ( .C (clk), .D (signal_13444), .Q (signal_13445) ) ;
    buf_clk cell_10915 ( .C (clk), .D (signal_13460), .Q (signal_13461) ) ;
    buf_clk cell_10931 ( .C (clk), .D (signal_13476), .Q (signal_13477) ) ;
    buf_clk cell_10947 ( .C (clk), .D (signal_13492), .Q (signal_13493) ) ;
    buf_clk cell_10963 ( .C (clk), .D (signal_13508), .Q (signal_13509) ) ;
    buf_clk cell_10979 ( .C (clk), .D (signal_13524), .Q (signal_13525) ) ;
    buf_clk cell_10995 ( .C (clk), .D (signal_13540), .Q (signal_13541) ) ;
    buf_clk cell_11011 ( .C (clk), .D (signal_13556), .Q (signal_13557) ) ;
    buf_clk cell_11027 ( .C (clk), .D (signal_13572), .Q (signal_13573) ) ;
    buf_clk cell_11043 ( .C (clk), .D (signal_13588), .Q (signal_13589) ) ;
    buf_clk cell_11059 ( .C (clk), .D (signal_13604), .Q (signal_13605) ) ;
    buf_clk cell_11075 ( .C (clk), .D (signal_13620), .Q (signal_13621) ) ;
    buf_clk cell_11091 ( .C (clk), .D (signal_13636), .Q (signal_13637) ) ;
    buf_clk cell_11107 ( .C (clk), .D (signal_13652), .Q (signal_13653) ) ;
    buf_clk cell_11123 ( .C (clk), .D (signal_13668), .Q (signal_13669) ) ;
    buf_clk cell_11139 ( .C (clk), .D (signal_13684), .Q (signal_13685) ) ;
    buf_clk cell_11155 ( .C (clk), .D (signal_13700), .Q (signal_13701) ) ;
    buf_clk cell_11171 ( .C (clk), .D (signal_13716), .Q (signal_13717) ) ;
    buf_clk cell_11187 ( .C (clk), .D (signal_13732), .Q (signal_13733) ) ;
    buf_clk cell_11203 ( .C (clk), .D (signal_13748), .Q (signal_13749) ) ;
    buf_clk cell_11219 ( .C (clk), .D (signal_13764), .Q (signal_13765) ) ;
    buf_clk cell_11235 ( .C (clk), .D (signal_13780), .Q (signal_13781) ) ;
    buf_clk cell_11251 ( .C (clk), .D (signal_13796), .Q (signal_13797) ) ;
    buf_clk cell_11267 ( .C (clk), .D (signal_13812), .Q (signal_13813) ) ;
    buf_clk cell_11283 ( .C (clk), .D (signal_13828), .Q (signal_13829) ) ;
    buf_clk cell_11299 ( .C (clk), .D (signal_13844), .Q (signal_13845) ) ;
    buf_clk cell_11315 ( .C (clk), .D (signal_13860), .Q (signal_13861) ) ;
    buf_clk cell_11331 ( .C (clk), .D (signal_13876), .Q (signal_13877) ) ;
    buf_clk cell_11347 ( .C (clk), .D (signal_13892), .Q (signal_13893) ) ;
    buf_clk cell_11363 ( .C (clk), .D (signal_13908), .Q (signal_13909) ) ;
    buf_clk cell_11379 ( .C (clk), .D (signal_13924), .Q (signal_13925) ) ;
    buf_clk cell_11395 ( .C (clk), .D (signal_13940), .Q (signal_13941) ) ;
    buf_clk cell_11411 ( .C (clk), .D (signal_13956), .Q (signal_13957) ) ;
    buf_clk cell_11427 ( .C (clk), .D (signal_13972), .Q (signal_13973) ) ;
    buf_clk cell_11443 ( .C (clk), .D (signal_13988), .Q (signal_13989) ) ;
    buf_clk cell_11459 ( .C (clk), .D (signal_14004), .Q (signal_14005) ) ;
    buf_clk cell_11475 ( .C (clk), .D (signal_14020), .Q (signal_14021) ) ;
    buf_clk cell_11491 ( .C (clk), .D (signal_14036), .Q (signal_14037) ) ;
    buf_clk cell_11507 ( .C (clk), .D (signal_14052), .Q (signal_14053) ) ;
    buf_clk cell_11523 ( .C (clk), .D (signal_14068), .Q (signal_14069) ) ;
    buf_clk cell_11539 ( .C (clk), .D (signal_14084), .Q (signal_14085) ) ;
    buf_clk cell_11555 ( .C (clk), .D (signal_14100), .Q (signal_14101) ) ;
    buf_clk cell_11571 ( .C (clk), .D (signal_14116), .Q (signal_14117) ) ;
    buf_clk cell_11587 ( .C (clk), .D (signal_14132), .Q (signal_14133) ) ;
    buf_clk cell_11603 ( .C (clk), .D (signal_14148), .Q (signal_14149) ) ;
    buf_clk cell_11619 ( .C (clk), .D (signal_14164), .Q (signal_14165) ) ;
    buf_clk cell_11635 ( .C (clk), .D (signal_14180), .Q (signal_14181) ) ;
    buf_clk cell_11651 ( .C (clk), .D (signal_14196), .Q (signal_14197) ) ;
    buf_clk cell_11667 ( .C (clk), .D (signal_14212), .Q (signal_14213) ) ;
    buf_clk cell_11683 ( .C (clk), .D (signal_14228), .Q (signal_14229) ) ;
    buf_clk cell_11699 ( .C (clk), .D (signal_14244), .Q (signal_14245) ) ;
    buf_clk cell_11715 ( .C (clk), .D (signal_14260), .Q (signal_14261) ) ;
    buf_clk cell_11731 ( .C (clk), .D (signal_14276), .Q (signal_14277) ) ;
    buf_clk cell_11747 ( .C (clk), .D (signal_14292), .Q (signal_14293) ) ;
    buf_clk cell_11763 ( .C (clk), .D (signal_14308), .Q (signal_14309) ) ;
    buf_clk cell_11779 ( .C (clk), .D (signal_14324), .Q (signal_14325) ) ;
    buf_clk cell_11795 ( .C (clk), .D (signal_14340), .Q (signal_14341) ) ;
    buf_clk cell_11811 ( .C (clk), .D (signal_14356), .Q (signal_14357) ) ;
    buf_clk cell_11827 ( .C (clk), .D (signal_14372), .Q (signal_14373) ) ;
    buf_clk cell_11843 ( .C (clk), .D (signal_14388), .Q (signal_14389) ) ;
    buf_clk cell_11859 ( .C (clk), .D (signal_14404), .Q (signal_14405) ) ;
    buf_clk cell_11875 ( .C (clk), .D (signal_14420), .Q (signal_14421) ) ;
    buf_clk cell_11891 ( .C (clk), .D (signal_14436), .Q (signal_14437) ) ;
    buf_clk cell_11907 ( .C (clk), .D (signal_14452), .Q (signal_14453) ) ;
    buf_clk cell_11923 ( .C (clk), .D (signal_14468), .Q (signal_14469) ) ;
    buf_clk cell_11939 ( .C (clk), .D (signal_14484), .Q (signal_14485) ) ;
    buf_clk cell_11955 ( .C (clk), .D (signal_14500), .Q (signal_14501) ) ;
    buf_clk cell_11971 ( .C (clk), .D (signal_14516), .Q (signal_14517) ) ;
    buf_clk cell_11987 ( .C (clk), .D (signal_14532), .Q (signal_14533) ) ;
    buf_clk cell_12003 ( .C (clk), .D (signal_14548), .Q (signal_14549) ) ;
    buf_clk cell_12019 ( .C (clk), .D (signal_14564), .Q (signal_14565) ) ;
    buf_clk cell_12035 ( .C (clk), .D (signal_14580), .Q (signal_14581) ) ;
    buf_clk cell_12051 ( .C (clk), .D (signal_14596), .Q (signal_14597) ) ;
    buf_clk cell_12067 ( .C (clk), .D (signal_14612), .Q (signal_14613) ) ;
    buf_clk cell_12083 ( .C (clk), .D (signal_14628), .Q (signal_14629) ) ;
    buf_clk cell_12099 ( .C (clk), .D (signal_14644), .Q (signal_14645) ) ;
    buf_clk cell_12115 ( .C (clk), .D (signal_14660), .Q (signal_14661) ) ;
    buf_clk cell_12131 ( .C (clk), .D (signal_14676), .Q (signal_14677) ) ;
    buf_clk cell_12147 ( .C (clk), .D (signal_14692), .Q (signal_14693) ) ;
    buf_clk cell_12163 ( .C (clk), .D (signal_14708), .Q (signal_14709) ) ;
    buf_clk cell_12179 ( .C (clk), .D (signal_14724), .Q (signal_14725) ) ;
    buf_clk cell_12195 ( .C (clk), .D (signal_14740), .Q (signal_14741) ) ;
    buf_clk cell_12211 ( .C (clk), .D (signal_14756), .Q (signal_14757) ) ;
    buf_clk cell_12227 ( .C (clk), .D (signal_14772), .Q (signal_14773) ) ;
    buf_clk cell_12243 ( .C (clk), .D (signal_14788), .Q (signal_14789) ) ;
    buf_clk cell_12259 ( .C (clk), .D (signal_14804), .Q (signal_14805) ) ;
    buf_clk cell_12275 ( .C (clk), .D (signal_14820), .Q (signal_14821) ) ;
    buf_clk cell_12291 ( .C (clk), .D (signal_14836), .Q (signal_14837) ) ;
    buf_clk cell_12307 ( .C (clk), .D (signal_14852), .Q (signal_14853) ) ;
    buf_clk cell_12323 ( .C (clk), .D (signal_14868), .Q (signal_14869) ) ;
    buf_clk cell_12339 ( .C (clk), .D (signal_14884), .Q (signal_14885) ) ;
    buf_clk cell_12355 ( .C (clk), .D (signal_14900), .Q (signal_14901) ) ;
    buf_clk cell_12371 ( .C (clk), .D (signal_14916), .Q (signal_14917) ) ;
    buf_clk cell_12387 ( .C (clk), .D (signal_14932), .Q (signal_14933) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1904 ( .s ({signal_4734, signal_4732}), .b ({signal_3477, signal_2022}), .a ({signal_3476, signal_2021}), .clk (clk), .r (Fresh[190]), .c ({signal_3699, signal_2172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1905 ( .s ({signal_4734, signal_4732}), .b ({signal_3479, signal_2024}), .a ({signal_3478, signal_2023}), .clk (clk), .r (Fresh[191]), .c ({signal_3700, signal_2173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1906 ( .s ({signal_4734, signal_4732}), .b ({signal_3481, signal_2026}), .a ({signal_3480, signal_2025}), .clk (clk), .r (Fresh[192]), .c ({signal_3701, signal_2174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1907 ( .s ({signal_4734, signal_4732}), .b ({signal_3482, signal_2027}), .a ({signal_4738, signal_4736}), .clk (clk), .r (Fresh[193]), .c ({signal_3702, signal_2175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1908 ( .s ({signal_4734, signal_4732}), .b ({signal_4742, signal_4740}), .a ({signal_3483, signal_2028}), .clk (clk), .r (Fresh[194]), .c ({signal_3703, signal_2176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1909 ( .s ({signal_4734, signal_4732}), .b ({signal_3485, signal_2030}), .a ({signal_3484, signal_2029}), .clk (clk), .r (Fresh[195]), .c ({signal_3704, signal_2177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1910 ( .s ({signal_4734, signal_4732}), .b ({signal_3487, signal_2032}), .a ({signal_3486, signal_2031}), .clk (clk), .r (Fresh[196]), .c ({signal_3705, signal_2178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1911 ( .s ({signal_4734, signal_4732}), .b ({signal_3489, signal_2034}), .a ({signal_3488, signal_2033}), .clk (clk), .r (Fresh[197]), .c ({signal_3706, signal_2179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1912 ( .s ({signal_4734, signal_4732}), .b ({signal_3492, signal_2037}), .a ({signal_3491, signal_2036}), .clk (clk), .r (Fresh[198]), .c ({signal_3707, signal_2180}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1913 ( .s ({signal_4734, signal_4732}), .b ({signal_3493, signal_2038}), .a ({signal_4746, signal_4744}), .clk (clk), .r (Fresh[199]), .c ({signal_3708, signal_2181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1914 ( .s ({signal_4734, signal_4732}), .b ({signal_3494, signal_2039}), .a ({signal_4750, signal_4748}), .clk (clk), .r (Fresh[200]), .c ({signal_3709, signal_2182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1915 ( .s ({signal_4734, signal_4732}), .b ({signal_3496, signal_2041}), .a ({signal_4754, signal_4752}), .clk (clk), .r (Fresh[201]), .c ({signal_3710, signal_2183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1916 ( .s ({signal_4734, signal_4732}), .b ({signal_3498, signal_2043}), .a ({signal_3478, signal_2023}), .clk (clk), .r (Fresh[202]), .c ({signal_3711, signal_2184}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1917 ( .s ({signal_4734, signal_4732}), .b ({signal_3500, signal_2045}), .a ({signal_3499, signal_2044}), .clk (clk), .r (Fresh[203]), .c ({signal_3712, signal_2185}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1918 ( .s ({signal_4734, signal_4732}), .b ({signal_4758, signal_4756}), .a ({signal_3501, signal_2046}), .clk (clk), .r (Fresh[204]), .c ({signal_3713, signal_2186}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1919 ( .s ({signal_4734, signal_4732}), .b ({signal_3503, signal_2048}), .a ({signal_3502, signal_2047}), .clk (clk), .r (Fresh[205]), .c ({signal_3714, signal_2187}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1920 ( .s ({signal_4734, signal_4732}), .b ({signal_3504, signal_2049}), .a ({signal_3483, signal_2028}), .clk (clk), .r (Fresh[206]), .c ({signal_3715, signal_2188}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1921 ( .s ({signal_4734, signal_4732}), .b ({signal_4762, signal_4760}), .a ({signal_3505, signal_2050}), .clk (clk), .r (Fresh[207]), .c ({signal_3716, signal_2189}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1922 ( .s ({signal_4734, signal_4732}), .b ({signal_4766, signal_4764}), .a ({signal_3506, signal_2051}), .clk (clk), .r (Fresh[208]), .c ({signal_3717, signal_2190}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1923 ( .s ({signal_4734, signal_4732}), .b ({signal_3508, signal_2053}), .a ({signal_3507, signal_2052}), .clk (clk), .r (Fresh[209]), .c ({signal_3718, signal_2191}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1924 ( .s ({signal_4734, signal_4732}), .b ({signal_3478, signal_2023}), .a ({signal_3509, signal_2054}), .clk (clk), .r (Fresh[210]), .c ({signal_3719, signal_2192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1925 ( .s ({signal_4734, signal_4732}), .b ({signal_3510, signal_2055}), .a ({signal_4770, signal_4768}), .clk (clk), .r (Fresh[211]), .c ({signal_3720, signal_2193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1926 ( .s ({signal_4734, signal_4732}), .b ({signal_3512, signal_2057}), .a ({signal_3511, signal_2056}), .clk (clk), .r (Fresh[212]), .c ({signal_3721, signal_2194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1927 ( .s ({signal_4734, signal_4732}), .b ({signal_3513, signal_2058}), .a ({signal_3510, signal_2055}), .clk (clk), .r (Fresh[213]), .c ({signal_3722, signal_2195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1928 ( .s ({signal_4734, signal_4732}), .b ({signal_3515, signal_2060}), .a ({signal_3514, signal_2059}), .clk (clk), .r (Fresh[214]), .c ({signal_3723, signal_2196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1929 ( .s ({signal_4734, signal_4732}), .b ({signal_3517, signal_2062}), .a ({signal_3516, signal_2061}), .clk (clk), .r (Fresh[215]), .c ({signal_3724, signal_2197}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1930 ( .s ({signal_4734, signal_4732}), .b ({signal_3518, signal_2063}), .a ({signal_4774, signal_4772}), .clk (clk), .r (Fresh[216]), .c ({signal_3725, signal_2198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1931 ( .s ({signal_4734, signal_4732}), .b ({signal_3519, signal_2064}), .a ({signal_3476, signal_2021}), .clk (clk), .r (Fresh[217]), .c ({signal_3726, signal_2199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1932 ( .s ({signal_4734, signal_4732}), .b ({signal_3521, signal_2066}), .a ({signal_3520, signal_2065}), .clk (clk), .r (Fresh[218]), .c ({signal_3727, signal_2200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1933 ( .s ({signal_4734, signal_4732}), .b ({signal_3523, signal_2068}), .a ({signal_3522, signal_2067}), .clk (clk), .r (Fresh[219]), .c ({signal_3728, signal_2201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1934 ( .s ({signal_4734, signal_4732}), .b ({signal_3525, signal_2070}), .a ({signal_3524, signal_2069}), .clk (clk), .r (Fresh[220]), .c ({signal_3729, signal_2202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1935 ( .s ({signal_4734, signal_4732}), .b ({signal_3527, signal_2072}), .a ({signal_3526, signal_2071}), .clk (clk), .r (Fresh[221]), .c ({signal_3730, signal_2203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1936 ( .s ({signal_4734, signal_4732}), .b ({signal_3529, signal_2074}), .a ({signal_3528, signal_2073}), .clk (clk), .r (Fresh[222]), .c ({signal_3731, signal_2204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1937 ( .s ({signal_4734, signal_4732}), .b ({signal_3531, signal_2076}), .a ({signal_3530, signal_2075}), .clk (clk), .r (Fresh[223]), .c ({signal_3732, signal_2205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1938 ( .s ({signal_4734, signal_4732}), .b ({signal_3533, signal_2078}), .a ({signal_3532, signal_2077}), .clk (clk), .r (Fresh[224]), .c ({signal_3733, signal_2206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1939 ( .s ({signal_4734, signal_4732}), .b ({signal_3506, signal_2051}), .a ({signal_3534, signal_2079}), .clk (clk), .r (Fresh[225]), .c ({signal_3734, signal_2207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1940 ( .s ({signal_4734, signal_4732}), .b ({signal_4778, signal_4776}), .a ({signal_3535, signal_2080}), .clk (clk), .r (Fresh[226]), .c ({signal_3735, signal_2208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1941 ( .s ({signal_4734, signal_4732}), .b ({signal_3478, signal_2023}), .a ({signal_3536, signal_2081}), .clk (clk), .r (Fresh[227]), .c ({signal_3736, signal_2209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1942 ( .s ({signal_4734, signal_4732}), .b ({signal_4750, signal_4748}), .a ({signal_3537, signal_2082}), .clk (clk), .r (Fresh[228]), .c ({signal_3737, signal_2210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1943 ( .s ({signal_4734, signal_4732}), .b ({signal_3538, signal_2083}), .a ({signal_4782, signal_4780}), .clk (clk), .r (Fresh[229]), .c ({signal_3738, signal_2211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1944 ( .s ({signal_4734, signal_4732}), .b ({signal_3540, signal_2085}), .a ({signal_3539, signal_2084}), .clk (clk), .r (Fresh[230]), .c ({signal_3739, signal_2212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1945 ( .s ({signal_4734, signal_4732}), .b ({signal_3526, signal_2071}), .a ({signal_3541, signal_2086}), .clk (clk), .r (Fresh[231]), .c ({signal_3740, signal_2213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1946 ( .s ({signal_4734, signal_4732}), .b ({signal_3529, signal_2074}), .a ({signal_4754, signal_4752}), .clk (clk), .r (Fresh[232]), .c ({signal_3741, signal_2214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1947 ( .s ({signal_4734, signal_4732}), .b ({signal_3542, signal_2087}), .a ({signal_3515, signal_2060}), .clk (clk), .r (Fresh[233]), .c ({signal_3742, signal_2215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1948 ( .s ({signal_4734, signal_4732}), .b ({signal_3544, signal_2089}), .a ({signal_3543, signal_2088}), .clk (clk), .r (Fresh[234]), .c ({signal_3743, signal_2216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1949 ( .s ({signal_4734, signal_4732}), .b ({signal_3546, signal_2091}), .a ({signal_3545, signal_2090}), .clk (clk), .r (Fresh[235]), .c ({signal_3744, signal_2217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1950 ( .s ({signal_4734, signal_4732}), .b ({signal_4786, signal_4784}), .a ({signal_3547, signal_2092}), .clk (clk), .r (Fresh[236]), .c ({signal_3745, signal_2218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1951 ( .s ({signal_4734, signal_4732}), .b ({signal_3549, signal_2094}), .a ({signal_3548, signal_2093}), .clk (clk), .r (Fresh[237]), .c ({signal_3746, signal_2219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1952 ( .s ({signal_4734, signal_4732}), .b ({signal_3551, signal_2096}), .a ({signal_3550, signal_2095}), .clk (clk), .r (Fresh[238]), .c ({signal_3747, signal_2220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1953 ( .s ({signal_4734, signal_4732}), .b ({signal_3512, signal_2057}), .a ({signal_3553, signal_2098}), .clk (clk), .r (Fresh[239]), .c ({signal_3748, signal_2221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1954 ( .s ({signal_4734, signal_4732}), .b ({signal_4790, signal_4788}), .a ({signal_3554, signal_2099}), .clk (clk), .r (Fresh[240]), .c ({signal_3749, signal_2222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1955 ( .s ({signal_4734, signal_4732}), .b ({signal_3555, signal_2100}), .a ({signal_3536, signal_2081}), .clk (clk), .r (Fresh[241]), .c ({signal_3750, signal_2223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1956 ( .s ({signal_4734, signal_4732}), .b ({signal_4794, signal_4792}), .a ({signal_3556, signal_2101}), .clk (clk), .r (Fresh[242]), .c ({signal_3751, signal_2224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1957 ( .s ({signal_4734, signal_4732}), .b ({signal_3558, signal_2103}), .a ({signal_3557, signal_2102}), .clk (clk), .r (Fresh[243]), .c ({signal_3752, signal_2225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1958 ( .s ({signal_4734, signal_4732}), .b ({signal_4798, signal_4796}), .a ({signal_3559, signal_2104}), .clk (clk), .r (Fresh[244]), .c ({signal_3753, signal_2226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1959 ( .s ({signal_4734, signal_4732}), .b ({signal_3560, signal_2105}), .a ({signal_3526, signal_2071}), .clk (clk), .r (Fresh[245]), .c ({signal_3754, signal_2227}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1960 ( .s ({signal_4734, signal_4732}), .b ({signal_3562, signal_2107}), .a ({signal_3561, signal_2106}), .clk (clk), .r (Fresh[246]), .c ({signal_3755, signal_2228}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1961 ( .s ({signal_4734, signal_4732}), .b ({signal_3556, signal_2101}), .a ({signal_3563, signal_2108}), .clk (clk), .r (Fresh[247]), .c ({signal_3756, signal_2229}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1962 ( .s ({signal_4734, signal_4732}), .b ({signal_4746, signal_4744}), .a ({signal_3564, signal_2109}), .clk (clk), .r (Fresh[248]), .c ({signal_3757, signal_2230}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1963 ( .s ({signal_4734, signal_4732}), .b ({signal_3566, signal_2111}), .a ({signal_3565, signal_2110}), .clk (clk), .r (Fresh[249]), .c ({signal_3758, signal_2231}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1964 ( .s ({signal_4734, signal_4732}), .b ({signal_3568, signal_2113}), .a ({signal_3567, signal_2112}), .clk (clk), .r (Fresh[250]), .c ({signal_3759, signal_2232}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1965 ( .s ({signal_4734, signal_4732}), .b ({signal_3569, signal_2114}), .a ({signal_4802, signal_4800}), .clk (clk), .r (Fresh[251]), .c ({signal_3760, signal_2233}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1966 ( .s ({signal_4734, signal_4732}), .b ({signal_3570, signal_2115}), .a ({signal_3566, signal_2111}), .clk (clk), .r (Fresh[252]), .c ({signal_3761, signal_2234}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1967 ( .s ({signal_4734, signal_4732}), .b ({signal_3525, signal_2070}), .a ({signal_3572, signal_2117}), .clk (clk), .r (Fresh[253]), .c ({signal_3762, signal_2235}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1968 ( .s ({signal_4734, signal_4732}), .b ({signal_3574, signal_2119}), .a ({signal_3573, signal_2118}), .clk (clk), .r (Fresh[254]), .c ({signal_3763, signal_2236}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1969 ( .s ({signal_4734, signal_4732}), .b ({signal_3576, signal_2121}), .a ({signal_3575, signal_2120}), .clk (clk), .r (Fresh[255]), .c ({signal_3764, signal_2237}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1970 ( .s ({signal_4734, signal_4732}), .b ({signal_3563, signal_2108}), .a ({signal_4806, signal_4804}), .clk (clk), .r (Fresh[256]), .c ({signal_3765, signal_2238}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1971 ( .s ({signal_4734, signal_4732}), .b ({signal_3542, signal_2087}), .a ({signal_4810, signal_4808}), .clk (clk), .r (Fresh[257]), .c ({signal_3766, signal_2239}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1972 ( .s ({signal_4734, signal_4732}), .b ({signal_4814, signal_4812}), .a ({signal_3577, signal_2122}), .clk (clk), .r (Fresh[258]), .c ({signal_3767, signal_2240}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1973 ( .s ({signal_4734, signal_4732}), .b ({signal_3566, signal_2111}), .a ({signal_3578, signal_2123}), .clk (clk), .r (Fresh[259]), .c ({signal_3768, signal_2241}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1974 ( .s ({signal_4734, signal_4732}), .b ({signal_3568, signal_2113}), .a ({signal_3536, signal_2081}), .clk (clk), .r (Fresh[260]), .c ({signal_3769, signal_2242}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1975 ( .s ({signal_4734, signal_4732}), .b ({signal_3579, signal_2124}), .a ({signal_4774, signal_4772}), .clk (clk), .r (Fresh[261]), .c ({signal_3770, signal_2243}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1976 ( .s ({signal_4734, signal_4732}), .b ({signal_3581, signal_2126}), .a ({signal_3580, signal_2125}), .clk (clk), .r (Fresh[262]), .c ({signal_3771, signal_2244}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1977 ( .s ({signal_4734, signal_4732}), .b ({signal_3523, signal_2068}), .a ({signal_3582, signal_2127}), .clk (clk), .r (Fresh[263]), .c ({signal_3772, signal_2245}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1978 ( .s ({signal_4734, signal_4732}), .b ({signal_3483, signal_2028}), .a ({signal_3583, signal_2128}), .clk (clk), .r (Fresh[264]), .c ({signal_3773, signal_2246}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1979 ( .s ({signal_4734, signal_4732}), .b ({signal_3585, signal_2130}), .a ({signal_3584, signal_2129}), .clk (clk), .r (Fresh[265]), .c ({signal_3774, signal_2247}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1980 ( .s ({signal_4734, signal_4732}), .b ({signal_3587, signal_2132}), .a ({signal_3586, signal_2131}), .clk (clk), .r (Fresh[266]), .c ({signal_3775, signal_2248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1981 ( .s ({signal_4734, signal_4732}), .b ({signal_3588, signal_2133}), .a ({signal_3504, signal_2049}), .clk (clk), .r (Fresh[267]), .c ({signal_3776, signal_2249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1982 ( .s ({signal_4734, signal_4732}), .b ({signal_3590, signal_2135}), .a ({signal_3589, signal_2134}), .clk (clk), .r (Fresh[268]), .c ({signal_3777, signal_2250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1983 ( .s ({signal_4734, signal_4732}), .b ({signal_3583, signal_2128}), .a ({signal_3579, signal_2124}), .clk (clk), .r (Fresh[269]), .c ({signal_3778, signal_2251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1984 ( .s ({signal_4734, signal_4732}), .b ({signal_3591, signal_2136}), .a ({signal_3554, signal_2099}), .clk (clk), .r (Fresh[270]), .c ({signal_3779, signal_2252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1985 ( .s ({signal_4734, signal_4732}), .b ({signal_3592, signal_2137}), .a ({signal_3527, signal_2072}), .clk (clk), .r (Fresh[271]), .c ({signal_3780, signal_2253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1986 ( .s ({signal_4734, signal_4732}), .b ({signal_3575, signal_2120}), .a ({signal_3593, signal_2138}), .clk (clk), .r (Fresh[272]), .c ({signal_3781, signal_2254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1987 ( .s ({signal_4734, signal_4732}), .b ({signal_3595, signal_2140}), .a ({signal_3594, signal_2139}), .clk (clk), .r (Fresh[273]), .c ({signal_3782, signal_2255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1988 ( .s ({signal_4734, signal_4732}), .b ({signal_3596, signal_2141}), .a ({signal_3583, signal_2128}), .clk (clk), .r (Fresh[274]), .c ({signal_3783, signal_2256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1989 ( .s ({signal_4734, signal_4732}), .b ({signal_3598, signal_2143}), .a ({signal_3597, signal_2142}), .clk (clk), .r (Fresh[275]), .c ({signal_3784, signal_2257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1990 ( .s ({signal_4734, signal_4732}), .b ({signal_3503, signal_2048}), .a ({signal_3599, signal_2144}), .clk (clk), .r (Fresh[276]), .c ({signal_3785, signal_2258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1991 ( .s ({signal_4734, signal_4732}), .b ({signal_3561, signal_2106}), .a ({signal_3543, signal_2088}), .clk (clk), .r (Fresh[277]), .c ({signal_3786, signal_2259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1992 ( .s ({signal_4734, signal_4732}), .b ({signal_3493, signal_2038}), .a ({signal_3600, signal_2145}), .clk (clk), .r (Fresh[278]), .c ({signal_3787, signal_2260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1993 ( .s ({signal_4734, signal_4732}), .b ({signal_3521, signal_2066}), .a ({signal_3503, signal_2048}), .clk (clk), .r (Fresh[279]), .c ({signal_3788, signal_2261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1994 ( .s ({signal_4734, signal_4732}), .b ({signal_3563, signal_2108}), .a ({signal_3539, signal_2084}), .clk (clk), .r (Fresh[280]), .c ({signal_3789, signal_2262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1995 ( .s ({signal_4734, signal_4732}), .b ({signal_4818, signal_4816}), .a ({signal_3518, signal_2063}), .clk (clk), .r (Fresh[281]), .c ({signal_3790, signal_2263}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1996 ( .s ({signal_4734, signal_4732}), .b ({signal_3537, signal_2082}), .a ({signal_4822, signal_4820}), .clk (clk), .r (Fresh[282]), .c ({signal_3791, signal_2264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1997 ( .s ({signal_4734, signal_4732}), .b ({signal_3479, signal_2024}), .a ({signal_4766, signal_4764}), .clk (clk), .r (Fresh[283]), .c ({signal_3792, signal_2265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1998 ( .s ({signal_4734, signal_4732}), .b ({signal_3498, signal_2043}), .a ({signal_4826, signal_4824}), .clk (clk), .r (Fresh[284]), .c ({signal_3793, signal_2266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1999 ( .s ({signal_4734, signal_4732}), .b ({signal_3604, signal_2149}), .a ({signal_3603, signal_2148}), .clk (clk), .r (Fresh[285]), .c ({signal_3794, signal_2267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2000 ( .s ({signal_4734, signal_4732}), .b ({signal_3606, signal_2151}), .a ({signal_3605, signal_2150}), .clk (clk), .r (Fresh[286]), .c ({signal_3795, signal_2268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2001 ( .s ({signal_4734, signal_4732}), .b ({signal_3608, signal_2153}), .a ({signal_3607, signal_2152}), .clk (clk), .r (Fresh[287]), .c ({signal_3796, signal_2269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2002 ( .s ({signal_4734, signal_4732}), .b ({signal_3561, signal_2106}), .a ({signal_3511, signal_2056}), .clk (clk), .r (Fresh[288]), .c ({signal_3797, signal_2270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2003 ( .s ({signal_4734, signal_4732}), .b ({signal_3581, signal_2126}), .a ({signal_3604, signal_2149}), .clk (clk), .r (Fresh[289]), .c ({signal_3798, signal_2271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2004 ( .s ({signal_4734, signal_4732}), .b ({signal_3609, signal_2154}), .a ({signal_3479, signal_2024}), .clk (clk), .r (Fresh[290]), .c ({signal_3799, signal_2272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2005 ( .s ({signal_4734, signal_4732}), .b ({signal_3555, signal_2100}), .a ({signal_3610, signal_2155}), .clk (clk), .r (Fresh[291]), .c ({signal_3800, signal_2273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2006 ( .s ({signal_4734, signal_4732}), .b ({signal_3612, signal_2157}), .a ({signal_3611, signal_2156}), .clk (clk), .r (Fresh[292]), .c ({signal_3801, signal_2274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2007 ( .s ({signal_4734, signal_4732}), .b ({signal_3578, signal_2123}), .a ({signal_3556, signal_2101}), .clk (clk), .r (Fresh[293]), .c ({signal_3802, signal_2275}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2008 ( .s ({signal_4734, signal_4732}), .b ({signal_3612, signal_2157}), .a ({signal_3551, signal_2096}), .clk (clk), .r (Fresh[294]), .c ({signal_3803, signal_2276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2009 ( .s ({signal_4734, signal_4732}), .b ({signal_4790, signal_4788}), .a ({signal_3613, signal_2158}), .clk (clk), .r (Fresh[295]), .c ({signal_3804, signal_2277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2010 ( .s ({signal_4734, signal_4732}), .b ({signal_4810, signal_4808}), .a ({signal_3515, signal_2060}), .clk (clk), .r (Fresh[296]), .c ({signal_3805, signal_2278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2011 ( .s ({signal_4734, signal_4732}), .b ({signal_3614, signal_2159}), .a ({signal_3537, signal_2082}), .clk (clk), .r (Fresh[297]), .c ({signal_3806, signal_2279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2012 ( .s ({signal_4734, signal_4732}), .b ({signal_3615, signal_2160}), .a ({signal_3592, signal_2137}), .clk (clk), .r (Fresh[298]), .c ({signal_3807, signal_2280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2013 ( .s ({signal_4734, signal_4732}), .b ({signal_3617, signal_2162}), .a ({signal_3616, signal_2161}), .clk (clk), .r (Fresh[299]), .c ({signal_3808, signal_2281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2014 ( .s ({signal_4734, signal_4732}), .b ({signal_3618, signal_2163}), .a ({signal_3532, signal_2077}), .clk (clk), .r (Fresh[300]), .c ({signal_3809, signal_2282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2015 ( .s ({signal_4734, signal_4732}), .b ({signal_3619, signal_2164}), .a ({signal_3513, signal_2058}), .clk (clk), .r (Fresh[301]), .c ({signal_3810, signal_2283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2016 ( .s ({signal_4734, signal_4732}), .b ({signal_3620, signal_2165}), .a ({signal_3588, signal_2133}), .clk (clk), .r (Fresh[302]), .c ({signal_3811, signal_2284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2017 ( .s ({signal_4734, signal_4732}), .b ({signal_3484, signal_2029}), .a ({signal_4830, signal_4828}), .clk (clk), .r (Fresh[303]), .c ({signal_3812, signal_2285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2018 ( .s ({signal_4734, signal_4732}), .b ({signal_3621, signal_2166}), .a ({signal_3566, signal_2111}), .clk (clk), .r (Fresh[304]), .c ({signal_3813, signal_2286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2019 ( .s ({signal_4734, signal_4732}), .b ({signal_3622, signal_2167}), .a ({signal_4834, signal_4832}), .clk (clk), .r (Fresh[305]), .c ({signal_3814, signal_2287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2020 ( .s ({signal_4734, signal_4732}), .b ({signal_3623, signal_2168}), .a ({signal_3517, signal_2062}), .clk (clk), .r (Fresh[306]), .c ({signal_3815, signal_2288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2021 ( .s ({signal_4734, signal_4732}), .b ({signal_3625, signal_2170}), .a ({signal_3624, signal_2169}), .clk (clk), .r (Fresh[307]), .c ({signal_3816, signal_2289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2022 ( .s ({signal_4734, signal_4732}), .b ({signal_3609, signal_2154}), .a ({signal_3586, signal_2131}), .clk (clk), .r (Fresh[308]), .c ({signal_3817, signal_2290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2023 ( .s ({signal_4734, signal_4732}), .b ({signal_4838, signal_4836}), .a ({signal_3626, signal_2171}), .clk (clk), .r (Fresh[309]), .c ({signal_3818, signal_2291}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2024 ( .s ({signal_4734, signal_4732}), .b ({signal_4842, signal_4840}), .a ({signal_3625, signal_2170}), .clk (clk), .r (Fresh[310]), .c ({signal_3819, signal_2292}) ) ;
    buf_clk cell_2304 ( .C (clk), .D (signal_4849), .Q (signal_4850) ) ;
    buf_clk cell_2312 ( .C (clk), .D (signal_4857), .Q (signal_4858) ) ;
    buf_clk cell_2314 ( .C (clk), .D (signal_4859), .Q (signal_4860) ) ;
    buf_clk cell_2316 ( .C (clk), .D (signal_4861), .Q (signal_4862) ) ;
    buf_clk cell_2318 ( .C (clk), .D (signal_4863), .Q (signal_4864) ) ;
    buf_clk cell_2320 ( .C (clk), .D (signal_4865), .Q (signal_4866) ) ;
    buf_clk cell_2322 ( .C (clk), .D (signal_4867), .Q (signal_4868) ) ;
    buf_clk cell_2324 ( .C (clk), .D (signal_4869), .Q (signal_4870) ) ;
    buf_clk cell_2326 ( .C (clk), .D (signal_4871), .Q (signal_4872) ) ;
    buf_clk cell_2328 ( .C (clk), .D (signal_4873), .Q (signal_4874) ) ;
    buf_clk cell_2330 ( .C (clk), .D (signal_4875), .Q (signal_4876) ) ;
    buf_clk cell_2332 ( .C (clk), .D (signal_4877), .Q (signal_4878) ) ;
    buf_clk cell_2334 ( .C (clk), .D (signal_4879), .Q (signal_4880) ) ;
    buf_clk cell_2336 ( .C (clk), .D (signal_4881), .Q (signal_4882) ) ;
    buf_clk cell_2338 ( .C (clk), .D (signal_4883), .Q (signal_4884) ) ;
    buf_clk cell_2340 ( .C (clk), .D (signal_4885), .Q (signal_4886) ) ;
    buf_clk cell_2348 ( .C (clk), .D (signal_4893), .Q (signal_4894) ) ;
    buf_clk cell_2358 ( .C (clk), .D (signal_4903), .Q (signal_4904) ) ;
    buf_clk cell_2368 ( .C (clk), .D (signal_4913), .Q (signal_4914) ) ;
    buf_clk cell_2380 ( .C (clk), .D (signal_4925), .Q (signal_4926) ) ;
    buf_clk cell_2392 ( .C (clk), .D (signal_4937), .Q (signal_4938) ) ;
    buf_clk cell_2408 ( .C (clk), .D (signal_4953), .Q (signal_4954) ) ;
    buf_clk cell_2424 ( .C (clk), .D (signal_4969), .Q (signal_4970) ) ;
    buf_clk cell_2440 ( .C (clk), .D (signal_4985), .Q (signal_4986) ) ;
    buf_clk cell_2456 ( .C (clk), .D (signal_5001), .Q (signal_5002) ) ;
    buf_clk cell_2472 ( .C (clk), .D (signal_5017), .Q (signal_5018) ) ;
    buf_clk cell_2488 ( .C (clk), .D (signal_5033), .Q (signal_5034) ) ;
    buf_clk cell_2504 ( .C (clk), .D (signal_5049), .Q (signal_5050) ) ;
    buf_clk cell_2520 ( .C (clk), .D (signal_5065), .Q (signal_5066) ) ;
    buf_clk cell_2536 ( .C (clk), .D (signal_5081), .Q (signal_5082) ) ;
    buf_clk cell_2552 ( .C (clk), .D (signal_5097), .Q (signal_5098) ) ;
    buf_clk cell_2568 ( .C (clk), .D (signal_5113), .Q (signal_5114) ) ;
    buf_clk cell_2584 ( .C (clk), .D (signal_5129), .Q (signal_5130) ) ;
    buf_clk cell_2600 ( .C (clk), .D (signal_5145), .Q (signal_5146) ) ;
    buf_clk cell_2616 ( .C (clk), .D (signal_5161), .Q (signal_5162) ) ;
    buf_clk cell_2632 ( .C (clk), .D (signal_5177), .Q (signal_5178) ) ;
    buf_clk cell_2648 ( .C (clk), .D (signal_5193), .Q (signal_5194) ) ;
    buf_clk cell_2664 ( .C (clk), .D (signal_5209), .Q (signal_5210) ) ;
    buf_clk cell_2680 ( .C (clk), .D (signal_5225), .Q (signal_5226) ) ;
    buf_clk cell_2696 ( .C (clk), .D (signal_5241), .Q (signal_5242) ) ;
    buf_clk cell_2712 ( .C (clk), .D (signal_5257), .Q (signal_5258) ) ;
    buf_clk cell_2728 ( .C (clk), .D (signal_5273), .Q (signal_5274) ) ;
    buf_clk cell_2744 ( .C (clk), .D (signal_5289), .Q (signal_5290) ) ;
    buf_clk cell_2760 ( .C (clk), .D (signal_5305), .Q (signal_5306) ) ;
    buf_clk cell_2776 ( .C (clk), .D (signal_5321), .Q (signal_5322) ) ;
    buf_clk cell_2792 ( .C (clk), .D (signal_5337), .Q (signal_5338) ) ;
    buf_clk cell_2808 ( .C (clk), .D (signal_5353), .Q (signal_5354) ) ;
    buf_clk cell_2824 ( .C (clk), .D (signal_5369), .Q (signal_5370) ) ;
    buf_clk cell_2840 ( .C (clk), .D (signal_5385), .Q (signal_5386) ) ;
    buf_clk cell_2856 ( .C (clk), .D (signal_5401), .Q (signal_5402) ) ;
    buf_clk cell_2872 ( .C (clk), .D (signal_5417), .Q (signal_5418) ) ;
    buf_clk cell_2888 ( .C (clk), .D (signal_5433), .Q (signal_5434) ) ;
    buf_clk cell_2904 ( .C (clk), .D (signal_5449), .Q (signal_5450) ) ;
    buf_clk cell_2920 ( .C (clk), .D (signal_5465), .Q (signal_5466) ) ;
    buf_clk cell_2936 ( .C (clk), .D (signal_5481), .Q (signal_5482) ) ;
    buf_clk cell_2952 ( .C (clk), .D (signal_5497), .Q (signal_5498) ) ;
    buf_clk cell_2968 ( .C (clk), .D (signal_5513), .Q (signal_5514) ) ;
    buf_clk cell_2984 ( .C (clk), .D (signal_5529), .Q (signal_5530) ) ;
    buf_clk cell_3000 ( .C (clk), .D (signal_5545), .Q (signal_5546) ) ;
    buf_clk cell_3016 ( .C (clk), .D (signal_5561), .Q (signal_5562) ) ;
    buf_clk cell_3032 ( .C (clk), .D (signal_5577), .Q (signal_5578) ) ;
    buf_clk cell_3048 ( .C (clk), .D (signal_5593), .Q (signal_5594) ) ;
    buf_clk cell_3064 ( .C (clk), .D (signal_5609), .Q (signal_5610) ) ;
    buf_clk cell_3080 ( .C (clk), .D (signal_5625), .Q (signal_5626) ) ;
    buf_clk cell_3096 ( .C (clk), .D (signal_5641), .Q (signal_5642) ) ;
    buf_clk cell_3112 ( .C (clk), .D (signal_5657), .Q (signal_5658) ) ;
    buf_clk cell_3128 ( .C (clk), .D (signal_5673), .Q (signal_5674) ) ;
    buf_clk cell_3144 ( .C (clk), .D (signal_5689), .Q (signal_5690) ) ;
    buf_clk cell_3160 ( .C (clk), .D (signal_5705), .Q (signal_5706) ) ;
    buf_clk cell_3176 ( .C (clk), .D (signal_5721), .Q (signal_5722) ) ;
    buf_clk cell_3192 ( .C (clk), .D (signal_5737), .Q (signal_5738) ) ;
    buf_clk cell_3208 ( .C (clk), .D (signal_5753), .Q (signal_5754) ) ;
    buf_clk cell_3224 ( .C (clk), .D (signal_5769), .Q (signal_5770) ) ;
    buf_clk cell_3240 ( .C (clk), .D (signal_5785), .Q (signal_5786) ) ;
    buf_clk cell_3256 ( .C (clk), .D (signal_5801), .Q (signal_5802) ) ;
    buf_clk cell_3272 ( .C (clk), .D (signal_5817), .Q (signal_5818) ) ;
    buf_clk cell_3288 ( .C (clk), .D (signal_5833), .Q (signal_5834) ) ;
    buf_clk cell_3304 ( .C (clk), .D (signal_5849), .Q (signal_5850) ) ;
    buf_clk cell_3320 ( .C (clk), .D (signal_5865), .Q (signal_5866) ) ;
    buf_clk cell_3336 ( .C (clk), .D (signal_5881), .Q (signal_5882) ) ;
    buf_clk cell_3352 ( .C (clk), .D (signal_5897), .Q (signal_5898) ) ;
    buf_clk cell_3368 ( .C (clk), .D (signal_5913), .Q (signal_5914) ) ;
    buf_clk cell_3384 ( .C (clk), .D (signal_5929), .Q (signal_5930) ) ;
    buf_clk cell_3400 ( .C (clk), .D (signal_5945), .Q (signal_5946) ) ;
    buf_clk cell_3416 ( .C (clk), .D (signal_5961), .Q (signal_5962) ) ;
    buf_clk cell_3432 ( .C (clk), .D (signal_5977), .Q (signal_5978) ) ;
    buf_clk cell_3448 ( .C (clk), .D (signal_5993), .Q (signal_5994) ) ;
    buf_clk cell_3464 ( .C (clk), .D (signal_6009), .Q (signal_6010) ) ;
    buf_clk cell_3480 ( .C (clk), .D (signal_6025), .Q (signal_6026) ) ;
    buf_clk cell_3496 ( .C (clk), .D (signal_6041), .Q (signal_6042) ) ;
    buf_clk cell_3512 ( .C (clk), .D (signal_6057), .Q (signal_6058) ) ;
    buf_clk cell_3528 ( .C (clk), .D (signal_6073), .Q (signal_6074) ) ;
    buf_clk cell_3544 ( .C (clk), .D (signal_6089), .Q (signal_6090) ) ;
    buf_clk cell_3560 ( .C (clk), .D (signal_6105), .Q (signal_6106) ) ;
    buf_clk cell_3576 ( .C (clk), .D (signal_6121), .Q (signal_6122) ) ;
    buf_clk cell_3592 ( .C (clk), .D (signal_6137), .Q (signal_6138) ) ;
    buf_clk cell_3608 ( .C (clk), .D (signal_6153), .Q (signal_6154) ) ;
    buf_clk cell_3624 ( .C (clk), .D (signal_6169), .Q (signal_6170) ) ;
    buf_clk cell_3640 ( .C (clk), .D (signal_6185), .Q (signal_6186) ) ;
    buf_clk cell_3656 ( .C (clk), .D (signal_6201), .Q (signal_6202) ) ;
    buf_clk cell_3672 ( .C (clk), .D (signal_6217), .Q (signal_6218) ) ;
    buf_clk cell_3688 ( .C (clk), .D (signal_6233), .Q (signal_6234) ) ;
    buf_clk cell_3704 ( .C (clk), .D (signal_6249), .Q (signal_6250) ) ;
    buf_clk cell_3720 ( .C (clk), .D (signal_6265), .Q (signal_6266) ) ;
    buf_clk cell_3736 ( .C (clk), .D (signal_6281), .Q (signal_6282) ) ;
    buf_clk cell_3752 ( .C (clk), .D (signal_6297), .Q (signal_6298) ) ;
    buf_clk cell_3768 ( .C (clk), .D (signal_6313), .Q (signal_6314) ) ;
    buf_clk cell_3784 ( .C (clk), .D (signal_6329), .Q (signal_6330) ) ;
    buf_clk cell_3800 ( .C (clk), .D (signal_6345), .Q (signal_6346) ) ;
    buf_clk cell_3816 ( .C (clk), .D (signal_6361), .Q (signal_6362) ) ;
    buf_clk cell_3832 ( .C (clk), .D (signal_6377), .Q (signal_6378) ) ;
    buf_clk cell_3848 ( .C (clk), .D (signal_6393), .Q (signal_6394) ) ;
    buf_clk cell_3864 ( .C (clk), .D (signal_6409), .Q (signal_6410) ) ;
    buf_clk cell_3880 ( .C (clk), .D (signal_6425), .Q (signal_6426) ) ;
    buf_clk cell_3896 ( .C (clk), .D (signal_6441), .Q (signal_6442) ) ;
    buf_clk cell_3912 ( .C (clk), .D (signal_6457), .Q (signal_6458) ) ;
    buf_clk cell_3928 ( .C (clk), .D (signal_6473), .Q (signal_6474) ) ;
    buf_clk cell_3944 ( .C (clk), .D (signal_6489), .Q (signal_6490) ) ;
    buf_clk cell_3960 ( .C (clk), .D (signal_6505), .Q (signal_6506) ) ;
    buf_clk cell_3976 ( .C (clk), .D (signal_6521), .Q (signal_6522) ) ;
    buf_clk cell_3992 ( .C (clk), .D (signal_6537), .Q (signal_6538) ) ;
    buf_clk cell_4008 ( .C (clk), .D (signal_6553), .Q (signal_6554) ) ;
    buf_clk cell_4024 ( .C (clk), .D (signal_6569), .Q (signal_6570) ) ;
    buf_clk cell_4040 ( .C (clk), .D (signal_6585), .Q (signal_6586) ) ;
    buf_clk cell_4056 ( .C (clk), .D (signal_6601), .Q (signal_6602) ) ;
    buf_clk cell_4072 ( .C (clk), .D (signal_6617), .Q (signal_6618) ) ;
    buf_clk cell_4088 ( .C (clk), .D (signal_6633), .Q (signal_6634) ) ;
    buf_clk cell_4104 ( .C (clk), .D (signal_6649), .Q (signal_6650) ) ;
    buf_clk cell_4120 ( .C (clk), .D (signal_6665), .Q (signal_6666) ) ;
    buf_clk cell_4136 ( .C (clk), .D (signal_6681), .Q (signal_6682) ) ;
    buf_clk cell_4152 ( .C (clk), .D (signal_6697), .Q (signal_6698) ) ;
    buf_clk cell_4168 ( .C (clk), .D (signal_6713), .Q (signal_6714) ) ;
    buf_clk cell_4184 ( .C (clk), .D (signal_6729), .Q (signal_6730) ) ;
    buf_clk cell_4200 ( .C (clk), .D (signal_6745), .Q (signal_6746) ) ;
    buf_clk cell_4216 ( .C (clk), .D (signal_6761), .Q (signal_6762) ) ;
    buf_clk cell_4232 ( .C (clk), .D (signal_6777), .Q (signal_6778) ) ;
    buf_clk cell_4248 ( .C (clk), .D (signal_6793), .Q (signal_6794) ) ;
    buf_clk cell_4264 ( .C (clk), .D (signal_6809), .Q (signal_6810) ) ;
    buf_clk cell_4280 ( .C (clk), .D (signal_6825), .Q (signal_6826) ) ;
    buf_clk cell_4296 ( .C (clk), .D (signal_6841), .Q (signal_6842) ) ;
    buf_clk cell_4312 ( .C (clk), .D (signal_6857), .Q (signal_6858) ) ;
    buf_clk cell_4328 ( .C (clk), .D (signal_6873), .Q (signal_6874) ) ;
    buf_clk cell_4344 ( .C (clk), .D (signal_6889), .Q (signal_6890) ) ;
    buf_clk cell_4360 ( .C (clk), .D (signal_6905), .Q (signal_6906) ) ;
    buf_clk cell_4376 ( .C (clk), .D (signal_6921), .Q (signal_6922) ) ;
    buf_clk cell_4392 ( .C (clk), .D (signal_6937), .Q (signal_6938) ) ;
    buf_clk cell_4408 ( .C (clk), .D (signal_6953), .Q (signal_6954) ) ;
    buf_clk cell_4422 ( .C (clk), .D (signal_6967), .Q (signal_6968) ) ;
    buf_clk cell_4436 ( .C (clk), .D (signal_6981), .Q (signal_6982) ) ;
    buf_clk cell_4452 ( .C (clk), .D (signal_6997), .Q (signal_6998) ) ;
    buf_clk cell_4468 ( .C (clk), .D (signal_7013), .Q (signal_7014) ) ;
    buf_clk cell_4484 ( .C (clk), .D (signal_7029), .Q (signal_7030) ) ;
    buf_clk cell_4500 ( .C (clk), .D (signal_7045), .Q (signal_7046) ) ;
    buf_clk cell_4516 ( .C (clk), .D (signal_7061), .Q (signal_7062) ) ;
    buf_clk cell_4532 ( .C (clk), .D (signal_7077), .Q (signal_7078) ) ;
    buf_clk cell_4548 ( .C (clk), .D (signal_7093), .Q (signal_7094) ) ;
    buf_clk cell_4564 ( .C (clk), .D (signal_7109), .Q (signal_7110) ) ;
    buf_clk cell_4580 ( .C (clk), .D (signal_7125), .Q (signal_7126) ) ;
    buf_clk cell_4596 ( .C (clk), .D (signal_7141), .Q (signal_7142) ) ;
    buf_clk cell_4612 ( .C (clk), .D (signal_7157), .Q (signal_7158) ) ;
    buf_clk cell_4628 ( .C (clk), .D (signal_7173), .Q (signal_7174) ) ;
    buf_clk cell_4644 ( .C (clk), .D (signal_7189), .Q (signal_7190) ) ;
    buf_clk cell_4660 ( .C (clk), .D (signal_7205), .Q (signal_7206) ) ;
    buf_clk cell_4676 ( .C (clk), .D (signal_7221), .Q (signal_7222) ) ;
    buf_clk cell_4692 ( .C (clk), .D (signal_7237), .Q (signal_7238) ) ;
    buf_clk cell_4708 ( .C (clk), .D (signal_7253), .Q (signal_7254) ) ;
    buf_clk cell_4724 ( .C (clk), .D (signal_7269), .Q (signal_7270) ) ;
    buf_clk cell_4740 ( .C (clk), .D (signal_7285), .Q (signal_7286) ) ;
    buf_clk cell_4756 ( .C (clk), .D (signal_7301), .Q (signal_7302) ) ;
    buf_clk cell_4772 ( .C (clk), .D (signal_7317), .Q (signal_7318) ) ;
    buf_clk cell_4788 ( .C (clk), .D (signal_7333), .Q (signal_7334) ) ;
    buf_clk cell_4804 ( .C (clk), .D (signal_7349), .Q (signal_7350) ) ;
    buf_clk cell_4820 ( .C (clk), .D (signal_7365), .Q (signal_7366) ) ;
    buf_clk cell_4836 ( .C (clk), .D (signal_7381), .Q (signal_7382) ) ;
    buf_clk cell_4852 ( .C (clk), .D (signal_7397), .Q (signal_7398) ) ;
    buf_clk cell_4868 ( .C (clk), .D (signal_7413), .Q (signal_7414) ) ;
    buf_clk cell_4884 ( .C (clk), .D (signal_7429), .Q (signal_7430) ) ;
    buf_clk cell_4900 ( .C (clk), .D (signal_7445), .Q (signal_7446) ) ;
    buf_clk cell_4916 ( .C (clk), .D (signal_7461), .Q (signal_7462) ) ;
    buf_clk cell_4932 ( .C (clk), .D (signal_7477), .Q (signal_7478) ) ;
    buf_clk cell_4948 ( .C (clk), .D (signal_7493), .Q (signal_7494) ) ;
    buf_clk cell_4964 ( .C (clk), .D (signal_7509), .Q (signal_7510) ) ;
    buf_clk cell_4980 ( .C (clk), .D (signal_7525), .Q (signal_7526) ) ;
    buf_clk cell_4996 ( .C (clk), .D (signal_7541), .Q (signal_7542) ) ;
    buf_clk cell_5012 ( .C (clk), .D (signal_7557), .Q (signal_7558) ) ;
    buf_clk cell_5028 ( .C (clk), .D (signal_7573), .Q (signal_7574) ) ;
    buf_clk cell_5044 ( .C (clk), .D (signal_7589), .Q (signal_7590) ) ;
    buf_clk cell_5060 ( .C (clk), .D (signal_7605), .Q (signal_7606) ) ;
    buf_clk cell_5076 ( .C (clk), .D (signal_7621), .Q (signal_7622) ) ;
    buf_clk cell_5092 ( .C (clk), .D (signal_7637), .Q (signal_7638) ) ;
    buf_clk cell_5108 ( .C (clk), .D (signal_7653), .Q (signal_7654) ) ;
    buf_clk cell_5124 ( .C (clk), .D (signal_7669), .Q (signal_7670) ) ;
    buf_clk cell_5140 ( .C (clk), .D (signal_7685), .Q (signal_7686) ) ;
    buf_clk cell_5156 ( .C (clk), .D (signal_7701), .Q (signal_7702) ) ;
    buf_clk cell_5172 ( .C (clk), .D (signal_7717), .Q (signal_7718) ) ;
    buf_clk cell_5188 ( .C (clk), .D (signal_7733), .Q (signal_7734) ) ;
    buf_clk cell_5204 ( .C (clk), .D (signal_7749), .Q (signal_7750) ) ;
    buf_clk cell_5220 ( .C (clk), .D (signal_7765), .Q (signal_7766) ) ;
    buf_clk cell_5236 ( .C (clk), .D (signal_7781), .Q (signal_7782) ) ;
    buf_clk cell_5252 ( .C (clk), .D (signal_7797), .Q (signal_7798) ) ;
    buf_clk cell_5268 ( .C (clk), .D (signal_7813), .Q (signal_7814) ) ;
    buf_clk cell_5284 ( .C (clk), .D (signal_7829), .Q (signal_7830) ) ;
    buf_clk cell_5300 ( .C (clk), .D (signal_7845), .Q (signal_7846) ) ;
    buf_clk cell_5316 ( .C (clk), .D (signal_7861), .Q (signal_7862) ) ;
    buf_clk cell_5332 ( .C (clk), .D (signal_7877), .Q (signal_7878) ) ;
    buf_clk cell_5348 ( .C (clk), .D (signal_7893), .Q (signal_7894) ) ;
    buf_clk cell_5364 ( .C (clk), .D (signal_7909), .Q (signal_7910) ) ;
    buf_clk cell_5380 ( .C (clk), .D (signal_7925), .Q (signal_7926) ) ;
    buf_clk cell_5396 ( .C (clk), .D (signal_7941), .Q (signal_7942) ) ;
    buf_clk cell_5412 ( .C (clk), .D (signal_7957), .Q (signal_7958) ) ;
    buf_clk cell_5428 ( .C (clk), .D (signal_7973), .Q (signal_7974) ) ;
    buf_clk cell_5444 ( .C (clk), .D (signal_7989), .Q (signal_7990) ) ;
    buf_clk cell_5460 ( .C (clk), .D (signal_8005), .Q (signal_8006) ) ;
    buf_clk cell_5476 ( .C (clk), .D (signal_8021), .Q (signal_8022) ) ;
    buf_clk cell_5492 ( .C (clk), .D (signal_8037), .Q (signal_8038) ) ;
    buf_clk cell_5508 ( .C (clk), .D (signal_8053), .Q (signal_8054) ) ;
    buf_clk cell_5524 ( .C (clk), .D (signal_8069), .Q (signal_8070) ) ;
    buf_clk cell_5540 ( .C (clk), .D (signal_8085), .Q (signal_8086) ) ;
    buf_clk cell_5556 ( .C (clk), .D (signal_8101), .Q (signal_8102) ) ;
    buf_clk cell_5572 ( .C (clk), .D (signal_8117), .Q (signal_8118) ) ;
    buf_clk cell_5588 ( .C (clk), .D (signal_8133), .Q (signal_8134) ) ;
    buf_clk cell_5604 ( .C (clk), .D (signal_8149), .Q (signal_8150) ) ;
    buf_clk cell_5620 ( .C (clk), .D (signal_8165), .Q (signal_8166) ) ;
    buf_clk cell_5636 ( .C (clk), .D (signal_8181), .Q (signal_8182) ) ;
    buf_clk cell_5652 ( .C (clk), .D (signal_8197), .Q (signal_8198) ) ;
    buf_clk cell_5668 ( .C (clk), .D (signal_8213), .Q (signal_8214) ) ;
    buf_clk cell_5684 ( .C (clk), .D (signal_8229), .Q (signal_8230) ) ;
    buf_clk cell_5700 ( .C (clk), .D (signal_8245), .Q (signal_8246) ) ;
    buf_clk cell_5716 ( .C (clk), .D (signal_8261), .Q (signal_8262) ) ;
    buf_clk cell_5732 ( .C (clk), .D (signal_8277), .Q (signal_8278) ) ;
    buf_clk cell_5748 ( .C (clk), .D (signal_8293), .Q (signal_8294) ) ;
    buf_clk cell_5764 ( .C (clk), .D (signal_8309), .Q (signal_8310) ) ;
    buf_clk cell_5780 ( .C (clk), .D (signal_8325), .Q (signal_8326) ) ;
    buf_clk cell_5796 ( .C (clk), .D (signal_8341), .Q (signal_8342) ) ;
    buf_clk cell_5812 ( .C (clk), .D (signal_8357), .Q (signal_8358) ) ;
    buf_clk cell_5828 ( .C (clk), .D (signal_8373), .Q (signal_8374) ) ;
    buf_clk cell_5844 ( .C (clk), .D (signal_8389), .Q (signal_8390) ) ;
    buf_clk cell_5860 ( .C (clk), .D (signal_8405), .Q (signal_8406) ) ;
    buf_clk cell_5876 ( .C (clk), .D (signal_8421), .Q (signal_8422) ) ;
    buf_clk cell_5892 ( .C (clk), .D (signal_8437), .Q (signal_8438) ) ;
    buf_clk cell_5908 ( .C (clk), .D (signal_8453), .Q (signal_8454) ) ;
    buf_clk cell_5924 ( .C (clk), .D (signal_8469), .Q (signal_8470) ) ;
    buf_clk cell_5940 ( .C (clk), .D (signal_8485), .Q (signal_8486) ) ;
    buf_clk cell_5956 ( .C (clk), .D (signal_8501), .Q (signal_8502) ) ;
    buf_clk cell_5972 ( .C (clk), .D (signal_8517), .Q (signal_8518) ) ;
    buf_clk cell_5988 ( .C (clk), .D (signal_8533), .Q (signal_8534) ) ;
    buf_clk cell_6004 ( .C (clk), .D (signal_8549), .Q (signal_8550) ) ;
    buf_clk cell_6020 ( .C (clk), .D (signal_8565), .Q (signal_8566) ) ;
    buf_clk cell_6036 ( .C (clk), .D (signal_8581), .Q (signal_8582) ) ;
    buf_clk cell_6052 ( .C (clk), .D (signal_8597), .Q (signal_8598) ) ;
    buf_clk cell_6068 ( .C (clk), .D (signal_8613), .Q (signal_8614) ) ;
    buf_clk cell_6084 ( .C (clk), .D (signal_8629), .Q (signal_8630) ) ;
    buf_clk cell_6100 ( .C (clk), .D (signal_8645), .Q (signal_8646) ) ;
    buf_clk cell_6116 ( .C (clk), .D (signal_8661), .Q (signal_8662) ) ;
    buf_clk cell_6132 ( .C (clk), .D (signal_8677), .Q (signal_8678) ) ;
    buf_clk cell_6148 ( .C (clk), .D (signal_8693), .Q (signal_8694) ) ;
    buf_clk cell_6164 ( .C (clk), .D (signal_8709), .Q (signal_8710) ) ;
    buf_clk cell_6180 ( .C (clk), .D (signal_8725), .Q (signal_8726) ) ;
    buf_clk cell_6196 ( .C (clk), .D (signal_8741), .Q (signal_8742) ) ;
    buf_clk cell_6212 ( .C (clk), .D (signal_8757), .Q (signal_8758) ) ;
    buf_clk cell_6228 ( .C (clk), .D (signal_8773), .Q (signal_8774) ) ;
    buf_clk cell_6244 ( .C (clk), .D (signal_8789), .Q (signal_8790) ) ;
    buf_clk cell_6260 ( .C (clk), .D (signal_8805), .Q (signal_8806) ) ;
    buf_clk cell_6276 ( .C (clk), .D (signal_8821), .Q (signal_8822) ) ;
    buf_clk cell_6292 ( .C (clk), .D (signal_8837), .Q (signal_8838) ) ;
    buf_clk cell_6308 ( .C (clk), .D (signal_8853), .Q (signal_8854) ) ;
    buf_clk cell_6324 ( .C (clk), .D (signal_8869), .Q (signal_8870) ) ;
    buf_clk cell_6340 ( .C (clk), .D (signal_8885), .Q (signal_8886) ) ;
    buf_clk cell_6356 ( .C (clk), .D (signal_8901), .Q (signal_8902) ) ;
    buf_clk cell_6372 ( .C (clk), .D (signal_8917), .Q (signal_8918) ) ;
    buf_clk cell_6388 ( .C (clk), .D (signal_8933), .Q (signal_8934) ) ;
    buf_clk cell_6404 ( .C (clk), .D (signal_8949), .Q (signal_8950) ) ;
    buf_clk cell_6420 ( .C (clk), .D (signal_8965), .Q (signal_8966) ) ;
    buf_clk cell_6436 ( .C (clk), .D (signal_8981), .Q (signal_8982) ) ;
    buf_clk cell_6452 ( .C (clk), .D (signal_8997), .Q (signal_8998) ) ;
    buf_clk cell_6468 ( .C (clk), .D (signal_9013), .Q (signal_9014) ) ;
    buf_clk cell_6484 ( .C (clk), .D (signal_9029), .Q (signal_9030) ) ;
    buf_clk cell_6500 ( .C (clk), .D (signal_9045), .Q (signal_9046) ) ;
    buf_clk cell_6516 ( .C (clk), .D (signal_9061), .Q (signal_9062) ) ;
    buf_clk cell_6532 ( .C (clk), .D (signal_9077), .Q (signal_9078) ) ;
    buf_clk cell_6548 ( .C (clk), .D (signal_9093), .Q (signal_9094) ) ;
    buf_clk cell_6564 ( .C (clk), .D (signal_9109), .Q (signal_9110) ) ;
    buf_clk cell_6580 ( .C (clk), .D (signal_9125), .Q (signal_9126) ) ;
    buf_clk cell_6596 ( .C (clk), .D (signal_9141), .Q (signal_9142) ) ;
    buf_clk cell_6612 ( .C (clk), .D (signal_9157), .Q (signal_9158) ) ;
    buf_clk cell_6628 ( .C (clk), .D (signal_9173), .Q (signal_9174) ) ;
    buf_clk cell_6644 ( .C (clk), .D (signal_9189), .Q (signal_9190) ) ;
    buf_clk cell_6660 ( .C (clk), .D (signal_9205), .Q (signal_9206) ) ;
    buf_clk cell_6676 ( .C (clk), .D (signal_9221), .Q (signal_9222) ) ;
    buf_clk cell_6692 ( .C (clk), .D (signal_9237), .Q (signal_9238) ) ;
    buf_clk cell_6708 ( .C (clk), .D (signal_9253), .Q (signal_9254) ) ;
    buf_clk cell_6724 ( .C (clk), .D (signal_9269), .Q (signal_9270) ) ;
    buf_clk cell_6740 ( .C (clk), .D (signal_9285), .Q (signal_9286) ) ;
    buf_clk cell_6756 ( .C (clk), .D (signal_9301), .Q (signal_9302) ) ;
    buf_clk cell_6772 ( .C (clk), .D (signal_9317), .Q (signal_9318) ) ;
    buf_clk cell_6788 ( .C (clk), .D (signal_9333), .Q (signal_9334) ) ;
    buf_clk cell_6804 ( .C (clk), .D (signal_9349), .Q (signal_9350) ) ;
    buf_clk cell_6820 ( .C (clk), .D (signal_9365), .Q (signal_9366) ) ;
    buf_clk cell_6836 ( .C (clk), .D (signal_9381), .Q (signal_9382) ) ;
    buf_clk cell_6852 ( .C (clk), .D (signal_9397), .Q (signal_9398) ) ;
    buf_clk cell_6868 ( .C (clk), .D (signal_9413), .Q (signal_9414) ) ;
    buf_clk cell_6884 ( .C (clk), .D (signal_9429), .Q (signal_9430) ) ;
    buf_clk cell_6900 ( .C (clk), .D (signal_9445), .Q (signal_9446) ) ;
    buf_clk cell_6916 ( .C (clk), .D (signal_9461), .Q (signal_9462) ) ;
    buf_clk cell_6932 ( .C (clk), .D (signal_9477), .Q (signal_9478) ) ;
    buf_clk cell_6948 ( .C (clk), .D (signal_9493), .Q (signal_9494) ) ;
    buf_clk cell_6964 ( .C (clk), .D (signal_9509), .Q (signal_9510) ) ;
    buf_clk cell_6980 ( .C (clk), .D (signal_9525), .Q (signal_9526) ) ;
    buf_clk cell_6996 ( .C (clk), .D (signal_9541), .Q (signal_9542) ) ;
    buf_clk cell_7012 ( .C (clk), .D (signal_9557), .Q (signal_9558) ) ;
    buf_clk cell_7028 ( .C (clk), .D (signal_9573), .Q (signal_9574) ) ;
    buf_clk cell_7044 ( .C (clk), .D (signal_9589), .Q (signal_9590) ) ;
    buf_clk cell_7060 ( .C (clk), .D (signal_9605), .Q (signal_9606) ) ;
    buf_clk cell_7076 ( .C (clk), .D (signal_9621), .Q (signal_9622) ) ;
    buf_clk cell_7092 ( .C (clk), .D (signal_9637), .Q (signal_9638) ) ;
    buf_clk cell_7108 ( .C (clk), .D (signal_9653), .Q (signal_9654) ) ;
    buf_clk cell_7124 ( .C (clk), .D (signal_9669), .Q (signal_9670) ) ;
    buf_clk cell_7140 ( .C (clk), .D (signal_9685), .Q (signal_9686) ) ;
    buf_clk cell_7156 ( .C (clk), .D (signal_9701), .Q (signal_9702) ) ;
    buf_clk cell_7172 ( .C (clk), .D (signal_9717), .Q (signal_9718) ) ;
    buf_clk cell_7188 ( .C (clk), .D (signal_9733), .Q (signal_9734) ) ;
    buf_clk cell_7204 ( .C (clk), .D (signal_9749), .Q (signal_9750) ) ;
    buf_clk cell_7220 ( .C (clk), .D (signal_9765), .Q (signal_9766) ) ;
    buf_clk cell_7236 ( .C (clk), .D (signal_9781), .Q (signal_9782) ) ;
    buf_clk cell_7252 ( .C (clk), .D (signal_9797), .Q (signal_9798) ) ;
    buf_clk cell_7268 ( .C (clk), .D (signal_9813), .Q (signal_9814) ) ;
    buf_clk cell_7284 ( .C (clk), .D (signal_9829), .Q (signal_9830) ) ;
    buf_clk cell_7300 ( .C (clk), .D (signal_9845), .Q (signal_9846) ) ;
    buf_clk cell_7316 ( .C (clk), .D (signal_9861), .Q (signal_9862) ) ;
    buf_clk cell_7332 ( .C (clk), .D (signal_9877), .Q (signal_9878) ) ;
    buf_clk cell_7348 ( .C (clk), .D (signal_9893), .Q (signal_9894) ) ;
    buf_clk cell_7364 ( .C (clk), .D (signal_9909), .Q (signal_9910) ) ;
    buf_clk cell_7380 ( .C (clk), .D (signal_9925), .Q (signal_9926) ) ;
    buf_clk cell_7396 ( .C (clk), .D (signal_9941), .Q (signal_9942) ) ;
    buf_clk cell_7412 ( .C (clk), .D (signal_9957), .Q (signal_9958) ) ;
    buf_clk cell_7428 ( .C (clk), .D (signal_9973), .Q (signal_9974) ) ;
    buf_clk cell_7444 ( .C (clk), .D (signal_9989), .Q (signal_9990) ) ;
    buf_clk cell_7460 ( .C (clk), .D (signal_10005), .Q (signal_10006) ) ;
    buf_clk cell_7476 ( .C (clk), .D (signal_10021), .Q (signal_10022) ) ;
    buf_clk cell_7492 ( .C (clk), .D (signal_10037), .Q (signal_10038) ) ;
    buf_clk cell_7508 ( .C (clk), .D (signal_10053), .Q (signal_10054) ) ;
    buf_clk cell_7524 ( .C (clk), .D (signal_10069), .Q (signal_10070) ) ;
    buf_clk cell_7540 ( .C (clk), .D (signal_10085), .Q (signal_10086) ) ;
    buf_clk cell_7556 ( .C (clk), .D (signal_10101), .Q (signal_10102) ) ;
    buf_clk cell_7572 ( .C (clk), .D (signal_10117), .Q (signal_10118) ) ;
    buf_clk cell_7588 ( .C (clk), .D (signal_10133), .Q (signal_10134) ) ;
    buf_clk cell_7604 ( .C (clk), .D (signal_10149), .Q (signal_10150) ) ;
    buf_clk cell_7620 ( .C (clk), .D (signal_10165), .Q (signal_10166) ) ;
    buf_clk cell_7636 ( .C (clk), .D (signal_10181), .Q (signal_10182) ) ;
    buf_clk cell_7652 ( .C (clk), .D (signal_10197), .Q (signal_10198) ) ;
    buf_clk cell_7668 ( .C (clk), .D (signal_10213), .Q (signal_10214) ) ;
    buf_clk cell_7684 ( .C (clk), .D (signal_10229), .Q (signal_10230) ) ;
    buf_clk cell_7700 ( .C (clk), .D (signal_10245), .Q (signal_10246) ) ;
    buf_clk cell_7716 ( .C (clk), .D (signal_10261), .Q (signal_10262) ) ;
    buf_clk cell_7732 ( .C (clk), .D (signal_10277), .Q (signal_10278) ) ;
    buf_clk cell_7748 ( .C (clk), .D (signal_10293), .Q (signal_10294) ) ;
    buf_clk cell_7764 ( .C (clk), .D (signal_10309), .Q (signal_10310) ) ;
    buf_clk cell_7780 ( .C (clk), .D (signal_10325), .Q (signal_10326) ) ;
    buf_clk cell_7796 ( .C (clk), .D (signal_10341), .Q (signal_10342) ) ;
    buf_clk cell_7812 ( .C (clk), .D (signal_10357), .Q (signal_10358) ) ;
    buf_clk cell_7828 ( .C (clk), .D (signal_10373), .Q (signal_10374) ) ;
    buf_clk cell_7844 ( .C (clk), .D (signal_10389), .Q (signal_10390) ) ;
    buf_clk cell_7860 ( .C (clk), .D (signal_10405), .Q (signal_10406) ) ;
    buf_clk cell_7876 ( .C (clk), .D (signal_10421), .Q (signal_10422) ) ;
    buf_clk cell_7892 ( .C (clk), .D (signal_10437), .Q (signal_10438) ) ;
    buf_clk cell_7908 ( .C (clk), .D (signal_10453), .Q (signal_10454) ) ;
    buf_clk cell_7924 ( .C (clk), .D (signal_10469), .Q (signal_10470) ) ;
    buf_clk cell_7940 ( .C (clk), .D (signal_10485), .Q (signal_10486) ) ;
    buf_clk cell_7956 ( .C (clk), .D (signal_10501), .Q (signal_10502) ) ;
    buf_clk cell_7972 ( .C (clk), .D (signal_10517), .Q (signal_10518) ) ;
    buf_clk cell_7988 ( .C (clk), .D (signal_10533), .Q (signal_10534) ) ;
    buf_clk cell_8004 ( .C (clk), .D (signal_10549), .Q (signal_10550) ) ;
    buf_clk cell_8020 ( .C (clk), .D (signal_10565), .Q (signal_10566) ) ;
    buf_clk cell_8036 ( .C (clk), .D (signal_10581), .Q (signal_10582) ) ;
    buf_clk cell_8052 ( .C (clk), .D (signal_10597), .Q (signal_10598) ) ;
    buf_clk cell_8068 ( .C (clk), .D (signal_10613), .Q (signal_10614) ) ;
    buf_clk cell_8084 ( .C (clk), .D (signal_10629), .Q (signal_10630) ) ;
    buf_clk cell_8100 ( .C (clk), .D (signal_10645), .Q (signal_10646) ) ;
    buf_clk cell_8116 ( .C (clk), .D (signal_10661), .Q (signal_10662) ) ;
    buf_clk cell_8132 ( .C (clk), .D (signal_10677), .Q (signal_10678) ) ;
    buf_clk cell_8148 ( .C (clk), .D (signal_10693), .Q (signal_10694) ) ;
    buf_clk cell_8164 ( .C (clk), .D (signal_10709), .Q (signal_10710) ) ;
    buf_clk cell_8180 ( .C (clk), .D (signal_10725), .Q (signal_10726) ) ;
    buf_clk cell_8196 ( .C (clk), .D (signal_10741), .Q (signal_10742) ) ;
    buf_clk cell_8212 ( .C (clk), .D (signal_10757), .Q (signal_10758) ) ;
    buf_clk cell_8228 ( .C (clk), .D (signal_10773), .Q (signal_10774) ) ;
    buf_clk cell_8244 ( .C (clk), .D (signal_10789), .Q (signal_10790) ) ;
    buf_clk cell_8260 ( .C (clk), .D (signal_10805), .Q (signal_10806) ) ;
    buf_clk cell_8276 ( .C (clk), .D (signal_10821), .Q (signal_10822) ) ;
    buf_clk cell_8292 ( .C (clk), .D (signal_10837), .Q (signal_10838) ) ;
    buf_clk cell_8308 ( .C (clk), .D (signal_10853), .Q (signal_10854) ) ;
    buf_clk cell_8324 ( .C (clk), .D (signal_10869), .Q (signal_10870) ) ;
    buf_clk cell_8340 ( .C (clk), .D (signal_10885), .Q (signal_10886) ) ;
    buf_clk cell_8356 ( .C (clk), .D (signal_10901), .Q (signal_10902) ) ;
    buf_clk cell_8372 ( .C (clk), .D (signal_10917), .Q (signal_10918) ) ;
    buf_clk cell_8388 ( .C (clk), .D (signal_10933), .Q (signal_10934) ) ;
    buf_clk cell_8404 ( .C (clk), .D (signal_10949), .Q (signal_10950) ) ;
    buf_clk cell_8420 ( .C (clk), .D (signal_10965), .Q (signal_10966) ) ;
    buf_clk cell_8436 ( .C (clk), .D (signal_10981), .Q (signal_10982) ) ;
    buf_clk cell_8452 ( .C (clk), .D (signal_10997), .Q (signal_10998) ) ;
    buf_clk cell_8468 ( .C (clk), .D (signal_11013), .Q (signal_11014) ) ;
    buf_clk cell_8484 ( .C (clk), .D (signal_11029), .Q (signal_11030) ) ;
    buf_clk cell_8500 ( .C (clk), .D (signal_11045), .Q (signal_11046) ) ;
    buf_clk cell_8516 ( .C (clk), .D (signal_11061), .Q (signal_11062) ) ;
    buf_clk cell_8532 ( .C (clk), .D (signal_11077), .Q (signal_11078) ) ;
    buf_clk cell_8548 ( .C (clk), .D (signal_11093), .Q (signal_11094) ) ;
    buf_clk cell_8564 ( .C (clk), .D (signal_11109), .Q (signal_11110) ) ;
    buf_clk cell_8580 ( .C (clk), .D (signal_11125), .Q (signal_11126) ) ;
    buf_clk cell_8596 ( .C (clk), .D (signal_11141), .Q (signal_11142) ) ;
    buf_clk cell_8612 ( .C (clk), .D (signal_11157), .Q (signal_11158) ) ;
    buf_clk cell_8628 ( .C (clk), .D (signal_11173), .Q (signal_11174) ) ;
    buf_clk cell_8644 ( .C (clk), .D (signal_11189), .Q (signal_11190) ) ;
    buf_clk cell_8660 ( .C (clk), .D (signal_11205), .Q (signal_11206) ) ;
    buf_clk cell_8676 ( .C (clk), .D (signal_11221), .Q (signal_11222) ) ;
    buf_clk cell_8692 ( .C (clk), .D (signal_11237), .Q (signal_11238) ) ;
    buf_clk cell_8708 ( .C (clk), .D (signal_11253), .Q (signal_11254) ) ;
    buf_clk cell_8724 ( .C (clk), .D (signal_11269), .Q (signal_11270) ) ;
    buf_clk cell_8740 ( .C (clk), .D (signal_11285), .Q (signal_11286) ) ;
    buf_clk cell_8756 ( .C (clk), .D (signal_11301), .Q (signal_11302) ) ;
    buf_clk cell_8772 ( .C (clk), .D (signal_11317), .Q (signal_11318) ) ;
    buf_clk cell_8788 ( .C (clk), .D (signal_11333), .Q (signal_11334) ) ;
    buf_clk cell_8804 ( .C (clk), .D (signal_11349), .Q (signal_11350) ) ;
    buf_clk cell_8820 ( .C (clk), .D (signal_11365), .Q (signal_11366) ) ;
    buf_clk cell_8836 ( .C (clk), .D (signal_11381), .Q (signal_11382) ) ;
    buf_clk cell_8852 ( .C (clk), .D (signal_11397), .Q (signal_11398) ) ;
    buf_clk cell_8868 ( .C (clk), .D (signal_11413), .Q (signal_11414) ) ;
    buf_clk cell_8884 ( .C (clk), .D (signal_11429), .Q (signal_11430) ) ;
    buf_clk cell_8900 ( .C (clk), .D (signal_11445), .Q (signal_11446) ) ;
    buf_clk cell_8916 ( .C (clk), .D (signal_11461), .Q (signal_11462) ) ;
    buf_clk cell_8932 ( .C (clk), .D (signal_11477), .Q (signal_11478) ) ;
    buf_clk cell_8948 ( .C (clk), .D (signal_11493), .Q (signal_11494) ) ;
    buf_clk cell_8964 ( .C (clk), .D (signal_11509), .Q (signal_11510) ) ;
    buf_clk cell_8980 ( .C (clk), .D (signal_11525), .Q (signal_11526) ) ;
    buf_clk cell_8996 ( .C (clk), .D (signal_11541), .Q (signal_11542) ) ;
    buf_clk cell_9012 ( .C (clk), .D (signal_11557), .Q (signal_11558) ) ;
    buf_clk cell_9028 ( .C (clk), .D (signal_11573), .Q (signal_11574) ) ;
    buf_clk cell_9044 ( .C (clk), .D (signal_11589), .Q (signal_11590) ) ;
    buf_clk cell_9060 ( .C (clk), .D (signal_11605), .Q (signal_11606) ) ;
    buf_clk cell_9076 ( .C (clk), .D (signal_11621), .Q (signal_11622) ) ;
    buf_clk cell_9092 ( .C (clk), .D (signal_11637), .Q (signal_11638) ) ;
    buf_clk cell_9108 ( .C (clk), .D (signal_11653), .Q (signal_11654) ) ;
    buf_clk cell_9124 ( .C (clk), .D (signal_11669), .Q (signal_11670) ) ;
    buf_clk cell_9140 ( .C (clk), .D (signal_11685), .Q (signal_11686) ) ;
    buf_clk cell_9156 ( .C (clk), .D (signal_11701), .Q (signal_11702) ) ;
    buf_clk cell_9172 ( .C (clk), .D (signal_11717), .Q (signal_11718) ) ;
    buf_clk cell_9188 ( .C (clk), .D (signal_11733), .Q (signal_11734) ) ;
    buf_clk cell_9204 ( .C (clk), .D (signal_11749), .Q (signal_11750) ) ;
    buf_clk cell_9220 ( .C (clk), .D (signal_11765), .Q (signal_11766) ) ;
    buf_clk cell_9236 ( .C (clk), .D (signal_11781), .Q (signal_11782) ) ;
    buf_clk cell_9252 ( .C (clk), .D (signal_11797), .Q (signal_11798) ) ;
    buf_clk cell_9268 ( .C (clk), .D (signal_11813), .Q (signal_11814) ) ;
    buf_clk cell_9284 ( .C (clk), .D (signal_11829), .Q (signal_11830) ) ;
    buf_clk cell_9300 ( .C (clk), .D (signal_11845), .Q (signal_11846) ) ;
    buf_clk cell_9316 ( .C (clk), .D (signal_11861), .Q (signal_11862) ) ;
    buf_clk cell_9332 ( .C (clk), .D (signal_11877), .Q (signal_11878) ) ;
    buf_clk cell_9348 ( .C (clk), .D (signal_11893), .Q (signal_11894) ) ;
    buf_clk cell_9364 ( .C (clk), .D (signal_11909), .Q (signal_11910) ) ;
    buf_clk cell_9380 ( .C (clk), .D (signal_11925), .Q (signal_11926) ) ;
    buf_clk cell_9396 ( .C (clk), .D (signal_11941), .Q (signal_11942) ) ;
    buf_clk cell_9412 ( .C (clk), .D (signal_11957), .Q (signal_11958) ) ;
    buf_clk cell_9428 ( .C (clk), .D (signal_11973), .Q (signal_11974) ) ;
    buf_clk cell_9444 ( .C (clk), .D (signal_11989), .Q (signal_11990) ) ;
    buf_clk cell_9460 ( .C (clk), .D (signal_12005), .Q (signal_12006) ) ;
    buf_clk cell_9476 ( .C (clk), .D (signal_12021), .Q (signal_12022) ) ;
    buf_clk cell_9492 ( .C (clk), .D (signal_12037), .Q (signal_12038) ) ;
    buf_clk cell_9508 ( .C (clk), .D (signal_12053), .Q (signal_12054) ) ;
    buf_clk cell_9524 ( .C (clk), .D (signal_12069), .Q (signal_12070) ) ;
    buf_clk cell_9540 ( .C (clk), .D (signal_12085), .Q (signal_12086) ) ;
    buf_clk cell_9556 ( .C (clk), .D (signal_12101), .Q (signal_12102) ) ;
    buf_clk cell_9572 ( .C (clk), .D (signal_12117), .Q (signal_12118) ) ;
    buf_clk cell_9588 ( .C (clk), .D (signal_12133), .Q (signal_12134) ) ;
    buf_clk cell_9604 ( .C (clk), .D (signal_12149), .Q (signal_12150) ) ;
    buf_clk cell_9620 ( .C (clk), .D (signal_12165), .Q (signal_12166) ) ;
    buf_clk cell_9636 ( .C (clk), .D (signal_12181), .Q (signal_12182) ) ;
    buf_clk cell_9652 ( .C (clk), .D (signal_12197), .Q (signal_12198) ) ;
    buf_clk cell_9668 ( .C (clk), .D (signal_12213), .Q (signal_12214) ) ;
    buf_clk cell_9684 ( .C (clk), .D (signal_12229), .Q (signal_12230) ) ;
    buf_clk cell_9700 ( .C (clk), .D (signal_12245), .Q (signal_12246) ) ;
    buf_clk cell_9716 ( .C (clk), .D (signal_12261), .Q (signal_12262) ) ;
    buf_clk cell_9732 ( .C (clk), .D (signal_12277), .Q (signal_12278) ) ;
    buf_clk cell_9748 ( .C (clk), .D (signal_12293), .Q (signal_12294) ) ;
    buf_clk cell_9764 ( .C (clk), .D (signal_12309), .Q (signal_12310) ) ;
    buf_clk cell_9780 ( .C (clk), .D (signal_12325), .Q (signal_12326) ) ;
    buf_clk cell_9796 ( .C (clk), .D (signal_12341), .Q (signal_12342) ) ;
    buf_clk cell_9812 ( .C (clk), .D (signal_12357), .Q (signal_12358) ) ;
    buf_clk cell_9828 ( .C (clk), .D (signal_12373), .Q (signal_12374) ) ;
    buf_clk cell_9844 ( .C (clk), .D (signal_12389), .Q (signal_12390) ) ;
    buf_clk cell_9860 ( .C (clk), .D (signal_12405), .Q (signal_12406) ) ;
    buf_clk cell_9876 ( .C (clk), .D (signal_12421), .Q (signal_12422) ) ;
    buf_clk cell_9892 ( .C (clk), .D (signal_12437), .Q (signal_12438) ) ;
    buf_clk cell_9908 ( .C (clk), .D (signal_12453), .Q (signal_12454) ) ;
    buf_clk cell_9924 ( .C (clk), .D (signal_12469), .Q (signal_12470) ) ;
    buf_clk cell_9940 ( .C (clk), .D (signal_12485), .Q (signal_12486) ) ;
    buf_clk cell_9956 ( .C (clk), .D (signal_12501), .Q (signal_12502) ) ;
    buf_clk cell_9972 ( .C (clk), .D (signal_12517), .Q (signal_12518) ) ;
    buf_clk cell_9988 ( .C (clk), .D (signal_12533), .Q (signal_12534) ) ;
    buf_clk cell_10004 ( .C (clk), .D (signal_12549), .Q (signal_12550) ) ;
    buf_clk cell_10020 ( .C (clk), .D (signal_12565), .Q (signal_12566) ) ;
    buf_clk cell_10036 ( .C (clk), .D (signal_12581), .Q (signal_12582) ) ;
    buf_clk cell_10052 ( .C (clk), .D (signal_12597), .Q (signal_12598) ) ;
    buf_clk cell_10068 ( .C (clk), .D (signal_12613), .Q (signal_12614) ) ;
    buf_clk cell_10084 ( .C (clk), .D (signal_12629), .Q (signal_12630) ) ;
    buf_clk cell_10100 ( .C (clk), .D (signal_12645), .Q (signal_12646) ) ;
    buf_clk cell_10116 ( .C (clk), .D (signal_12661), .Q (signal_12662) ) ;
    buf_clk cell_10132 ( .C (clk), .D (signal_12677), .Q (signal_12678) ) ;
    buf_clk cell_10148 ( .C (clk), .D (signal_12693), .Q (signal_12694) ) ;
    buf_clk cell_10164 ( .C (clk), .D (signal_12709), .Q (signal_12710) ) ;
    buf_clk cell_10180 ( .C (clk), .D (signal_12725), .Q (signal_12726) ) ;
    buf_clk cell_10196 ( .C (clk), .D (signal_12741), .Q (signal_12742) ) ;
    buf_clk cell_10212 ( .C (clk), .D (signal_12757), .Q (signal_12758) ) ;
    buf_clk cell_10228 ( .C (clk), .D (signal_12773), .Q (signal_12774) ) ;
    buf_clk cell_10244 ( .C (clk), .D (signal_12789), .Q (signal_12790) ) ;
    buf_clk cell_10260 ( .C (clk), .D (signal_12805), .Q (signal_12806) ) ;
    buf_clk cell_10276 ( .C (clk), .D (signal_12821), .Q (signal_12822) ) ;
    buf_clk cell_10292 ( .C (clk), .D (signal_12837), .Q (signal_12838) ) ;
    buf_clk cell_10308 ( .C (clk), .D (signal_12853), .Q (signal_12854) ) ;
    buf_clk cell_10324 ( .C (clk), .D (signal_12869), .Q (signal_12870) ) ;
    buf_clk cell_10340 ( .C (clk), .D (signal_12885), .Q (signal_12886) ) ;
    buf_clk cell_10356 ( .C (clk), .D (signal_12901), .Q (signal_12902) ) ;
    buf_clk cell_10372 ( .C (clk), .D (signal_12917), .Q (signal_12918) ) ;
    buf_clk cell_10388 ( .C (clk), .D (signal_12933), .Q (signal_12934) ) ;
    buf_clk cell_10404 ( .C (clk), .D (signal_12949), .Q (signal_12950) ) ;
    buf_clk cell_10420 ( .C (clk), .D (signal_12965), .Q (signal_12966) ) ;
    buf_clk cell_10436 ( .C (clk), .D (signal_12981), .Q (signal_12982) ) ;
    buf_clk cell_10452 ( .C (clk), .D (signal_12997), .Q (signal_12998) ) ;
    buf_clk cell_10468 ( .C (clk), .D (signal_13013), .Q (signal_13014) ) ;
    buf_clk cell_10484 ( .C (clk), .D (signal_13029), .Q (signal_13030) ) ;
    buf_clk cell_10500 ( .C (clk), .D (signal_13045), .Q (signal_13046) ) ;
    buf_clk cell_10516 ( .C (clk), .D (signal_13061), .Q (signal_13062) ) ;
    buf_clk cell_10532 ( .C (clk), .D (signal_13077), .Q (signal_13078) ) ;
    buf_clk cell_10548 ( .C (clk), .D (signal_13093), .Q (signal_13094) ) ;
    buf_clk cell_10564 ( .C (clk), .D (signal_13109), .Q (signal_13110) ) ;
    buf_clk cell_10580 ( .C (clk), .D (signal_13125), .Q (signal_13126) ) ;
    buf_clk cell_10596 ( .C (clk), .D (signal_13141), .Q (signal_13142) ) ;
    buf_clk cell_10612 ( .C (clk), .D (signal_13157), .Q (signal_13158) ) ;
    buf_clk cell_10628 ( .C (clk), .D (signal_13173), .Q (signal_13174) ) ;
    buf_clk cell_10644 ( .C (clk), .D (signal_13189), .Q (signal_13190) ) ;
    buf_clk cell_10660 ( .C (clk), .D (signal_13205), .Q (signal_13206) ) ;
    buf_clk cell_10676 ( .C (clk), .D (signal_13221), .Q (signal_13222) ) ;
    buf_clk cell_10692 ( .C (clk), .D (signal_13237), .Q (signal_13238) ) ;
    buf_clk cell_10708 ( .C (clk), .D (signal_13253), .Q (signal_13254) ) ;
    buf_clk cell_10724 ( .C (clk), .D (signal_13269), .Q (signal_13270) ) ;
    buf_clk cell_10740 ( .C (clk), .D (signal_13285), .Q (signal_13286) ) ;
    buf_clk cell_10756 ( .C (clk), .D (signal_13301), .Q (signal_13302) ) ;
    buf_clk cell_10772 ( .C (clk), .D (signal_13317), .Q (signal_13318) ) ;
    buf_clk cell_10788 ( .C (clk), .D (signal_13333), .Q (signal_13334) ) ;
    buf_clk cell_10804 ( .C (clk), .D (signal_13349), .Q (signal_13350) ) ;
    buf_clk cell_10820 ( .C (clk), .D (signal_13365), .Q (signal_13366) ) ;
    buf_clk cell_10836 ( .C (clk), .D (signal_13381), .Q (signal_13382) ) ;
    buf_clk cell_10852 ( .C (clk), .D (signal_13397), .Q (signal_13398) ) ;
    buf_clk cell_10868 ( .C (clk), .D (signal_13413), .Q (signal_13414) ) ;
    buf_clk cell_10884 ( .C (clk), .D (signal_13429), .Q (signal_13430) ) ;
    buf_clk cell_10900 ( .C (clk), .D (signal_13445), .Q (signal_13446) ) ;
    buf_clk cell_10916 ( .C (clk), .D (signal_13461), .Q (signal_13462) ) ;
    buf_clk cell_10932 ( .C (clk), .D (signal_13477), .Q (signal_13478) ) ;
    buf_clk cell_10948 ( .C (clk), .D (signal_13493), .Q (signal_13494) ) ;
    buf_clk cell_10964 ( .C (clk), .D (signal_13509), .Q (signal_13510) ) ;
    buf_clk cell_10980 ( .C (clk), .D (signal_13525), .Q (signal_13526) ) ;
    buf_clk cell_10996 ( .C (clk), .D (signal_13541), .Q (signal_13542) ) ;
    buf_clk cell_11012 ( .C (clk), .D (signal_13557), .Q (signal_13558) ) ;
    buf_clk cell_11028 ( .C (clk), .D (signal_13573), .Q (signal_13574) ) ;
    buf_clk cell_11044 ( .C (clk), .D (signal_13589), .Q (signal_13590) ) ;
    buf_clk cell_11060 ( .C (clk), .D (signal_13605), .Q (signal_13606) ) ;
    buf_clk cell_11076 ( .C (clk), .D (signal_13621), .Q (signal_13622) ) ;
    buf_clk cell_11092 ( .C (clk), .D (signal_13637), .Q (signal_13638) ) ;
    buf_clk cell_11108 ( .C (clk), .D (signal_13653), .Q (signal_13654) ) ;
    buf_clk cell_11124 ( .C (clk), .D (signal_13669), .Q (signal_13670) ) ;
    buf_clk cell_11140 ( .C (clk), .D (signal_13685), .Q (signal_13686) ) ;
    buf_clk cell_11156 ( .C (clk), .D (signal_13701), .Q (signal_13702) ) ;
    buf_clk cell_11172 ( .C (clk), .D (signal_13717), .Q (signal_13718) ) ;
    buf_clk cell_11188 ( .C (clk), .D (signal_13733), .Q (signal_13734) ) ;
    buf_clk cell_11204 ( .C (clk), .D (signal_13749), .Q (signal_13750) ) ;
    buf_clk cell_11220 ( .C (clk), .D (signal_13765), .Q (signal_13766) ) ;
    buf_clk cell_11236 ( .C (clk), .D (signal_13781), .Q (signal_13782) ) ;
    buf_clk cell_11252 ( .C (clk), .D (signal_13797), .Q (signal_13798) ) ;
    buf_clk cell_11268 ( .C (clk), .D (signal_13813), .Q (signal_13814) ) ;
    buf_clk cell_11284 ( .C (clk), .D (signal_13829), .Q (signal_13830) ) ;
    buf_clk cell_11300 ( .C (clk), .D (signal_13845), .Q (signal_13846) ) ;
    buf_clk cell_11316 ( .C (clk), .D (signal_13861), .Q (signal_13862) ) ;
    buf_clk cell_11332 ( .C (clk), .D (signal_13877), .Q (signal_13878) ) ;
    buf_clk cell_11348 ( .C (clk), .D (signal_13893), .Q (signal_13894) ) ;
    buf_clk cell_11364 ( .C (clk), .D (signal_13909), .Q (signal_13910) ) ;
    buf_clk cell_11380 ( .C (clk), .D (signal_13925), .Q (signal_13926) ) ;
    buf_clk cell_11396 ( .C (clk), .D (signal_13941), .Q (signal_13942) ) ;
    buf_clk cell_11412 ( .C (clk), .D (signal_13957), .Q (signal_13958) ) ;
    buf_clk cell_11428 ( .C (clk), .D (signal_13973), .Q (signal_13974) ) ;
    buf_clk cell_11444 ( .C (clk), .D (signal_13989), .Q (signal_13990) ) ;
    buf_clk cell_11460 ( .C (clk), .D (signal_14005), .Q (signal_14006) ) ;
    buf_clk cell_11476 ( .C (clk), .D (signal_14021), .Q (signal_14022) ) ;
    buf_clk cell_11492 ( .C (clk), .D (signal_14037), .Q (signal_14038) ) ;
    buf_clk cell_11508 ( .C (clk), .D (signal_14053), .Q (signal_14054) ) ;
    buf_clk cell_11524 ( .C (clk), .D (signal_14069), .Q (signal_14070) ) ;
    buf_clk cell_11540 ( .C (clk), .D (signal_14085), .Q (signal_14086) ) ;
    buf_clk cell_11556 ( .C (clk), .D (signal_14101), .Q (signal_14102) ) ;
    buf_clk cell_11572 ( .C (clk), .D (signal_14117), .Q (signal_14118) ) ;
    buf_clk cell_11588 ( .C (clk), .D (signal_14133), .Q (signal_14134) ) ;
    buf_clk cell_11604 ( .C (clk), .D (signal_14149), .Q (signal_14150) ) ;
    buf_clk cell_11620 ( .C (clk), .D (signal_14165), .Q (signal_14166) ) ;
    buf_clk cell_11636 ( .C (clk), .D (signal_14181), .Q (signal_14182) ) ;
    buf_clk cell_11652 ( .C (clk), .D (signal_14197), .Q (signal_14198) ) ;
    buf_clk cell_11668 ( .C (clk), .D (signal_14213), .Q (signal_14214) ) ;
    buf_clk cell_11684 ( .C (clk), .D (signal_14229), .Q (signal_14230) ) ;
    buf_clk cell_11700 ( .C (clk), .D (signal_14245), .Q (signal_14246) ) ;
    buf_clk cell_11716 ( .C (clk), .D (signal_14261), .Q (signal_14262) ) ;
    buf_clk cell_11732 ( .C (clk), .D (signal_14277), .Q (signal_14278) ) ;
    buf_clk cell_11748 ( .C (clk), .D (signal_14293), .Q (signal_14294) ) ;
    buf_clk cell_11764 ( .C (clk), .D (signal_14309), .Q (signal_14310) ) ;
    buf_clk cell_11780 ( .C (clk), .D (signal_14325), .Q (signal_14326) ) ;
    buf_clk cell_11796 ( .C (clk), .D (signal_14341), .Q (signal_14342) ) ;
    buf_clk cell_11812 ( .C (clk), .D (signal_14357), .Q (signal_14358) ) ;
    buf_clk cell_11828 ( .C (clk), .D (signal_14373), .Q (signal_14374) ) ;
    buf_clk cell_11844 ( .C (clk), .D (signal_14389), .Q (signal_14390) ) ;
    buf_clk cell_11860 ( .C (clk), .D (signal_14405), .Q (signal_14406) ) ;
    buf_clk cell_11876 ( .C (clk), .D (signal_14421), .Q (signal_14422) ) ;
    buf_clk cell_11892 ( .C (clk), .D (signal_14437), .Q (signal_14438) ) ;
    buf_clk cell_11908 ( .C (clk), .D (signal_14453), .Q (signal_14454) ) ;
    buf_clk cell_11924 ( .C (clk), .D (signal_14469), .Q (signal_14470) ) ;
    buf_clk cell_11940 ( .C (clk), .D (signal_14485), .Q (signal_14486) ) ;
    buf_clk cell_11956 ( .C (clk), .D (signal_14501), .Q (signal_14502) ) ;
    buf_clk cell_11972 ( .C (clk), .D (signal_14517), .Q (signal_14518) ) ;
    buf_clk cell_11988 ( .C (clk), .D (signal_14533), .Q (signal_14534) ) ;
    buf_clk cell_12004 ( .C (clk), .D (signal_14549), .Q (signal_14550) ) ;
    buf_clk cell_12020 ( .C (clk), .D (signal_14565), .Q (signal_14566) ) ;
    buf_clk cell_12036 ( .C (clk), .D (signal_14581), .Q (signal_14582) ) ;
    buf_clk cell_12052 ( .C (clk), .D (signal_14597), .Q (signal_14598) ) ;
    buf_clk cell_12068 ( .C (clk), .D (signal_14613), .Q (signal_14614) ) ;
    buf_clk cell_12084 ( .C (clk), .D (signal_14629), .Q (signal_14630) ) ;
    buf_clk cell_12100 ( .C (clk), .D (signal_14645), .Q (signal_14646) ) ;
    buf_clk cell_12116 ( .C (clk), .D (signal_14661), .Q (signal_14662) ) ;
    buf_clk cell_12132 ( .C (clk), .D (signal_14677), .Q (signal_14678) ) ;
    buf_clk cell_12148 ( .C (clk), .D (signal_14693), .Q (signal_14694) ) ;
    buf_clk cell_12164 ( .C (clk), .D (signal_14709), .Q (signal_14710) ) ;
    buf_clk cell_12180 ( .C (clk), .D (signal_14725), .Q (signal_14726) ) ;
    buf_clk cell_12196 ( .C (clk), .D (signal_14741), .Q (signal_14742) ) ;
    buf_clk cell_12212 ( .C (clk), .D (signal_14757), .Q (signal_14758) ) ;
    buf_clk cell_12228 ( .C (clk), .D (signal_14773), .Q (signal_14774) ) ;
    buf_clk cell_12244 ( .C (clk), .D (signal_14789), .Q (signal_14790) ) ;
    buf_clk cell_12260 ( .C (clk), .D (signal_14805), .Q (signal_14806) ) ;
    buf_clk cell_12276 ( .C (clk), .D (signal_14821), .Q (signal_14822) ) ;
    buf_clk cell_12292 ( .C (clk), .D (signal_14837), .Q (signal_14838) ) ;
    buf_clk cell_12308 ( .C (clk), .D (signal_14853), .Q (signal_14854) ) ;
    buf_clk cell_12324 ( .C (clk), .D (signal_14869), .Q (signal_14870) ) ;
    buf_clk cell_12340 ( .C (clk), .D (signal_14885), .Q (signal_14886) ) ;
    buf_clk cell_12356 ( .C (clk), .D (signal_14901), .Q (signal_14902) ) ;
    buf_clk cell_12372 ( .C (clk), .D (signal_14917), .Q (signal_14918) ) ;
    buf_clk cell_12388 ( .C (clk), .D (signal_14933), .Q (signal_14934) ) ;

    /* cells in depth 9 */
    buf_clk cell_2349 ( .C (clk), .D (signal_4894), .Q (signal_4895) ) ;
    buf_clk cell_2359 ( .C (clk), .D (signal_4904), .Q (signal_4905) ) ;
    buf_clk cell_2369 ( .C (clk), .D (signal_4914), .Q (signal_4915) ) ;
    buf_clk cell_2381 ( .C (clk), .D (signal_4926), .Q (signal_4927) ) ;
    buf_clk cell_2393 ( .C (clk), .D (signal_4938), .Q (signal_4939) ) ;
    buf_clk cell_2409 ( .C (clk), .D (signal_4954), .Q (signal_4955) ) ;
    buf_clk cell_2425 ( .C (clk), .D (signal_4970), .Q (signal_4971) ) ;
    buf_clk cell_2441 ( .C (clk), .D (signal_4986), .Q (signal_4987) ) ;
    buf_clk cell_2457 ( .C (clk), .D (signal_5002), .Q (signal_5003) ) ;
    buf_clk cell_2473 ( .C (clk), .D (signal_5018), .Q (signal_5019) ) ;
    buf_clk cell_2489 ( .C (clk), .D (signal_5034), .Q (signal_5035) ) ;
    buf_clk cell_2505 ( .C (clk), .D (signal_5050), .Q (signal_5051) ) ;
    buf_clk cell_2521 ( .C (clk), .D (signal_5066), .Q (signal_5067) ) ;
    buf_clk cell_2537 ( .C (clk), .D (signal_5082), .Q (signal_5083) ) ;
    buf_clk cell_2553 ( .C (clk), .D (signal_5098), .Q (signal_5099) ) ;
    buf_clk cell_2569 ( .C (clk), .D (signal_5114), .Q (signal_5115) ) ;
    buf_clk cell_2585 ( .C (clk), .D (signal_5130), .Q (signal_5131) ) ;
    buf_clk cell_2601 ( .C (clk), .D (signal_5146), .Q (signal_5147) ) ;
    buf_clk cell_2617 ( .C (clk), .D (signal_5162), .Q (signal_5163) ) ;
    buf_clk cell_2633 ( .C (clk), .D (signal_5178), .Q (signal_5179) ) ;
    buf_clk cell_2649 ( .C (clk), .D (signal_5194), .Q (signal_5195) ) ;
    buf_clk cell_2665 ( .C (clk), .D (signal_5210), .Q (signal_5211) ) ;
    buf_clk cell_2681 ( .C (clk), .D (signal_5226), .Q (signal_5227) ) ;
    buf_clk cell_2697 ( .C (clk), .D (signal_5242), .Q (signal_5243) ) ;
    buf_clk cell_2713 ( .C (clk), .D (signal_5258), .Q (signal_5259) ) ;
    buf_clk cell_2729 ( .C (clk), .D (signal_5274), .Q (signal_5275) ) ;
    buf_clk cell_2745 ( .C (clk), .D (signal_5290), .Q (signal_5291) ) ;
    buf_clk cell_2761 ( .C (clk), .D (signal_5306), .Q (signal_5307) ) ;
    buf_clk cell_2777 ( .C (clk), .D (signal_5322), .Q (signal_5323) ) ;
    buf_clk cell_2793 ( .C (clk), .D (signal_5338), .Q (signal_5339) ) ;
    buf_clk cell_2809 ( .C (clk), .D (signal_5354), .Q (signal_5355) ) ;
    buf_clk cell_2825 ( .C (clk), .D (signal_5370), .Q (signal_5371) ) ;
    buf_clk cell_2841 ( .C (clk), .D (signal_5386), .Q (signal_5387) ) ;
    buf_clk cell_2857 ( .C (clk), .D (signal_5402), .Q (signal_5403) ) ;
    buf_clk cell_2873 ( .C (clk), .D (signal_5418), .Q (signal_5419) ) ;
    buf_clk cell_2889 ( .C (clk), .D (signal_5434), .Q (signal_5435) ) ;
    buf_clk cell_2905 ( .C (clk), .D (signal_5450), .Q (signal_5451) ) ;
    buf_clk cell_2921 ( .C (clk), .D (signal_5466), .Q (signal_5467) ) ;
    buf_clk cell_2937 ( .C (clk), .D (signal_5482), .Q (signal_5483) ) ;
    buf_clk cell_2953 ( .C (clk), .D (signal_5498), .Q (signal_5499) ) ;
    buf_clk cell_2969 ( .C (clk), .D (signal_5514), .Q (signal_5515) ) ;
    buf_clk cell_2985 ( .C (clk), .D (signal_5530), .Q (signal_5531) ) ;
    buf_clk cell_3001 ( .C (clk), .D (signal_5546), .Q (signal_5547) ) ;
    buf_clk cell_3017 ( .C (clk), .D (signal_5562), .Q (signal_5563) ) ;
    buf_clk cell_3033 ( .C (clk), .D (signal_5578), .Q (signal_5579) ) ;
    buf_clk cell_3049 ( .C (clk), .D (signal_5594), .Q (signal_5595) ) ;
    buf_clk cell_3065 ( .C (clk), .D (signal_5610), .Q (signal_5611) ) ;
    buf_clk cell_3081 ( .C (clk), .D (signal_5626), .Q (signal_5627) ) ;
    buf_clk cell_3097 ( .C (clk), .D (signal_5642), .Q (signal_5643) ) ;
    buf_clk cell_3113 ( .C (clk), .D (signal_5658), .Q (signal_5659) ) ;
    buf_clk cell_3129 ( .C (clk), .D (signal_5674), .Q (signal_5675) ) ;
    buf_clk cell_3145 ( .C (clk), .D (signal_5690), .Q (signal_5691) ) ;
    buf_clk cell_3161 ( .C (clk), .D (signal_5706), .Q (signal_5707) ) ;
    buf_clk cell_3177 ( .C (clk), .D (signal_5722), .Q (signal_5723) ) ;
    buf_clk cell_3193 ( .C (clk), .D (signal_5738), .Q (signal_5739) ) ;
    buf_clk cell_3209 ( .C (clk), .D (signal_5754), .Q (signal_5755) ) ;
    buf_clk cell_3225 ( .C (clk), .D (signal_5770), .Q (signal_5771) ) ;
    buf_clk cell_3241 ( .C (clk), .D (signal_5786), .Q (signal_5787) ) ;
    buf_clk cell_3257 ( .C (clk), .D (signal_5802), .Q (signal_5803) ) ;
    buf_clk cell_3273 ( .C (clk), .D (signal_5818), .Q (signal_5819) ) ;
    buf_clk cell_3289 ( .C (clk), .D (signal_5834), .Q (signal_5835) ) ;
    buf_clk cell_3305 ( .C (clk), .D (signal_5850), .Q (signal_5851) ) ;
    buf_clk cell_3321 ( .C (clk), .D (signal_5866), .Q (signal_5867) ) ;
    buf_clk cell_3337 ( .C (clk), .D (signal_5882), .Q (signal_5883) ) ;
    buf_clk cell_3353 ( .C (clk), .D (signal_5898), .Q (signal_5899) ) ;
    buf_clk cell_3369 ( .C (clk), .D (signal_5914), .Q (signal_5915) ) ;
    buf_clk cell_3385 ( .C (clk), .D (signal_5930), .Q (signal_5931) ) ;
    buf_clk cell_3401 ( .C (clk), .D (signal_5946), .Q (signal_5947) ) ;
    buf_clk cell_3417 ( .C (clk), .D (signal_5962), .Q (signal_5963) ) ;
    buf_clk cell_3433 ( .C (clk), .D (signal_5978), .Q (signal_5979) ) ;
    buf_clk cell_3449 ( .C (clk), .D (signal_5994), .Q (signal_5995) ) ;
    buf_clk cell_3465 ( .C (clk), .D (signal_6010), .Q (signal_6011) ) ;
    buf_clk cell_3481 ( .C (clk), .D (signal_6026), .Q (signal_6027) ) ;
    buf_clk cell_3497 ( .C (clk), .D (signal_6042), .Q (signal_6043) ) ;
    buf_clk cell_3513 ( .C (clk), .D (signal_6058), .Q (signal_6059) ) ;
    buf_clk cell_3529 ( .C (clk), .D (signal_6074), .Q (signal_6075) ) ;
    buf_clk cell_3545 ( .C (clk), .D (signal_6090), .Q (signal_6091) ) ;
    buf_clk cell_3561 ( .C (clk), .D (signal_6106), .Q (signal_6107) ) ;
    buf_clk cell_3577 ( .C (clk), .D (signal_6122), .Q (signal_6123) ) ;
    buf_clk cell_3593 ( .C (clk), .D (signal_6138), .Q (signal_6139) ) ;
    buf_clk cell_3609 ( .C (clk), .D (signal_6154), .Q (signal_6155) ) ;
    buf_clk cell_3625 ( .C (clk), .D (signal_6170), .Q (signal_6171) ) ;
    buf_clk cell_3641 ( .C (clk), .D (signal_6186), .Q (signal_6187) ) ;
    buf_clk cell_3657 ( .C (clk), .D (signal_6202), .Q (signal_6203) ) ;
    buf_clk cell_3673 ( .C (clk), .D (signal_6218), .Q (signal_6219) ) ;
    buf_clk cell_3689 ( .C (clk), .D (signal_6234), .Q (signal_6235) ) ;
    buf_clk cell_3705 ( .C (clk), .D (signal_6250), .Q (signal_6251) ) ;
    buf_clk cell_3721 ( .C (clk), .D (signal_6266), .Q (signal_6267) ) ;
    buf_clk cell_3737 ( .C (clk), .D (signal_6282), .Q (signal_6283) ) ;
    buf_clk cell_3753 ( .C (clk), .D (signal_6298), .Q (signal_6299) ) ;
    buf_clk cell_3769 ( .C (clk), .D (signal_6314), .Q (signal_6315) ) ;
    buf_clk cell_3785 ( .C (clk), .D (signal_6330), .Q (signal_6331) ) ;
    buf_clk cell_3801 ( .C (clk), .D (signal_6346), .Q (signal_6347) ) ;
    buf_clk cell_3817 ( .C (clk), .D (signal_6362), .Q (signal_6363) ) ;
    buf_clk cell_3833 ( .C (clk), .D (signal_6378), .Q (signal_6379) ) ;
    buf_clk cell_3849 ( .C (clk), .D (signal_6394), .Q (signal_6395) ) ;
    buf_clk cell_3865 ( .C (clk), .D (signal_6410), .Q (signal_6411) ) ;
    buf_clk cell_3881 ( .C (clk), .D (signal_6426), .Q (signal_6427) ) ;
    buf_clk cell_3897 ( .C (clk), .D (signal_6442), .Q (signal_6443) ) ;
    buf_clk cell_3913 ( .C (clk), .D (signal_6458), .Q (signal_6459) ) ;
    buf_clk cell_3929 ( .C (clk), .D (signal_6474), .Q (signal_6475) ) ;
    buf_clk cell_3945 ( .C (clk), .D (signal_6490), .Q (signal_6491) ) ;
    buf_clk cell_3961 ( .C (clk), .D (signal_6506), .Q (signal_6507) ) ;
    buf_clk cell_3977 ( .C (clk), .D (signal_6522), .Q (signal_6523) ) ;
    buf_clk cell_3993 ( .C (clk), .D (signal_6538), .Q (signal_6539) ) ;
    buf_clk cell_4009 ( .C (clk), .D (signal_6554), .Q (signal_6555) ) ;
    buf_clk cell_4025 ( .C (clk), .D (signal_6570), .Q (signal_6571) ) ;
    buf_clk cell_4041 ( .C (clk), .D (signal_6586), .Q (signal_6587) ) ;
    buf_clk cell_4057 ( .C (clk), .D (signal_6602), .Q (signal_6603) ) ;
    buf_clk cell_4073 ( .C (clk), .D (signal_6618), .Q (signal_6619) ) ;
    buf_clk cell_4089 ( .C (clk), .D (signal_6634), .Q (signal_6635) ) ;
    buf_clk cell_4105 ( .C (clk), .D (signal_6650), .Q (signal_6651) ) ;
    buf_clk cell_4121 ( .C (clk), .D (signal_6666), .Q (signal_6667) ) ;
    buf_clk cell_4137 ( .C (clk), .D (signal_6682), .Q (signal_6683) ) ;
    buf_clk cell_4153 ( .C (clk), .D (signal_6698), .Q (signal_6699) ) ;
    buf_clk cell_4169 ( .C (clk), .D (signal_6714), .Q (signal_6715) ) ;
    buf_clk cell_4185 ( .C (clk), .D (signal_6730), .Q (signal_6731) ) ;
    buf_clk cell_4201 ( .C (clk), .D (signal_6746), .Q (signal_6747) ) ;
    buf_clk cell_4217 ( .C (clk), .D (signal_6762), .Q (signal_6763) ) ;
    buf_clk cell_4233 ( .C (clk), .D (signal_6778), .Q (signal_6779) ) ;
    buf_clk cell_4249 ( .C (clk), .D (signal_6794), .Q (signal_6795) ) ;
    buf_clk cell_4265 ( .C (clk), .D (signal_6810), .Q (signal_6811) ) ;
    buf_clk cell_4281 ( .C (clk), .D (signal_6826), .Q (signal_6827) ) ;
    buf_clk cell_4297 ( .C (clk), .D (signal_6842), .Q (signal_6843) ) ;
    buf_clk cell_4313 ( .C (clk), .D (signal_6858), .Q (signal_6859) ) ;
    buf_clk cell_4329 ( .C (clk), .D (signal_6874), .Q (signal_6875) ) ;
    buf_clk cell_4345 ( .C (clk), .D (signal_6890), .Q (signal_6891) ) ;
    buf_clk cell_4361 ( .C (clk), .D (signal_6906), .Q (signal_6907) ) ;
    buf_clk cell_4377 ( .C (clk), .D (signal_6922), .Q (signal_6923) ) ;
    buf_clk cell_4393 ( .C (clk), .D (signal_6938), .Q (signal_6939) ) ;
    buf_clk cell_4409 ( .C (clk), .D (signal_6954), .Q (signal_6955) ) ;
    buf_clk cell_4423 ( .C (clk), .D (signal_6968), .Q (signal_6969) ) ;
    buf_clk cell_4437 ( .C (clk), .D (signal_6982), .Q (signal_6983) ) ;
    buf_clk cell_4453 ( .C (clk), .D (signal_6998), .Q (signal_6999) ) ;
    buf_clk cell_4469 ( .C (clk), .D (signal_7014), .Q (signal_7015) ) ;
    buf_clk cell_4485 ( .C (clk), .D (signal_7030), .Q (signal_7031) ) ;
    buf_clk cell_4501 ( .C (clk), .D (signal_7046), .Q (signal_7047) ) ;
    buf_clk cell_4517 ( .C (clk), .D (signal_7062), .Q (signal_7063) ) ;
    buf_clk cell_4533 ( .C (clk), .D (signal_7078), .Q (signal_7079) ) ;
    buf_clk cell_4549 ( .C (clk), .D (signal_7094), .Q (signal_7095) ) ;
    buf_clk cell_4565 ( .C (clk), .D (signal_7110), .Q (signal_7111) ) ;
    buf_clk cell_4581 ( .C (clk), .D (signal_7126), .Q (signal_7127) ) ;
    buf_clk cell_4597 ( .C (clk), .D (signal_7142), .Q (signal_7143) ) ;
    buf_clk cell_4613 ( .C (clk), .D (signal_7158), .Q (signal_7159) ) ;
    buf_clk cell_4629 ( .C (clk), .D (signal_7174), .Q (signal_7175) ) ;
    buf_clk cell_4645 ( .C (clk), .D (signal_7190), .Q (signal_7191) ) ;
    buf_clk cell_4661 ( .C (clk), .D (signal_7206), .Q (signal_7207) ) ;
    buf_clk cell_4677 ( .C (clk), .D (signal_7222), .Q (signal_7223) ) ;
    buf_clk cell_4693 ( .C (clk), .D (signal_7238), .Q (signal_7239) ) ;
    buf_clk cell_4709 ( .C (clk), .D (signal_7254), .Q (signal_7255) ) ;
    buf_clk cell_4725 ( .C (clk), .D (signal_7270), .Q (signal_7271) ) ;
    buf_clk cell_4741 ( .C (clk), .D (signal_7286), .Q (signal_7287) ) ;
    buf_clk cell_4757 ( .C (clk), .D (signal_7302), .Q (signal_7303) ) ;
    buf_clk cell_4773 ( .C (clk), .D (signal_7318), .Q (signal_7319) ) ;
    buf_clk cell_4789 ( .C (clk), .D (signal_7334), .Q (signal_7335) ) ;
    buf_clk cell_4805 ( .C (clk), .D (signal_7350), .Q (signal_7351) ) ;
    buf_clk cell_4821 ( .C (clk), .D (signal_7366), .Q (signal_7367) ) ;
    buf_clk cell_4837 ( .C (clk), .D (signal_7382), .Q (signal_7383) ) ;
    buf_clk cell_4853 ( .C (clk), .D (signal_7398), .Q (signal_7399) ) ;
    buf_clk cell_4869 ( .C (clk), .D (signal_7414), .Q (signal_7415) ) ;
    buf_clk cell_4885 ( .C (clk), .D (signal_7430), .Q (signal_7431) ) ;
    buf_clk cell_4901 ( .C (clk), .D (signal_7446), .Q (signal_7447) ) ;
    buf_clk cell_4917 ( .C (clk), .D (signal_7462), .Q (signal_7463) ) ;
    buf_clk cell_4933 ( .C (clk), .D (signal_7478), .Q (signal_7479) ) ;
    buf_clk cell_4949 ( .C (clk), .D (signal_7494), .Q (signal_7495) ) ;
    buf_clk cell_4965 ( .C (clk), .D (signal_7510), .Q (signal_7511) ) ;
    buf_clk cell_4981 ( .C (clk), .D (signal_7526), .Q (signal_7527) ) ;
    buf_clk cell_4997 ( .C (clk), .D (signal_7542), .Q (signal_7543) ) ;
    buf_clk cell_5013 ( .C (clk), .D (signal_7558), .Q (signal_7559) ) ;
    buf_clk cell_5029 ( .C (clk), .D (signal_7574), .Q (signal_7575) ) ;
    buf_clk cell_5045 ( .C (clk), .D (signal_7590), .Q (signal_7591) ) ;
    buf_clk cell_5061 ( .C (clk), .D (signal_7606), .Q (signal_7607) ) ;
    buf_clk cell_5077 ( .C (clk), .D (signal_7622), .Q (signal_7623) ) ;
    buf_clk cell_5093 ( .C (clk), .D (signal_7638), .Q (signal_7639) ) ;
    buf_clk cell_5109 ( .C (clk), .D (signal_7654), .Q (signal_7655) ) ;
    buf_clk cell_5125 ( .C (clk), .D (signal_7670), .Q (signal_7671) ) ;
    buf_clk cell_5141 ( .C (clk), .D (signal_7686), .Q (signal_7687) ) ;
    buf_clk cell_5157 ( .C (clk), .D (signal_7702), .Q (signal_7703) ) ;
    buf_clk cell_5173 ( .C (clk), .D (signal_7718), .Q (signal_7719) ) ;
    buf_clk cell_5189 ( .C (clk), .D (signal_7734), .Q (signal_7735) ) ;
    buf_clk cell_5205 ( .C (clk), .D (signal_7750), .Q (signal_7751) ) ;
    buf_clk cell_5221 ( .C (clk), .D (signal_7766), .Q (signal_7767) ) ;
    buf_clk cell_5237 ( .C (clk), .D (signal_7782), .Q (signal_7783) ) ;
    buf_clk cell_5253 ( .C (clk), .D (signal_7798), .Q (signal_7799) ) ;
    buf_clk cell_5269 ( .C (clk), .D (signal_7814), .Q (signal_7815) ) ;
    buf_clk cell_5285 ( .C (clk), .D (signal_7830), .Q (signal_7831) ) ;
    buf_clk cell_5301 ( .C (clk), .D (signal_7846), .Q (signal_7847) ) ;
    buf_clk cell_5317 ( .C (clk), .D (signal_7862), .Q (signal_7863) ) ;
    buf_clk cell_5333 ( .C (clk), .D (signal_7878), .Q (signal_7879) ) ;
    buf_clk cell_5349 ( .C (clk), .D (signal_7894), .Q (signal_7895) ) ;
    buf_clk cell_5365 ( .C (clk), .D (signal_7910), .Q (signal_7911) ) ;
    buf_clk cell_5381 ( .C (clk), .D (signal_7926), .Q (signal_7927) ) ;
    buf_clk cell_5397 ( .C (clk), .D (signal_7942), .Q (signal_7943) ) ;
    buf_clk cell_5413 ( .C (clk), .D (signal_7958), .Q (signal_7959) ) ;
    buf_clk cell_5429 ( .C (clk), .D (signal_7974), .Q (signal_7975) ) ;
    buf_clk cell_5445 ( .C (clk), .D (signal_7990), .Q (signal_7991) ) ;
    buf_clk cell_5461 ( .C (clk), .D (signal_8006), .Q (signal_8007) ) ;
    buf_clk cell_5477 ( .C (clk), .D (signal_8022), .Q (signal_8023) ) ;
    buf_clk cell_5493 ( .C (clk), .D (signal_8038), .Q (signal_8039) ) ;
    buf_clk cell_5509 ( .C (clk), .D (signal_8054), .Q (signal_8055) ) ;
    buf_clk cell_5525 ( .C (clk), .D (signal_8070), .Q (signal_8071) ) ;
    buf_clk cell_5541 ( .C (clk), .D (signal_8086), .Q (signal_8087) ) ;
    buf_clk cell_5557 ( .C (clk), .D (signal_8102), .Q (signal_8103) ) ;
    buf_clk cell_5573 ( .C (clk), .D (signal_8118), .Q (signal_8119) ) ;
    buf_clk cell_5589 ( .C (clk), .D (signal_8134), .Q (signal_8135) ) ;
    buf_clk cell_5605 ( .C (clk), .D (signal_8150), .Q (signal_8151) ) ;
    buf_clk cell_5621 ( .C (clk), .D (signal_8166), .Q (signal_8167) ) ;
    buf_clk cell_5637 ( .C (clk), .D (signal_8182), .Q (signal_8183) ) ;
    buf_clk cell_5653 ( .C (clk), .D (signal_8198), .Q (signal_8199) ) ;
    buf_clk cell_5669 ( .C (clk), .D (signal_8214), .Q (signal_8215) ) ;
    buf_clk cell_5685 ( .C (clk), .D (signal_8230), .Q (signal_8231) ) ;
    buf_clk cell_5701 ( .C (clk), .D (signal_8246), .Q (signal_8247) ) ;
    buf_clk cell_5717 ( .C (clk), .D (signal_8262), .Q (signal_8263) ) ;
    buf_clk cell_5733 ( .C (clk), .D (signal_8278), .Q (signal_8279) ) ;
    buf_clk cell_5749 ( .C (clk), .D (signal_8294), .Q (signal_8295) ) ;
    buf_clk cell_5765 ( .C (clk), .D (signal_8310), .Q (signal_8311) ) ;
    buf_clk cell_5781 ( .C (clk), .D (signal_8326), .Q (signal_8327) ) ;
    buf_clk cell_5797 ( .C (clk), .D (signal_8342), .Q (signal_8343) ) ;
    buf_clk cell_5813 ( .C (clk), .D (signal_8358), .Q (signal_8359) ) ;
    buf_clk cell_5829 ( .C (clk), .D (signal_8374), .Q (signal_8375) ) ;
    buf_clk cell_5845 ( .C (clk), .D (signal_8390), .Q (signal_8391) ) ;
    buf_clk cell_5861 ( .C (clk), .D (signal_8406), .Q (signal_8407) ) ;
    buf_clk cell_5877 ( .C (clk), .D (signal_8422), .Q (signal_8423) ) ;
    buf_clk cell_5893 ( .C (clk), .D (signal_8438), .Q (signal_8439) ) ;
    buf_clk cell_5909 ( .C (clk), .D (signal_8454), .Q (signal_8455) ) ;
    buf_clk cell_5925 ( .C (clk), .D (signal_8470), .Q (signal_8471) ) ;
    buf_clk cell_5941 ( .C (clk), .D (signal_8486), .Q (signal_8487) ) ;
    buf_clk cell_5957 ( .C (clk), .D (signal_8502), .Q (signal_8503) ) ;
    buf_clk cell_5973 ( .C (clk), .D (signal_8518), .Q (signal_8519) ) ;
    buf_clk cell_5989 ( .C (clk), .D (signal_8534), .Q (signal_8535) ) ;
    buf_clk cell_6005 ( .C (clk), .D (signal_8550), .Q (signal_8551) ) ;
    buf_clk cell_6021 ( .C (clk), .D (signal_8566), .Q (signal_8567) ) ;
    buf_clk cell_6037 ( .C (clk), .D (signal_8582), .Q (signal_8583) ) ;
    buf_clk cell_6053 ( .C (clk), .D (signal_8598), .Q (signal_8599) ) ;
    buf_clk cell_6069 ( .C (clk), .D (signal_8614), .Q (signal_8615) ) ;
    buf_clk cell_6085 ( .C (clk), .D (signal_8630), .Q (signal_8631) ) ;
    buf_clk cell_6101 ( .C (clk), .D (signal_8646), .Q (signal_8647) ) ;
    buf_clk cell_6117 ( .C (clk), .D (signal_8662), .Q (signal_8663) ) ;
    buf_clk cell_6133 ( .C (clk), .D (signal_8678), .Q (signal_8679) ) ;
    buf_clk cell_6149 ( .C (clk), .D (signal_8694), .Q (signal_8695) ) ;
    buf_clk cell_6165 ( .C (clk), .D (signal_8710), .Q (signal_8711) ) ;
    buf_clk cell_6181 ( .C (clk), .D (signal_8726), .Q (signal_8727) ) ;
    buf_clk cell_6197 ( .C (clk), .D (signal_8742), .Q (signal_8743) ) ;
    buf_clk cell_6213 ( .C (clk), .D (signal_8758), .Q (signal_8759) ) ;
    buf_clk cell_6229 ( .C (clk), .D (signal_8774), .Q (signal_8775) ) ;
    buf_clk cell_6245 ( .C (clk), .D (signal_8790), .Q (signal_8791) ) ;
    buf_clk cell_6261 ( .C (clk), .D (signal_8806), .Q (signal_8807) ) ;
    buf_clk cell_6277 ( .C (clk), .D (signal_8822), .Q (signal_8823) ) ;
    buf_clk cell_6293 ( .C (clk), .D (signal_8838), .Q (signal_8839) ) ;
    buf_clk cell_6309 ( .C (clk), .D (signal_8854), .Q (signal_8855) ) ;
    buf_clk cell_6325 ( .C (clk), .D (signal_8870), .Q (signal_8871) ) ;
    buf_clk cell_6341 ( .C (clk), .D (signal_8886), .Q (signal_8887) ) ;
    buf_clk cell_6357 ( .C (clk), .D (signal_8902), .Q (signal_8903) ) ;
    buf_clk cell_6373 ( .C (clk), .D (signal_8918), .Q (signal_8919) ) ;
    buf_clk cell_6389 ( .C (clk), .D (signal_8934), .Q (signal_8935) ) ;
    buf_clk cell_6405 ( .C (clk), .D (signal_8950), .Q (signal_8951) ) ;
    buf_clk cell_6421 ( .C (clk), .D (signal_8966), .Q (signal_8967) ) ;
    buf_clk cell_6437 ( .C (clk), .D (signal_8982), .Q (signal_8983) ) ;
    buf_clk cell_6453 ( .C (clk), .D (signal_8998), .Q (signal_8999) ) ;
    buf_clk cell_6469 ( .C (clk), .D (signal_9014), .Q (signal_9015) ) ;
    buf_clk cell_6485 ( .C (clk), .D (signal_9030), .Q (signal_9031) ) ;
    buf_clk cell_6501 ( .C (clk), .D (signal_9046), .Q (signal_9047) ) ;
    buf_clk cell_6517 ( .C (clk), .D (signal_9062), .Q (signal_9063) ) ;
    buf_clk cell_6533 ( .C (clk), .D (signal_9078), .Q (signal_9079) ) ;
    buf_clk cell_6549 ( .C (clk), .D (signal_9094), .Q (signal_9095) ) ;
    buf_clk cell_6565 ( .C (clk), .D (signal_9110), .Q (signal_9111) ) ;
    buf_clk cell_6581 ( .C (clk), .D (signal_9126), .Q (signal_9127) ) ;
    buf_clk cell_6597 ( .C (clk), .D (signal_9142), .Q (signal_9143) ) ;
    buf_clk cell_6613 ( .C (clk), .D (signal_9158), .Q (signal_9159) ) ;
    buf_clk cell_6629 ( .C (clk), .D (signal_9174), .Q (signal_9175) ) ;
    buf_clk cell_6645 ( .C (clk), .D (signal_9190), .Q (signal_9191) ) ;
    buf_clk cell_6661 ( .C (clk), .D (signal_9206), .Q (signal_9207) ) ;
    buf_clk cell_6677 ( .C (clk), .D (signal_9222), .Q (signal_9223) ) ;
    buf_clk cell_6693 ( .C (clk), .D (signal_9238), .Q (signal_9239) ) ;
    buf_clk cell_6709 ( .C (clk), .D (signal_9254), .Q (signal_9255) ) ;
    buf_clk cell_6725 ( .C (clk), .D (signal_9270), .Q (signal_9271) ) ;
    buf_clk cell_6741 ( .C (clk), .D (signal_9286), .Q (signal_9287) ) ;
    buf_clk cell_6757 ( .C (clk), .D (signal_9302), .Q (signal_9303) ) ;
    buf_clk cell_6773 ( .C (clk), .D (signal_9318), .Q (signal_9319) ) ;
    buf_clk cell_6789 ( .C (clk), .D (signal_9334), .Q (signal_9335) ) ;
    buf_clk cell_6805 ( .C (clk), .D (signal_9350), .Q (signal_9351) ) ;
    buf_clk cell_6821 ( .C (clk), .D (signal_9366), .Q (signal_9367) ) ;
    buf_clk cell_6837 ( .C (clk), .D (signal_9382), .Q (signal_9383) ) ;
    buf_clk cell_6853 ( .C (clk), .D (signal_9398), .Q (signal_9399) ) ;
    buf_clk cell_6869 ( .C (clk), .D (signal_9414), .Q (signal_9415) ) ;
    buf_clk cell_6885 ( .C (clk), .D (signal_9430), .Q (signal_9431) ) ;
    buf_clk cell_6901 ( .C (clk), .D (signal_9446), .Q (signal_9447) ) ;
    buf_clk cell_6917 ( .C (clk), .D (signal_9462), .Q (signal_9463) ) ;
    buf_clk cell_6933 ( .C (clk), .D (signal_9478), .Q (signal_9479) ) ;
    buf_clk cell_6949 ( .C (clk), .D (signal_9494), .Q (signal_9495) ) ;
    buf_clk cell_6965 ( .C (clk), .D (signal_9510), .Q (signal_9511) ) ;
    buf_clk cell_6981 ( .C (clk), .D (signal_9526), .Q (signal_9527) ) ;
    buf_clk cell_6997 ( .C (clk), .D (signal_9542), .Q (signal_9543) ) ;
    buf_clk cell_7013 ( .C (clk), .D (signal_9558), .Q (signal_9559) ) ;
    buf_clk cell_7029 ( .C (clk), .D (signal_9574), .Q (signal_9575) ) ;
    buf_clk cell_7045 ( .C (clk), .D (signal_9590), .Q (signal_9591) ) ;
    buf_clk cell_7061 ( .C (clk), .D (signal_9606), .Q (signal_9607) ) ;
    buf_clk cell_7077 ( .C (clk), .D (signal_9622), .Q (signal_9623) ) ;
    buf_clk cell_7093 ( .C (clk), .D (signal_9638), .Q (signal_9639) ) ;
    buf_clk cell_7109 ( .C (clk), .D (signal_9654), .Q (signal_9655) ) ;
    buf_clk cell_7125 ( .C (clk), .D (signal_9670), .Q (signal_9671) ) ;
    buf_clk cell_7141 ( .C (clk), .D (signal_9686), .Q (signal_9687) ) ;
    buf_clk cell_7157 ( .C (clk), .D (signal_9702), .Q (signal_9703) ) ;
    buf_clk cell_7173 ( .C (clk), .D (signal_9718), .Q (signal_9719) ) ;
    buf_clk cell_7189 ( .C (clk), .D (signal_9734), .Q (signal_9735) ) ;
    buf_clk cell_7205 ( .C (clk), .D (signal_9750), .Q (signal_9751) ) ;
    buf_clk cell_7221 ( .C (clk), .D (signal_9766), .Q (signal_9767) ) ;
    buf_clk cell_7237 ( .C (clk), .D (signal_9782), .Q (signal_9783) ) ;
    buf_clk cell_7253 ( .C (clk), .D (signal_9798), .Q (signal_9799) ) ;
    buf_clk cell_7269 ( .C (clk), .D (signal_9814), .Q (signal_9815) ) ;
    buf_clk cell_7285 ( .C (clk), .D (signal_9830), .Q (signal_9831) ) ;
    buf_clk cell_7301 ( .C (clk), .D (signal_9846), .Q (signal_9847) ) ;
    buf_clk cell_7317 ( .C (clk), .D (signal_9862), .Q (signal_9863) ) ;
    buf_clk cell_7333 ( .C (clk), .D (signal_9878), .Q (signal_9879) ) ;
    buf_clk cell_7349 ( .C (clk), .D (signal_9894), .Q (signal_9895) ) ;
    buf_clk cell_7365 ( .C (clk), .D (signal_9910), .Q (signal_9911) ) ;
    buf_clk cell_7381 ( .C (clk), .D (signal_9926), .Q (signal_9927) ) ;
    buf_clk cell_7397 ( .C (clk), .D (signal_9942), .Q (signal_9943) ) ;
    buf_clk cell_7413 ( .C (clk), .D (signal_9958), .Q (signal_9959) ) ;
    buf_clk cell_7429 ( .C (clk), .D (signal_9974), .Q (signal_9975) ) ;
    buf_clk cell_7445 ( .C (clk), .D (signal_9990), .Q (signal_9991) ) ;
    buf_clk cell_7461 ( .C (clk), .D (signal_10006), .Q (signal_10007) ) ;
    buf_clk cell_7477 ( .C (clk), .D (signal_10022), .Q (signal_10023) ) ;
    buf_clk cell_7493 ( .C (clk), .D (signal_10038), .Q (signal_10039) ) ;
    buf_clk cell_7509 ( .C (clk), .D (signal_10054), .Q (signal_10055) ) ;
    buf_clk cell_7525 ( .C (clk), .D (signal_10070), .Q (signal_10071) ) ;
    buf_clk cell_7541 ( .C (clk), .D (signal_10086), .Q (signal_10087) ) ;
    buf_clk cell_7557 ( .C (clk), .D (signal_10102), .Q (signal_10103) ) ;
    buf_clk cell_7573 ( .C (clk), .D (signal_10118), .Q (signal_10119) ) ;
    buf_clk cell_7589 ( .C (clk), .D (signal_10134), .Q (signal_10135) ) ;
    buf_clk cell_7605 ( .C (clk), .D (signal_10150), .Q (signal_10151) ) ;
    buf_clk cell_7621 ( .C (clk), .D (signal_10166), .Q (signal_10167) ) ;
    buf_clk cell_7637 ( .C (clk), .D (signal_10182), .Q (signal_10183) ) ;
    buf_clk cell_7653 ( .C (clk), .D (signal_10198), .Q (signal_10199) ) ;
    buf_clk cell_7669 ( .C (clk), .D (signal_10214), .Q (signal_10215) ) ;
    buf_clk cell_7685 ( .C (clk), .D (signal_10230), .Q (signal_10231) ) ;
    buf_clk cell_7701 ( .C (clk), .D (signal_10246), .Q (signal_10247) ) ;
    buf_clk cell_7717 ( .C (clk), .D (signal_10262), .Q (signal_10263) ) ;
    buf_clk cell_7733 ( .C (clk), .D (signal_10278), .Q (signal_10279) ) ;
    buf_clk cell_7749 ( .C (clk), .D (signal_10294), .Q (signal_10295) ) ;
    buf_clk cell_7765 ( .C (clk), .D (signal_10310), .Q (signal_10311) ) ;
    buf_clk cell_7781 ( .C (clk), .D (signal_10326), .Q (signal_10327) ) ;
    buf_clk cell_7797 ( .C (clk), .D (signal_10342), .Q (signal_10343) ) ;
    buf_clk cell_7813 ( .C (clk), .D (signal_10358), .Q (signal_10359) ) ;
    buf_clk cell_7829 ( .C (clk), .D (signal_10374), .Q (signal_10375) ) ;
    buf_clk cell_7845 ( .C (clk), .D (signal_10390), .Q (signal_10391) ) ;
    buf_clk cell_7861 ( .C (clk), .D (signal_10406), .Q (signal_10407) ) ;
    buf_clk cell_7877 ( .C (clk), .D (signal_10422), .Q (signal_10423) ) ;
    buf_clk cell_7893 ( .C (clk), .D (signal_10438), .Q (signal_10439) ) ;
    buf_clk cell_7909 ( .C (clk), .D (signal_10454), .Q (signal_10455) ) ;
    buf_clk cell_7925 ( .C (clk), .D (signal_10470), .Q (signal_10471) ) ;
    buf_clk cell_7941 ( .C (clk), .D (signal_10486), .Q (signal_10487) ) ;
    buf_clk cell_7957 ( .C (clk), .D (signal_10502), .Q (signal_10503) ) ;
    buf_clk cell_7973 ( .C (clk), .D (signal_10518), .Q (signal_10519) ) ;
    buf_clk cell_7989 ( .C (clk), .D (signal_10534), .Q (signal_10535) ) ;
    buf_clk cell_8005 ( .C (clk), .D (signal_10550), .Q (signal_10551) ) ;
    buf_clk cell_8021 ( .C (clk), .D (signal_10566), .Q (signal_10567) ) ;
    buf_clk cell_8037 ( .C (clk), .D (signal_10582), .Q (signal_10583) ) ;
    buf_clk cell_8053 ( .C (clk), .D (signal_10598), .Q (signal_10599) ) ;
    buf_clk cell_8069 ( .C (clk), .D (signal_10614), .Q (signal_10615) ) ;
    buf_clk cell_8085 ( .C (clk), .D (signal_10630), .Q (signal_10631) ) ;
    buf_clk cell_8101 ( .C (clk), .D (signal_10646), .Q (signal_10647) ) ;
    buf_clk cell_8117 ( .C (clk), .D (signal_10662), .Q (signal_10663) ) ;
    buf_clk cell_8133 ( .C (clk), .D (signal_10678), .Q (signal_10679) ) ;
    buf_clk cell_8149 ( .C (clk), .D (signal_10694), .Q (signal_10695) ) ;
    buf_clk cell_8165 ( .C (clk), .D (signal_10710), .Q (signal_10711) ) ;
    buf_clk cell_8181 ( .C (clk), .D (signal_10726), .Q (signal_10727) ) ;
    buf_clk cell_8197 ( .C (clk), .D (signal_10742), .Q (signal_10743) ) ;
    buf_clk cell_8213 ( .C (clk), .D (signal_10758), .Q (signal_10759) ) ;
    buf_clk cell_8229 ( .C (clk), .D (signal_10774), .Q (signal_10775) ) ;
    buf_clk cell_8245 ( .C (clk), .D (signal_10790), .Q (signal_10791) ) ;
    buf_clk cell_8261 ( .C (clk), .D (signal_10806), .Q (signal_10807) ) ;
    buf_clk cell_8277 ( .C (clk), .D (signal_10822), .Q (signal_10823) ) ;
    buf_clk cell_8293 ( .C (clk), .D (signal_10838), .Q (signal_10839) ) ;
    buf_clk cell_8309 ( .C (clk), .D (signal_10854), .Q (signal_10855) ) ;
    buf_clk cell_8325 ( .C (clk), .D (signal_10870), .Q (signal_10871) ) ;
    buf_clk cell_8341 ( .C (clk), .D (signal_10886), .Q (signal_10887) ) ;
    buf_clk cell_8357 ( .C (clk), .D (signal_10902), .Q (signal_10903) ) ;
    buf_clk cell_8373 ( .C (clk), .D (signal_10918), .Q (signal_10919) ) ;
    buf_clk cell_8389 ( .C (clk), .D (signal_10934), .Q (signal_10935) ) ;
    buf_clk cell_8405 ( .C (clk), .D (signal_10950), .Q (signal_10951) ) ;
    buf_clk cell_8421 ( .C (clk), .D (signal_10966), .Q (signal_10967) ) ;
    buf_clk cell_8437 ( .C (clk), .D (signal_10982), .Q (signal_10983) ) ;
    buf_clk cell_8453 ( .C (clk), .D (signal_10998), .Q (signal_10999) ) ;
    buf_clk cell_8469 ( .C (clk), .D (signal_11014), .Q (signal_11015) ) ;
    buf_clk cell_8485 ( .C (clk), .D (signal_11030), .Q (signal_11031) ) ;
    buf_clk cell_8501 ( .C (clk), .D (signal_11046), .Q (signal_11047) ) ;
    buf_clk cell_8517 ( .C (clk), .D (signal_11062), .Q (signal_11063) ) ;
    buf_clk cell_8533 ( .C (clk), .D (signal_11078), .Q (signal_11079) ) ;
    buf_clk cell_8549 ( .C (clk), .D (signal_11094), .Q (signal_11095) ) ;
    buf_clk cell_8565 ( .C (clk), .D (signal_11110), .Q (signal_11111) ) ;
    buf_clk cell_8581 ( .C (clk), .D (signal_11126), .Q (signal_11127) ) ;
    buf_clk cell_8597 ( .C (clk), .D (signal_11142), .Q (signal_11143) ) ;
    buf_clk cell_8613 ( .C (clk), .D (signal_11158), .Q (signal_11159) ) ;
    buf_clk cell_8629 ( .C (clk), .D (signal_11174), .Q (signal_11175) ) ;
    buf_clk cell_8645 ( .C (clk), .D (signal_11190), .Q (signal_11191) ) ;
    buf_clk cell_8661 ( .C (clk), .D (signal_11206), .Q (signal_11207) ) ;
    buf_clk cell_8677 ( .C (clk), .D (signal_11222), .Q (signal_11223) ) ;
    buf_clk cell_8693 ( .C (clk), .D (signal_11238), .Q (signal_11239) ) ;
    buf_clk cell_8709 ( .C (clk), .D (signal_11254), .Q (signal_11255) ) ;
    buf_clk cell_8725 ( .C (clk), .D (signal_11270), .Q (signal_11271) ) ;
    buf_clk cell_8741 ( .C (clk), .D (signal_11286), .Q (signal_11287) ) ;
    buf_clk cell_8757 ( .C (clk), .D (signal_11302), .Q (signal_11303) ) ;
    buf_clk cell_8773 ( .C (clk), .D (signal_11318), .Q (signal_11319) ) ;
    buf_clk cell_8789 ( .C (clk), .D (signal_11334), .Q (signal_11335) ) ;
    buf_clk cell_8805 ( .C (clk), .D (signal_11350), .Q (signal_11351) ) ;
    buf_clk cell_8821 ( .C (clk), .D (signal_11366), .Q (signal_11367) ) ;
    buf_clk cell_8837 ( .C (clk), .D (signal_11382), .Q (signal_11383) ) ;
    buf_clk cell_8853 ( .C (clk), .D (signal_11398), .Q (signal_11399) ) ;
    buf_clk cell_8869 ( .C (clk), .D (signal_11414), .Q (signal_11415) ) ;
    buf_clk cell_8885 ( .C (clk), .D (signal_11430), .Q (signal_11431) ) ;
    buf_clk cell_8901 ( .C (clk), .D (signal_11446), .Q (signal_11447) ) ;
    buf_clk cell_8917 ( .C (clk), .D (signal_11462), .Q (signal_11463) ) ;
    buf_clk cell_8933 ( .C (clk), .D (signal_11478), .Q (signal_11479) ) ;
    buf_clk cell_8949 ( .C (clk), .D (signal_11494), .Q (signal_11495) ) ;
    buf_clk cell_8965 ( .C (clk), .D (signal_11510), .Q (signal_11511) ) ;
    buf_clk cell_8981 ( .C (clk), .D (signal_11526), .Q (signal_11527) ) ;
    buf_clk cell_8997 ( .C (clk), .D (signal_11542), .Q (signal_11543) ) ;
    buf_clk cell_9013 ( .C (clk), .D (signal_11558), .Q (signal_11559) ) ;
    buf_clk cell_9029 ( .C (clk), .D (signal_11574), .Q (signal_11575) ) ;
    buf_clk cell_9045 ( .C (clk), .D (signal_11590), .Q (signal_11591) ) ;
    buf_clk cell_9061 ( .C (clk), .D (signal_11606), .Q (signal_11607) ) ;
    buf_clk cell_9077 ( .C (clk), .D (signal_11622), .Q (signal_11623) ) ;
    buf_clk cell_9093 ( .C (clk), .D (signal_11638), .Q (signal_11639) ) ;
    buf_clk cell_9109 ( .C (clk), .D (signal_11654), .Q (signal_11655) ) ;
    buf_clk cell_9125 ( .C (clk), .D (signal_11670), .Q (signal_11671) ) ;
    buf_clk cell_9141 ( .C (clk), .D (signal_11686), .Q (signal_11687) ) ;
    buf_clk cell_9157 ( .C (clk), .D (signal_11702), .Q (signal_11703) ) ;
    buf_clk cell_9173 ( .C (clk), .D (signal_11718), .Q (signal_11719) ) ;
    buf_clk cell_9189 ( .C (clk), .D (signal_11734), .Q (signal_11735) ) ;
    buf_clk cell_9205 ( .C (clk), .D (signal_11750), .Q (signal_11751) ) ;
    buf_clk cell_9221 ( .C (clk), .D (signal_11766), .Q (signal_11767) ) ;
    buf_clk cell_9237 ( .C (clk), .D (signal_11782), .Q (signal_11783) ) ;
    buf_clk cell_9253 ( .C (clk), .D (signal_11798), .Q (signal_11799) ) ;
    buf_clk cell_9269 ( .C (clk), .D (signal_11814), .Q (signal_11815) ) ;
    buf_clk cell_9285 ( .C (clk), .D (signal_11830), .Q (signal_11831) ) ;
    buf_clk cell_9301 ( .C (clk), .D (signal_11846), .Q (signal_11847) ) ;
    buf_clk cell_9317 ( .C (clk), .D (signal_11862), .Q (signal_11863) ) ;
    buf_clk cell_9333 ( .C (clk), .D (signal_11878), .Q (signal_11879) ) ;
    buf_clk cell_9349 ( .C (clk), .D (signal_11894), .Q (signal_11895) ) ;
    buf_clk cell_9365 ( .C (clk), .D (signal_11910), .Q (signal_11911) ) ;
    buf_clk cell_9381 ( .C (clk), .D (signal_11926), .Q (signal_11927) ) ;
    buf_clk cell_9397 ( .C (clk), .D (signal_11942), .Q (signal_11943) ) ;
    buf_clk cell_9413 ( .C (clk), .D (signal_11958), .Q (signal_11959) ) ;
    buf_clk cell_9429 ( .C (clk), .D (signal_11974), .Q (signal_11975) ) ;
    buf_clk cell_9445 ( .C (clk), .D (signal_11990), .Q (signal_11991) ) ;
    buf_clk cell_9461 ( .C (clk), .D (signal_12006), .Q (signal_12007) ) ;
    buf_clk cell_9477 ( .C (clk), .D (signal_12022), .Q (signal_12023) ) ;
    buf_clk cell_9493 ( .C (clk), .D (signal_12038), .Q (signal_12039) ) ;
    buf_clk cell_9509 ( .C (clk), .D (signal_12054), .Q (signal_12055) ) ;
    buf_clk cell_9525 ( .C (clk), .D (signal_12070), .Q (signal_12071) ) ;
    buf_clk cell_9541 ( .C (clk), .D (signal_12086), .Q (signal_12087) ) ;
    buf_clk cell_9557 ( .C (clk), .D (signal_12102), .Q (signal_12103) ) ;
    buf_clk cell_9573 ( .C (clk), .D (signal_12118), .Q (signal_12119) ) ;
    buf_clk cell_9589 ( .C (clk), .D (signal_12134), .Q (signal_12135) ) ;
    buf_clk cell_9605 ( .C (clk), .D (signal_12150), .Q (signal_12151) ) ;
    buf_clk cell_9621 ( .C (clk), .D (signal_12166), .Q (signal_12167) ) ;
    buf_clk cell_9637 ( .C (clk), .D (signal_12182), .Q (signal_12183) ) ;
    buf_clk cell_9653 ( .C (clk), .D (signal_12198), .Q (signal_12199) ) ;
    buf_clk cell_9669 ( .C (clk), .D (signal_12214), .Q (signal_12215) ) ;
    buf_clk cell_9685 ( .C (clk), .D (signal_12230), .Q (signal_12231) ) ;
    buf_clk cell_9701 ( .C (clk), .D (signal_12246), .Q (signal_12247) ) ;
    buf_clk cell_9717 ( .C (clk), .D (signal_12262), .Q (signal_12263) ) ;
    buf_clk cell_9733 ( .C (clk), .D (signal_12278), .Q (signal_12279) ) ;
    buf_clk cell_9749 ( .C (clk), .D (signal_12294), .Q (signal_12295) ) ;
    buf_clk cell_9765 ( .C (clk), .D (signal_12310), .Q (signal_12311) ) ;
    buf_clk cell_9781 ( .C (clk), .D (signal_12326), .Q (signal_12327) ) ;
    buf_clk cell_9797 ( .C (clk), .D (signal_12342), .Q (signal_12343) ) ;
    buf_clk cell_9813 ( .C (clk), .D (signal_12358), .Q (signal_12359) ) ;
    buf_clk cell_9829 ( .C (clk), .D (signal_12374), .Q (signal_12375) ) ;
    buf_clk cell_9845 ( .C (clk), .D (signal_12390), .Q (signal_12391) ) ;
    buf_clk cell_9861 ( .C (clk), .D (signal_12406), .Q (signal_12407) ) ;
    buf_clk cell_9877 ( .C (clk), .D (signal_12422), .Q (signal_12423) ) ;
    buf_clk cell_9893 ( .C (clk), .D (signal_12438), .Q (signal_12439) ) ;
    buf_clk cell_9909 ( .C (clk), .D (signal_12454), .Q (signal_12455) ) ;
    buf_clk cell_9925 ( .C (clk), .D (signal_12470), .Q (signal_12471) ) ;
    buf_clk cell_9941 ( .C (clk), .D (signal_12486), .Q (signal_12487) ) ;
    buf_clk cell_9957 ( .C (clk), .D (signal_12502), .Q (signal_12503) ) ;
    buf_clk cell_9973 ( .C (clk), .D (signal_12518), .Q (signal_12519) ) ;
    buf_clk cell_9989 ( .C (clk), .D (signal_12534), .Q (signal_12535) ) ;
    buf_clk cell_10005 ( .C (clk), .D (signal_12550), .Q (signal_12551) ) ;
    buf_clk cell_10021 ( .C (clk), .D (signal_12566), .Q (signal_12567) ) ;
    buf_clk cell_10037 ( .C (clk), .D (signal_12582), .Q (signal_12583) ) ;
    buf_clk cell_10053 ( .C (clk), .D (signal_12598), .Q (signal_12599) ) ;
    buf_clk cell_10069 ( .C (clk), .D (signal_12614), .Q (signal_12615) ) ;
    buf_clk cell_10085 ( .C (clk), .D (signal_12630), .Q (signal_12631) ) ;
    buf_clk cell_10101 ( .C (clk), .D (signal_12646), .Q (signal_12647) ) ;
    buf_clk cell_10117 ( .C (clk), .D (signal_12662), .Q (signal_12663) ) ;
    buf_clk cell_10133 ( .C (clk), .D (signal_12678), .Q (signal_12679) ) ;
    buf_clk cell_10149 ( .C (clk), .D (signal_12694), .Q (signal_12695) ) ;
    buf_clk cell_10165 ( .C (clk), .D (signal_12710), .Q (signal_12711) ) ;
    buf_clk cell_10181 ( .C (clk), .D (signal_12726), .Q (signal_12727) ) ;
    buf_clk cell_10197 ( .C (clk), .D (signal_12742), .Q (signal_12743) ) ;
    buf_clk cell_10213 ( .C (clk), .D (signal_12758), .Q (signal_12759) ) ;
    buf_clk cell_10229 ( .C (clk), .D (signal_12774), .Q (signal_12775) ) ;
    buf_clk cell_10245 ( .C (clk), .D (signal_12790), .Q (signal_12791) ) ;
    buf_clk cell_10261 ( .C (clk), .D (signal_12806), .Q (signal_12807) ) ;
    buf_clk cell_10277 ( .C (clk), .D (signal_12822), .Q (signal_12823) ) ;
    buf_clk cell_10293 ( .C (clk), .D (signal_12838), .Q (signal_12839) ) ;
    buf_clk cell_10309 ( .C (clk), .D (signal_12854), .Q (signal_12855) ) ;
    buf_clk cell_10325 ( .C (clk), .D (signal_12870), .Q (signal_12871) ) ;
    buf_clk cell_10341 ( .C (clk), .D (signal_12886), .Q (signal_12887) ) ;
    buf_clk cell_10357 ( .C (clk), .D (signal_12902), .Q (signal_12903) ) ;
    buf_clk cell_10373 ( .C (clk), .D (signal_12918), .Q (signal_12919) ) ;
    buf_clk cell_10389 ( .C (clk), .D (signal_12934), .Q (signal_12935) ) ;
    buf_clk cell_10405 ( .C (clk), .D (signal_12950), .Q (signal_12951) ) ;
    buf_clk cell_10421 ( .C (clk), .D (signal_12966), .Q (signal_12967) ) ;
    buf_clk cell_10437 ( .C (clk), .D (signal_12982), .Q (signal_12983) ) ;
    buf_clk cell_10453 ( .C (clk), .D (signal_12998), .Q (signal_12999) ) ;
    buf_clk cell_10469 ( .C (clk), .D (signal_13014), .Q (signal_13015) ) ;
    buf_clk cell_10485 ( .C (clk), .D (signal_13030), .Q (signal_13031) ) ;
    buf_clk cell_10501 ( .C (clk), .D (signal_13046), .Q (signal_13047) ) ;
    buf_clk cell_10517 ( .C (clk), .D (signal_13062), .Q (signal_13063) ) ;
    buf_clk cell_10533 ( .C (clk), .D (signal_13078), .Q (signal_13079) ) ;
    buf_clk cell_10549 ( .C (clk), .D (signal_13094), .Q (signal_13095) ) ;
    buf_clk cell_10565 ( .C (clk), .D (signal_13110), .Q (signal_13111) ) ;
    buf_clk cell_10581 ( .C (clk), .D (signal_13126), .Q (signal_13127) ) ;
    buf_clk cell_10597 ( .C (clk), .D (signal_13142), .Q (signal_13143) ) ;
    buf_clk cell_10613 ( .C (clk), .D (signal_13158), .Q (signal_13159) ) ;
    buf_clk cell_10629 ( .C (clk), .D (signal_13174), .Q (signal_13175) ) ;
    buf_clk cell_10645 ( .C (clk), .D (signal_13190), .Q (signal_13191) ) ;
    buf_clk cell_10661 ( .C (clk), .D (signal_13206), .Q (signal_13207) ) ;
    buf_clk cell_10677 ( .C (clk), .D (signal_13222), .Q (signal_13223) ) ;
    buf_clk cell_10693 ( .C (clk), .D (signal_13238), .Q (signal_13239) ) ;
    buf_clk cell_10709 ( .C (clk), .D (signal_13254), .Q (signal_13255) ) ;
    buf_clk cell_10725 ( .C (clk), .D (signal_13270), .Q (signal_13271) ) ;
    buf_clk cell_10741 ( .C (clk), .D (signal_13286), .Q (signal_13287) ) ;
    buf_clk cell_10757 ( .C (clk), .D (signal_13302), .Q (signal_13303) ) ;
    buf_clk cell_10773 ( .C (clk), .D (signal_13318), .Q (signal_13319) ) ;
    buf_clk cell_10789 ( .C (clk), .D (signal_13334), .Q (signal_13335) ) ;
    buf_clk cell_10805 ( .C (clk), .D (signal_13350), .Q (signal_13351) ) ;
    buf_clk cell_10821 ( .C (clk), .D (signal_13366), .Q (signal_13367) ) ;
    buf_clk cell_10837 ( .C (clk), .D (signal_13382), .Q (signal_13383) ) ;
    buf_clk cell_10853 ( .C (clk), .D (signal_13398), .Q (signal_13399) ) ;
    buf_clk cell_10869 ( .C (clk), .D (signal_13414), .Q (signal_13415) ) ;
    buf_clk cell_10885 ( .C (clk), .D (signal_13430), .Q (signal_13431) ) ;
    buf_clk cell_10901 ( .C (clk), .D (signal_13446), .Q (signal_13447) ) ;
    buf_clk cell_10917 ( .C (clk), .D (signal_13462), .Q (signal_13463) ) ;
    buf_clk cell_10933 ( .C (clk), .D (signal_13478), .Q (signal_13479) ) ;
    buf_clk cell_10949 ( .C (clk), .D (signal_13494), .Q (signal_13495) ) ;
    buf_clk cell_10965 ( .C (clk), .D (signal_13510), .Q (signal_13511) ) ;
    buf_clk cell_10981 ( .C (clk), .D (signal_13526), .Q (signal_13527) ) ;
    buf_clk cell_10997 ( .C (clk), .D (signal_13542), .Q (signal_13543) ) ;
    buf_clk cell_11013 ( .C (clk), .D (signal_13558), .Q (signal_13559) ) ;
    buf_clk cell_11029 ( .C (clk), .D (signal_13574), .Q (signal_13575) ) ;
    buf_clk cell_11045 ( .C (clk), .D (signal_13590), .Q (signal_13591) ) ;
    buf_clk cell_11061 ( .C (clk), .D (signal_13606), .Q (signal_13607) ) ;
    buf_clk cell_11077 ( .C (clk), .D (signal_13622), .Q (signal_13623) ) ;
    buf_clk cell_11093 ( .C (clk), .D (signal_13638), .Q (signal_13639) ) ;
    buf_clk cell_11109 ( .C (clk), .D (signal_13654), .Q (signal_13655) ) ;
    buf_clk cell_11125 ( .C (clk), .D (signal_13670), .Q (signal_13671) ) ;
    buf_clk cell_11141 ( .C (clk), .D (signal_13686), .Q (signal_13687) ) ;
    buf_clk cell_11157 ( .C (clk), .D (signal_13702), .Q (signal_13703) ) ;
    buf_clk cell_11173 ( .C (clk), .D (signal_13718), .Q (signal_13719) ) ;
    buf_clk cell_11189 ( .C (clk), .D (signal_13734), .Q (signal_13735) ) ;
    buf_clk cell_11205 ( .C (clk), .D (signal_13750), .Q (signal_13751) ) ;
    buf_clk cell_11221 ( .C (clk), .D (signal_13766), .Q (signal_13767) ) ;
    buf_clk cell_11237 ( .C (clk), .D (signal_13782), .Q (signal_13783) ) ;
    buf_clk cell_11253 ( .C (clk), .D (signal_13798), .Q (signal_13799) ) ;
    buf_clk cell_11269 ( .C (clk), .D (signal_13814), .Q (signal_13815) ) ;
    buf_clk cell_11285 ( .C (clk), .D (signal_13830), .Q (signal_13831) ) ;
    buf_clk cell_11301 ( .C (clk), .D (signal_13846), .Q (signal_13847) ) ;
    buf_clk cell_11317 ( .C (clk), .D (signal_13862), .Q (signal_13863) ) ;
    buf_clk cell_11333 ( .C (clk), .D (signal_13878), .Q (signal_13879) ) ;
    buf_clk cell_11349 ( .C (clk), .D (signal_13894), .Q (signal_13895) ) ;
    buf_clk cell_11365 ( .C (clk), .D (signal_13910), .Q (signal_13911) ) ;
    buf_clk cell_11381 ( .C (clk), .D (signal_13926), .Q (signal_13927) ) ;
    buf_clk cell_11397 ( .C (clk), .D (signal_13942), .Q (signal_13943) ) ;
    buf_clk cell_11413 ( .C (clk), .D (signal_13958), .Q (signal_13959) ) ;
    buf_clk cell_11429 ( .C (clk), .D (signal_13974), .Q (signal_13975) ) ;
    buf_clk cell_11445 ( .C (clk), .D (signal_13990), .Q (signal_13991) ) ;
    buf_clk cell_11461 ( .C (clk), .D (signal_14006), .Q (signal_14007) ) ;
    buf_clk cell_11477 ( .C (clk), .D (signal_14022), .Q (signal_14023) ) ;
    buf_clk cell_11493 ( .C (clk), .D (signal_14038), .Q (signal_14039) ) ;
    buf_clk cell_11509 ( .C (clk), .D (signal_14054), .Q (signal_14055) ) ;
    buf_clk cell_11525 ( .C (clk), .D (signal_14070), .Q (signal_14071) ) ;
    buf_clk cell_11541 ( .C (clk), .D (signal_14086), .Q (signal_14087) ) ;
    buf_clk cell_11557 ( .C (clk), .D (signal_14102), .Q (signal_14103) ) ;
    buf_clk cell_11573 ( .C (clk), .D (signal_14118), .Q (signal_14119) ) ;
    buf_clk cell_11589 ( .C (clk), .D (signal_14134), .Q (signal_14135) ) ;
    buf_clk cell_11605 ( .C (clk), .D (signal_14150), .Q (signal_14151) ) ;
    buf_clk cell_11621 ( .C (clk), .D (signal_14166), .Q (signal_14167) ) ;
    buf_clk cell_11637 ( .C (clk), .D (signal_14182), .Q (signal_14183) ) ;
    buf_clk cell_11653 ( .C (clk), .D (signal_14198), .Q (signal_14199) ) ;
    buf_clk cell_11669 ( .C (clk), .D (signal_14214), .Q (signal_14215) ) ;
    buf_clk cell_11685 ( .C (clk), .D (signal_14230), .Q (signal_14231) ) ;
    buf_clk cell_11701 ( .C (clk), .D (signal_14246), .Q (signal_14247) ) ;
    buf_clk cell_11717 ( .C (clk), .D (signal_14262), .Q (signal_14263) ) ;
    buf_clk cell_11733 ( .C (clk), .D (signal_14278), .Q (signal_14279) ) ;
    buf_clk cell_11749 ( .C (clk), .D (signal_14294), .Q (signal_14295) ) ;
    buf_clk cell_11765 ( .C (clk), .D (signal_14310), .Q (signal_14311) ) ;
    buf_clk cell_11781 ( .C (clk), .D (signal_14326), .Q (signal_14327) ) ;
    buf_clk cell_11797 ( .C (clk), .D (signal_14342), .Q (signal_14343) ) ;
    buf_clk cell_11813 ( .C (clk), .D (signal_14358), .Q (signal_14359) ) ;
    buf_clk cell_11829 ( .C (clk), .D (signal_14374), .Q (signal_14375) ) ;
    buf_clk cell_11845 ( .C (clk), .D (signal_14390), .Q (signal_14391) ) ;
    buf_clk cell_11861 ( .C (clk), .D (signal_14406), .Q (signal_14407) ) ;
    buf_clk cell_11877 ( .C (clk), .D (signal_14422), .Q (signal_14423) ) ;
    buf_clk cell_11893 ( .C (clk), .D (signal_14438), .Q (signal_14439) ) ;
    buf_clk cell_11909 ( .C (clk), .D (signal_14454), .Q (signal_14455) ) ;
    buf_clk cell_11925 ( .C (clk), .D (signal_14470), .Q (signal_14471) ) ;
    buf_clk cell_11941 ( .C (clk), .D (signal_14486), .Q (signal_14487) ) ;
    buf_clk cell_11957 ( .C (clk), .D (signal_14502), .Q (signal_14503) ) ;
    buf_clk cell_11973 ( .C (clk), .D (signal_14518), .Q (signal_14519) ) ;
    buf_clk cell_11989 ( .C (clk), .D (signal_14534), .Q (signal_14535) ) ;
    buf_clk cell_12005 ( .C (clk), .D (signal_14550), .Q (signal_14551) ) ;
    buf_clk cell_12021 ( .C (clk), .D (signal_14566), .Q (signal_14567) ) ;
    buf_clk cell_12037 ( .C (clk), .D (signal_14582), .Q (signal_14583) ) ;
    buf_clk cell_12053 ( .C (clk), .D (signal_14598), .Q (signal_14599) ) ;
    buf_clk cell_12069 ( .C (clk), .D (signal_14614), .Q (signal_14615) ) ;
    buf_clk cell_12085 ( .C (clk), .D (signal_14630), .Q (signal_14631) ) ;
    buf_clk cell_12101 ( .C (clk), .D (signal_14646), .Q (signal_14647) ) ;
    buf_clk cell_12117 ( .C (clk), .D (signal_14662), .Q (signal_14663) ) ;
    buf_clk cell_12133 ( .C (clk), .D (signal_14678), .Q (signal_14679) ) ;
    buf_clk cell_12149 ( .C (clk), .D (signal_14694), .Q (signal_14695) ) ;
    buf_clk cell_12165 ( .C (clk), .D (signal_14710), .Q (signal_14711) ) ;
    buf_clk cell_12181 ( .C (clk), .D (signal_14726), .Q (signal_14727) ) ;
    buf_clk cell_12197 ( .C (clk), .D (signal_14742), .Q (signal_14743) ) ;
    buf_clk cell_12213 ( .C (clk), .D (signal_14758), .Q (signal_14759) ) ;
    buf_clk cell_12229 ( .C (clk), .D (signal_14774), .Q (signal_14775) ) ;
    buf_clk cell_12245 ( .C (clk), .D (signal_14790), .Q (signal_14791) ) ;
    buf_clk cell_12261 ( .C (clk), .D (signal_14806), .Q (signal_14807) ) ;
    buf_clk cell_12277 ( .C (clk), .D (signal_14822), .Q (signal_14823) ) ;
    buf_clk cell_12293 ( .C (clk), .D (signal_14838), .Q (signal_14839) ) ;
    buf_clk cell_12309 ( .C (clk), .D (signal_14854), .Q (signal_14855) ) ;
    buf_clk cell_12325 ( .C (clk), .D (signal_14870), .Q (signal_14871) ) ;
    buf_clk cell_12341 ( .C (clk), .D (signal_14886), .Q (signal_14887) ) ;
    buf_clk cell_12357 ( .C (clk), .D (signal_14902), .Q (signal_14903) ) ;
    buf_clk cell_12373 ( .C (clk), .D (signal_14918), .Q (signal_14919) ) ;
    buf_clk cell_12389 ( .C (clk), .D (signal_14934), .Q (signal_14935) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2025 ( .s ({signal_4858, signal_4850}), .b ({signal_3700, signal_2173}), .a ({signal_3699, signal_2172}), .clk (clk), .r (Fresh[311]), .c ({signal_3956, signal_2293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2026 ( .s ({signal_4858, signal_4850}), .b ({signal_3702, signal_2175}), .a ({signal_3701, signal_2174}), .clk (clk), .r (Fresh[312]), .c ({signal_3957, signal_2294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2027 ( .s ({signal_4858, signal_4850}), .b ({signal_3704, signal_2177}), .a ({signal_3703, signal_2176}), .clk (clk), .r (Fresh[313]), .c ({signal_3958, signal_2295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2028 ( .s ({signal_4858, signal_4850}), .b ({signal_3706, signal_2179}), .a ({signal_3705, signal_2178}), .clk (clk), .r (Fresh[314]), .c ({signal_3959, signal_2296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2029 ( .s ({signal_4858, signal_4850}), .b ({signal_3707, signal_2180}), .a ({signal_4862, signal_4860}), .clk (clk), .r (Fresh[315]), .c ({signal_3960, signal_2297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2030 ( .s ({signal_4858, signal_4850}), .b ({signal_3709, signal_2182}), .a ({signal_3708, signal_2181}), .clk (clk), .r (Fresh[316]), .c ({signal_3961, signal_2298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2031 ( .s ({signal_4858, signal_4850}), .b ({signal_3710, signal_2183}), .a ({signal_4866, signal_4864}), .clk (clk), .r (Fresh[317]), .c ({signal_3962, signal_2299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2032 ( .s ({signal_4858, signal_4850}), .b ({signal_3711, signal_2184}), .a ({signal_4870, signal_4868}), .clk (clk), .r (Fresh[318]), .c ({signal_3963, signal_2300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2033 ( .s ({signal_4858, signal_4850}), .b ({signal_3713, signal_2186}), .a ({signal_3712, signal_2185}), .clk (clk), .r (Fresh[319]), .c ({signal_3964, signal_2301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2034 ( .s ({signal_4858, signal_4850}), .b ({signal_3715, signal_2188}), .a ({signal_3714, signal_2187}), .clk (clk), .r (Fresh[320]), .c ({signal_3965, signal_2302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2035 ( .s ({signal_4858, signal_4850}), .b ({signal_3717, signal_2190}), .a ({signal_3716, signal_2189}), .clk (clk), .r (Fresh[321]), .c ({signal_3966, signal_2303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2036 ( .s ({signal_4858, signal_4850}), .b ({signal_3719, signal_2192}), .a ({signal_3718, signal_2191}), .clk (clk), .r (Fresh[322]), .c ({signal_3967, signal_2304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2037 ( .s ({signal_4858, signal_4850}), .b ({signal_3721, signal_2194}), .a ({signal_3720, signal_2193}), .clk (clk), .r (Fresh[323]), .c ({signal_3968, signal_2305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2038 ( .s ({signal_4858, signal_4850}), .b ({signal_3723, signal_2196}), .a ({signal_3722, signal_2195}), .clk (clk), .r (Fresh[324]), .c ({signal_3969, signal_2306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2039 ( .s ({signal_4858, signal_4850}), .b ({signal_3725, signal_2198}), .a ({signal_3724, signal_2197}), .clk (clk), .r (Fresh[325]), .c ({signal_3970, signal_2307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2040 ( .s ({signal_4858, signal_4850}), .b ({signal_3727, signal_2200}), .a ({signal_3726, signal_2199}), .clk (clk), .r (Fresh[326]), .c ({signal_3971, signal_2308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2041 ( .s ({signal_4858, signal_4850}), .b ({signal_3729, signal_2202}), .a ({signal_3728, signal_2201}), .clk (clk), .r (Fresh[327]), .c ({signal_3972, signal_2309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2042 ( .s ({signal_4858, signal_4850}), .b ({signal_3731, signal_2204}), .a ({signal_3730, signal_2203}), .clk (clk), .r (Fresh[328]), .c ({signal_3973, signal_2310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2043 ( .s ({signal_4858, signal_4850}), .b ({signal_3733, signal_2206}), .a ({signal_3732, signal_2205}), .clk (clk), .r (Fresh[329]), .c ({signal_3974, signal_2311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2044 ( .s ({signal_4858, signal_4850}), .b ({signal_3735, signal_2208}), .a ({signal_3734, signal_2207}), .clk (clk), .r (Fresh[330]), .c ({signal_3975, signal_2312}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2045 ( .s ({signal_4858, signal_4850}), .b ({signal_3737, signal_2210}), .a ({signal_3736, signal_2209}), .clk (clk), .r (Fresh[331]), .c ({signal_3976, signal_2313}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2046 ( .s ({signal_4858, signal_4850}), .b ({signal_3739, signal_2212}), .a ({signal_3738, signal_2211}), .clk (clk), .r (Fresh[332]), .c ({signal_3977, signal_2314}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2047 ( .s ({signal_4858, signal_4850}), .b ({signal_3741, signal_2214}), .a ({signal_3740, signal_2213}), .clk (clk), .r (Fresh[333]), .c ({signal_3978, signal_2315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2048 ( .s ({signal_4858, signal_4850}), .b ({signal_3743, signal_2216}), .a ({signal_3742, signal_2215}), .clk (clk), .r (Fresh[334]), .c ({signal_3979, signal_2316}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2049 ( .s ({signal_4858, signal_4850}), .b ({signal_3745, signal_2218}), .a ({signal_3744, signal_2217}), .clk (clk), .r (Fresh[335]), .c ({signal_3980, signal_2317}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2050 ( .s ({signal_4858, signal_4850}), .b ({signal_3747, signal_2220}), .a ({signal_3746, signal_2219}), .clk (clk), .r (Fresh[336]), .c ({signal_3981, signal_2318}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2051 ( .s ({signal_4858, signal_4850}), .b ({signal_3748, signal_2221}), .a ({signal_4874, signal_4872}), .clk (clk), .r (Fresh[337]), .c ({signal_3982, signal_2319}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2052 ( .s ({signal_4858, signal_4850}), .b ({signal_3750, signal_2223}), .a ({signal_3749, signal_2222}), .clk (clk), .r (Fresh[338]), .c ({signal_3983, signal_2320}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2053 ( .s ({signal_4858, signal_4850}), .b ({signal_3752, signal_2225}), .a ({signal_3751, signal_2224}), .clk (clk), .r (Fresh[339]), .c ({signal_3984, signal_2321}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2054 ( .s ({signal_4858, signal_4850}), .b ({signal_3754, signal_2227}), .a ({signal_3753, signal_2226}), .clk (clk), .r (Fresh[340]), .c ({signal_3985, signal_2322}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2055 ( .s ({signal_4858, signal_4850}), .b ({signal_3756, signal_2229}), .a ({signal_3755, signal_2228}), .clk (clk), .r (Fresh[341]), .c ({signal_3986, signal_2323}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2056 ( .s ({signal_4858, signal_4850}), .b ({signal_3758, signal_2231}), .a ({signal_3757, signal_2230}), .clk (clk), .r (Fresh[342]), .c ({signal_3987, signal_2324}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2057 ( .s ({signal_4858, signal_4850}), .b ({signal_3760, signal_2233}), .a ({signal_3759, signal_2232}), .clk (clk), .r (Fresh[343]), .c ({signal_3988, signal_2325}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2058 ( .s ({signal_4858, signal_4850}), .b ({signal_4878, signal_4876}), .a ({signal_3761, signal_2234}), .clk (clk), .r (Fresh[344]), .c ({signal_3989, signal_2326}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2059 ( .s ({signal_4858, signal_4850}), .b ({signal_3763, signal_2236}), .a ({signal_3762, signal_2235}), .clk (clk), .r (Fresh[345]), .c ({signal_3990, signal_2327}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2060 ( .s ({signal_4858, signal_4850}), .b ({signal_3765, signal_2238}), .a ({signal_3764, signal_2237}), .clk (clk), .r (Fresh[346]), .c ({signal_3991, signal_2328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2061 ( .s ({signal_4858, signal_4850}), .b ({signal_3767, signal_2240}), .a ({signal_3766, signal_2239}), .clk (clk), .r (Fresh[347]), .c ({signal_3992, signal_2329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2062 ( .s ({signal_4858, signal_4850}), .b ({signal_3769, signal_2242}), .a ({signal_3768, signal_2241}), .clk (clk), .r (Fresh[348]), .c ({signal_3993, signal_2330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2063 ( .s ({signal_4858, signal_4850}), .b ({signal_3771, signal_2244}), .a ({signal_3770, signal_2243}), .clk (clk), .r (Fresh[349]), .c ({signal_3994, signal_2331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2064 ( .s ({signal_4858, signal_4850}), .b ({signal_3773, signal_2246}), .a ({signal_3772, signal_2245}), .clk (clk), .r (Fresh[350]), .c ({signal_3995, signal_2332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2065 ( .s ({signal_4858, signal_4850}), .b ({signal_3775, signal_2248}), .a ({signal_3774, signal_2247}), .clk (clk), .r (Fresh[351]), .c ({signal_3996, signal_2333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2066 ( .s ({signal_4858, signal_4850}), .b ({signal_3777, signal_2250}), .a ({signal_3776, signal_2249}), .clk (clk), .r (Fresh[352]), .c ({signal_3997, signal_2334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2067 ( .s ({signal_4858, signal_4850}), .b ({signal_3779, signal_2252}), .a ({signal_3778, signal_2251}), .clk (clk), .r (Fresh[353]), .c ({signal_3998, signal_2335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2068 ( .s ({signal_4858, signal_4850}), .b ({signal_3781, signal_2254}), .a ({signal_3780, signal_2253}), .clk (clk), .r (Fresh[354]), .c ({signal_3999, signal_2336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2069 ( .s ({signal_4858, signal_4850}), .b ({signal_3783, signal_2256}), .a ({signal_3782, signal_2255}), .clk (clk), .r (Fresh[355]), .c ({signal_4000, signal_2337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2070 ( .s ({signal_4858, signal_4850}), .b ({signal_3785, signal_2258}), .a ({signal_3784, signal_2257}), .clk (clk), .r (Fresh[356]), .c ({signal_4001, signal_2338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2071 ( .s ({signal_4858, signal_4850}), .b ({signal_3787, signal_2260}), .a ({signal_3786, signal_2259}), .clk (clk), .r (Fresh[357]), .c ({signal_4002, signal_2339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2072 ( .s ({signal_4858, signal_4850}), .b ({signal_3789, signal_2262}), .a ({signal_3788, signal_2261}), .clk (clk), .r (Fresh[358]), .c ({signal_4003, signal_2340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2073 ( .s ({signal_4858, signal_4850}), .b ({signal_3791, signal_2264}), .a ({signal_3790, signal_2263}), .clk (clk), .r (Fresh[359]), .c ({signal_4004, signal_2341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2074 ( .s ({signal_4858, signal_4850}), .b ({signal_3792, signal_2265}), .a ({signal_4882, signal_4880}), .clk (clk), .r (Fresh[360]), .c ({signal_4005, signal_2342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2075 ( .s ({signal_4858, signal_4850}), .b ({signal_4886, signal_4884}), .a ({signal_3793, signal_2266}), .clk (clk), .r (Fresh[361]), .c ({signal_4006, signal_2343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2076 ( .s ({signal_4858, signal_4850}), .b ({signal_3795, signal_2268}), .a ({signal_3794, signal_2267}), .clk (clk), .r (Fresh[362]), .c ({signal_4007, signal_2344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2077 ( .s ({signal_4858, signal_4850}), .b ({signal_3797, signal_2270}), .a ({signal_3796, signal_2269}), .clk (clk), .r (Fresh[363]), .c ({signal_4008, signal_2345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2078 ( .s ({signal_4858, signal_4850}), .b ({signal_3799, signal_2272}), .a ({signal_3798, signal_2271}), .clk (clk), .r (Fresh[364]), .c ({signal_4009, signal_2346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2079 ( .s ({signal_4858, signal_4850}), .b ({signal_3801, signal_2274}), .a ({signal_3800, signal_2273}), .clk (clk), .r (Fresh[365]), .c ({signal_4010, signal_2347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2080 ( .s ({signal_4858, signal_4850}), .b ({signal_3803, signal_2276}), .a ({signal_3802, signal_2275}), .clk (clk), .r (Fresh[366]), .c ({signal_4011, signal_2348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2081 ( .s ({signal_4858, signal_4850}), .b ({signal_3805, signal_2278}), .a ({signal_3804, signal_2277}), .clk (clk), .r (Fresh[367]), .c ({signal_4012, signal_2349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2082 ( .s ({signal_4858, signal_4850}), .b ({signal_3807, signal_2280}), .a ({signal_3806, signal_2279}), .clk (clk), .r (Fresh[368]), .c ({signal_4013, signal_2350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2083 ( .s ({signal_4858, signal_4850}), .b ({signal_3809, signal_2282}), .a ({signal_3808, signal_2281}), .clk (clk), .r (Fresh[369]), .c ({signal_4014, signal_2351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2084 ( .s ({signal_4858, signal_4850}), .b ({signal_3811, signal_2284}), .a ({signal_3810, signal_2283}), .clk (clk), .r (Fresh[370]), .c ({signal_4015, signal_2352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2085 ( .s ({signal_4858, signal_4850}), .b ({signal_3813, signal_2286}), .a ({signal_3812, signal_2285}), .clk (clk), .r (Fresh[371]), .c ({signal_4016, signal_2353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2086 ( .s ({signal_4858, signal_4850}), .b ({signal_3815, signal_2288}), .a ({signal_3814, signal_2287}), .clk (clk), .r (Fresh[372]), .c ({signal_4017, signal_2354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2087 ( .s ({signal_4858, signal_4850}), .b ({signal_3817, signal_2290}), .a ({signal_3816, signal_2289}), .clk (clk), .r (Fresh[373]), .c ({signal_4018, signal_2355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2088 ( .s ({signal_4858, signal_4850}), .b ({signal_3819, signal_2292}), .a ({signal_3818, signal_2291}), .clk (clk), .r (Fresh[374]), .c ({signal_4019, signal_2356}) ) ;
    buf_clk cell_2350 ( .C (clk), .D (signal_4895), .Q (signal_4896) ) ;
    buf_clk cell_2360 ( .C (clk), .D (signal_4905), .Q (signal_4906) ) ;
    buf_clk cell_2370 ( .C (clk), .D (signal_4915), .Q (signal_4916) ) ;
    buf_clk cell_2382 ( .C (clk), .D (signal_4927), .Q (signal_4928) ) ;
    buf_clk cell_2394 ( .C (clk), .D (signal_4939), .Q (signal_4940) ) ;
    buf_clk cell_2410 ( .C (clk), .D (signal_4955), .Q (signal_4956) ) ;
    buf_clk cell_2426 ( .C (clk), .D (signal_4971), .Q (signal_4972) ) ;
    buf_clk cell_2442 ( .C (clk), .D (signal_4987), .Q (signal_4988) ) ;
    buf_clk cell_2458 ( .C (clk), .D (signal_5003), .Q (signal_5004) ) ;
    buf_clk cell_2474 ( .C (clk), .D (signal_5019), .Q (signal_5020) ) ;
    buf_clk cell_2490 ( .C (clk), .D (signal_5035), .Q (signal_5036) ) ;
    buf_clk cell_2506 ( .C (clk), .D (signal_5051), .Q (signal_5052) ) ;
    buf_clk cell_2522 ( .C (clk), .D (signal_5067), .Q (signal_5068) ) ;
    buf_clk cell_2538 ( .C (clk), .D (signal_5083), .Q (signal_5084) ) ;
    buf_clk cell_2554 ( .C (clk), .D (signal_5099), .Q (signal_5100) ) ;
    buf_clk cell_2570 ( .C (clk), .D (signal_5115), .Q (signal_5116) ) ;
    buf_clk cell_2586 ( .C (clk), .D (signal_5131), .Q (signal_5132) ) ;
    buf_clk cell_2602 ( .C (clk), .D (signal_5147), .Q (signal_5148) ) ;
    buf_clk cell_2618 ( .C (clk), .D (signal_5163), .Q (signal_5164) ) ;
    buf_clk cell_2634 ( .C (clk), .D (signal_5179), .Q (signal_5180) ) ;
    buf_clk cell_2650 ( .C (clk), .D (signal_5195), .Q (signal_5196) ) ;
    buf_clk cell_2666 ( .C (clk), .D (signal_5211), .Q (signal_5212) ) ;
    buf_clk cell_2682 ( .C (clk), .D (signal_5227), .Q (signal_5228) ) ;
    buf_clk cell_2698 ( .C (clk), .D (signal_5243), .Q (signal_5244) ) ;
    buf_clk cell_2714 ( .C (clk), .D (signal_5259), .Q (signal_5260) ) ;
    buf_clk cell_2730 ( .C (clk), .D (signal_5275), .Q (signal_5276) ) ;
    buf_clk cell_2746 ( .C (clk), .D (signal_5291), .Q (signal_5292) ) ;
    buf_clk cell_2762 ( .C (clk), .D (signal_5307), .Q (signal_5308) ) ;
    buf_clk cell_2778 ( .C (clk), .D (signal_5323), .Q (signal_5324) ) ;
    buf_clk cell_2794 ( .C (clk), .D (signal_5339), .Q (signal_5340) ) ;
    buf_clk cell_2810 ( .C (clk), .D (signal_5355), .Q (signal_5356) ) ;
    buf_clk cell_2826 ( .C (clk), .D (signal_5371), .Q (signal_5372) ) ;
    buf_clk cell_2842 ( .C (clk), .D (signal_5387), .Q (signal_5388) ) ;
    buf_clk cell_2858 ( .C (clk), .D (signal_5403), .Q (signal_5404) ) ;
    buf_clk cell_2874 ( .C (clk), .D (signal_5419), .Q (signal_5420) ) ;
    buf_clk cell_2890 ( .C (clk), .D (signal_5435), .Q (signal_5436) ) ;
    buf_clk cell_2906 ( .C (clk), .D (signal_5451), .Q (signal_5452) ) ;
    buf_clk cell_2922 ( .C (clk), .D (signal_5467), .Q (signal_5468) ) ;
    buf_clk cell_2938 ( .C (clk), .D (signal_5483), .Q (signal_5484) ) ;
    buf_clk cell_2954 ( .C (clk), .D (signal_5499), .Q (signal_5500) ) ;
    buf_clk cell_2970 ( .C (clk), .D (signal_5515), .Q (signal_5516) ) ;
    buf_clk cell_2986 ( .C (clk), .D (signal_5531), .Q (signal_5532) ) ;
    buf_clk cell_3002 ( .C (clk), .D (signal_5547), .Q (signal_5548) ) ;
    buf_clk cell_3018 ( .C (clk), .D (signal_5563), .Q (signal_5564) ) ;
    buf_clk cell_3034 ( .C (clk), .D (signal_5579), .Q (signal_5580) ) ;
    buf_clk cell_3050 ( .C (clk), .D (signal_5595), .Q (signal_5596) ) ;
    buf_clk cell_3066 ( .C (clk), .D (signal_5611), .Q (signal_5612) ) ;
    buf_clk cell_3082 ( .C (clk), .D (signal_5627), .Q (signal_5628) ) ;
    buf_clk cell_3098 ( .C (clk), .D (signal_5643), .Q (signal_5644) ) ;
    buf_clk cell_3114 ( .C (clk), .D (signal_5659), .Q (signal_5660) ) ;
    buf_clk cell_3130 ( .C (clk), .D (signal_5675), .Q (signal_5676) ) ;
    buf_clk cell_3146 ( .C (clk), .D (signal_5691), .Q (signal_5692) ) ;
    buf_clk cell_3162 ( .C (clk), .D (signal_5707), .Q (signal_5708) ) ;
    buf_clk cell_3178 ( .C (clk), .D (signal_5723), .Q (signal_5724) ) ;
    buf_clk cell_3194 ( .C (clk), .D (signal_5739), .Q (signal_5740) ) ;
    buf_clk cell_3210 ( .C (clk), .D (signal_5755), .Q (signal_5756) ) ;
    buf_clk cell_3226 ( .C (clk), .D (signal_5771), .Q (signal_5772) ) ;
    buf_clk cell_3242 ( .C (clk), .D (signal_5787), .Q (signal_5788) ) ;
    buf_clk cell_3258 ( .C (clk), .D (signal_5803), .Q (signal_5804) ) ;
    buf_clk cell_3274 ( .C (clk), .D (signal_5819), .Q (signal_5820) ) ;
    buf_clk cell_3290 ( .C (clk), .D (signal_5835), .Q (signal_5836) ) ;
    buf_clk cell_3306 ( .C (clk), .D (signal_5851), .Q (signal_5852) ) ;
    buf_clk cell_3322 ( .C (clk), .D (signal_5867), .Q (signal_5868) ) ;
    buf_clk cell_3338 ( .C (clk), .D (signal_5883), .Q (signal_5884) ) ;
    buf_clk cell_3354 ( .C (clk), .D (signal_5899), .Q (signal_5900) ) ;
    buf_clk cell_3370 ( .C (clk), .D (signal_5915), .Q (signal_5916) ) ;
    buf_clk cell_3386 ( .C (clk), .D (signal_5931), .Q (signal_5932) ) ;
    buf_clk cell_3402 ( .C (clk), .D (signal_5947), .Q (signal_5948) ) ;
    buf_clk cell_3418 ( .C (clk), .D (signal_5963), .Q (signal_5964) ) ;
    buf_clk cell_3434 ( .C (clk), .D (signal_5979), .Q (signal_5980) ) ;
    buf_clk cell_3450 ( .C (clk), .D (signal_5995), .Q (signal_5996) ) ;
    buf_clk cell_3466 ( .C (clk), .D (signal_6011), .Q (signal_6012) ) ;
    buf_clk cell_3482 ( .C (clk), .D (signal_6027), .Q (signal_6028) ) ;
    buf_clk cell_3498 ( .C (clk), .D (signal_6043), .Q (signal_6044) ) ;
    buf_clk cell_3514 ( .C (clk), .D (signal_6059), .Q (signal_6060) ) ;
    buf_clk cell_3530 ( .C (clk), .D (signal_6075), .Q (signal_6076) ) ;
    buf_clk cell_3546 ( .C (clk), .D (signal_6091), .Q (signal_6092) ) ;
    buf_clk cell_3562 ( .C (clk), .D (signal_6107), .Q (signal_6108) ) ;
    buf_clk cell_3578 ( .C (clk), .D (signal_6123), .Q (signal_6124) ) ;
    buf_clk cell_3594 ( .C (clk), .D (signal_6139), .Q (signal_6140) ) ;
    buf_clk cell_3610 ( .C (clk), .D (signal_6155), .Q (signal_6156) ) ;
    buf_clk cell_3626 ( .C (clk), .D (signal_6171), .Q (signal_6172) ) ;
    buf_clk cell_3642 ( .C (clk), .D (signal_6187), .Q (signal_6188) ) ;
    buf_clk cell_3658 ( .C (clk), .D (signal_6203), .Q (signal_6204) ) ;
    buf_clk cell_3674 ( .C (clk), .D (signal_6219), .Q (signal_6220) ) ;
    buf_clk cell_3690 ( .C (clk), .D (signal_6235), .Q (signal_6236) ) ;
    buf_clk cell_3706 ( .C (clk), .D (signal_6251), .Q (signal_6252) ) ;
    buf_clk cell_3722 ( .C (clk), .D (signal_6267), .Q (signal_6268) ) ;
    buf_clk cell_3738 ( .C (clk), .D (signal_6283), .Q (signal_6284) ) ;
    buf_clk cell_3754 ( .C (clk), .D (signal_6299), .Q (signal_6300) ) ;
    buf_clk cell_3770 ( .C (clk), .D (signal_6315), .Q (signal_6316) ) ;
    buf_clk cell_3786 ( .C (clk), .D (signal_6331), .Q (signal_6332) ) ;
    buf_clk cell_3802 ( .C (clk), .D (signal_6347), .Q (signal_6348) ) ;
    buf_clk cell_3818 ( .C (clk), .D (signal_6363), .Q (signal_6364) ) ;
    buf_clk cell_3834 ( .C (clk), .D (signal_6379), .Q (signal_6380) ) ;
    buf_clk cell_3850 ( .C (clk), .D (signal_6395), .Q (signal_6396) ) ;
    buf_clk cell_3866 ( .C (clk), .D (signal_6411), .Q (signal_6412) ) ;
    buf_clk cell_3882 ( .C (clk), .D (signal_6427), .Q (signal_6428) ) ;
    buf_clk cell_3898 ( .C (clk), .D (signal_6443), .Q (signal_6444) ) ;
    buf_clk cell_3914 ( .C (clk), .D (signal_6459), .Q (signal_6460) ) ;
    buf_clk cell_3930 ( .C (clk), .D (signal_6475), .Q (signal_6476) ) ;
    buf_clk cell_3946 ( .C (clk), .D (signal_6491), .Q (signal_6492) ) ;
    buf_clk cell_3962 ( .C (clk), .D (signal_6507), .Q (signal_6508) ) ;
    buf_clk cell_3978 ( .C (clk), .D (signal_6523), .Q (signal_6524) ) ;
    buf_clk cell_3994 ( .C (clk), .D (signal_6539), .Q (signal_6540) ) ;
    buf_clk cell_4010 ( .C (clk), .D (signal_6555), .Q (signal_6556) ) ;
    buf_clk cell_4026 ( .C (clk), .D (signal_6571), .Q (signal_6572) ) ;
    buf_clk cell_4042 ( .C (clk), .D (signal_6587), .Q (signal_6588) ) ;
    buf_clk cell_4058 ( .C (clk), .D (signal_6603), .Q (signal_6604) ) ;
    buf_clk cell_4074 ( .C (clk), .D (signal_6619), .Q (signal_6620) ) ;
    buf_clk cell_4090 ( .C (clk), .D (signal_6635), .Q (signal_6636) ) ;
    buf_clk cell_4106 ( .C (clk), .D (signal_6651), .Q (signal_6652) ) ;
    buf_clk cell_4122 ( .C (clk), .D (signal_6667), .Q (signal_6668) ) ;
    buf_clk cell_4138 ( .C (clk), .D (signal_6683), .Q (signal_6684) ) ;
    buf_clk cell_4154 ( .C (clk), .D (signal_6699), .Q (signal_6700) ) ;
    buf_clk cell_4170 ( .C (clk), .D (signal_6715), .Q (signal_6716) ) ;
    buf_clk cell_4186 ( .C (clk), .D (signal_6731), .Q (signal_6732) ) ;
    buf_clk cell_4202 ( .C (clk), .D (signal_6747), .Q (signal_6748) ) ;
    buf_clk cell_4218 ( .C (clk), .D (signal_6763), .Q (signal_6764) ) ;
    buf_clk cell_4234 ( .C (clk), .D (signal_6779), .Q (signal_6780) ) ;
    buf_clk cell_4250 ( .C (clk), .D (signal_6795), .Q (signal_6796) ) ;
    buf_clk cell_4266 ( .C (clk), .D (signal_6811), .Q (signal_6812) ) ;
    buf_clk cell_4282 ( .C (clk), .D (signal_6827), .Q (signal_6828) ) ;
    buf_clk cell_4298 ( .C (clk), .D (signal_6843), .Q (signal_6844) ) ;
    buf_clk cell_4314 ( .C (clk), .D (signal_6859), .Q (signal_6860) ) ;
    buf_clk cell_4330 ( .C (clk), .D (signal_6875), .Q (signal_6876) ) ;
    buf_clk cell_4346 ( .C (clk), .D (signal_6891), .Q (signal_6892) ) ;
    buf_clk cell_4362 ( .C (clk), .D (signal_6907), .Q (signal_6908) ) ;
    buf_clk cell_4378 ( .C (clk), .D (signal_6923), .Q (signal_6924) ) ;
    buf_clk cell_4394 ( .C (clk), .D (signal_6939), .Q (signal_6940) ) ;
    buf_clk cell_4410 ( .C (clk), .D (signal_6955), .Q (signal_6956) ) ;
    buf_clk cell_4424 ( .C (clk), .D (signal_6969), .Q (signal_6970) ) ;
    buf_clk cell_4438 ( .C (clk), .D (signal_6983), .Q (signal_6984) ) ;
    buf_clk cell_4454 ( .C (clk), .D (signal_6999), .Q (signal_7000) ) ;
    buf_clk cell_4470 ( .C (clk), .D (signal_7015), .Q (signal_7016) ) ;
    buf_clk cell_4486 ( .C (clk), .D (signal_7031), .Q (signal_7032) ) ;
    buf_clk cell_4502 ( .C (clk), .D (signal_7047), .Q (signal_7048) ) ;
    buf_clk cell_4518 ( .C (clk), .D (signal_7063), .Q (signal_7064) ) ;
    buf_clk cell_4534 ( .C (clk), .D (signal_7079), .Q (signal_7080) ) ;
    buf_clk cell_4550 ( .C (clk), .D (signal_7095), .Q (signal_7096) ) ;
    buf_clk cell_4566 ( .C (clk), .D (signal_7111), .Q (signal_7112) ) ;
    buf_clk cell_4582 ( .C (clk), .D (signal_7127), .Q (signal_7128) ) ;
    buf_clk cell_4598 ( .C (clk), .D (signal_7143), .Q (signal_7144) ) ;
    buf_clk cell_4614 ( .C (clk), .D (signal_7159), .Q (signal_7160) ) ;
    buf_clk cell_4630 ( .C (clk), .D (signal_7175), .Q (signal_7176) ) ;
    buf_clk cell_4646 ( .C (clk), .D (signal_7191), .Q (signal_7192) ) ;
    buf_clk cell_4662 ( .C (clk), .D (signal_7207), .Q (signal_7208) ) ;
    buf_clk cell_4678 ( .C (clk), .D (signal_7223), .Q (signal_7224) ) ;
    buf_clk cell_4694 ( .C (clk), .D (signal_7239), .Q (signal_7240) ) ;
    buf_clk cell_4710 ( .C (clk), .D (signal_7255), .Q (signal_7256) ) ;
    buf_clk cell_4726 ( .C (clk), .D (signal_7271), .Q (signal_7272) ) ;
    buf_clk cell_4742 ( .C (clk), .D (signal_7287), .Q (signal_7288) ) ;
    buf_clk cell_4758 ( .C (clk), .D (signal_7303), .Q (signal_7304) ) ;
    buf_clk cell_4774 ( .C (clk), .D (signal_7319), .Q (signal_7320) ) ;
    buf_clk cell_4790 ( .C (clk), .D (signal_7335), .Q (signal_7336) ) ;
    buf_clk cell_4806 ( .C (clk), .D (signal_7351), .Q (signal_7352) ) ;
    buf_clk cell_4822 ( .C (clk), .D (signal_7367), .Q (signal_7368) ) ;
    buf_clk cell_4838 ( .C (clk), .D (signal_7383), .Q (signal_7384) ) ;
    buf_clk cell_4854 ( .C (clk), .D (signal_7399), .Q (signal_7400) ) ;
    buf_clk cell_4870 ( .C (clk), .D (signal_7415), .Q (signal_7416) ) ;
    buf_clk cell_4886 ( .C (clk), .D (signal_7431), .Q (signal_7432) ) ;
    buf_clk cell_4902 ( .C (clk), .D (signal_7447), .Q (signal_7448) ) ;
    buf_clk cell_4918 ( .C (clk), .D (signal_7463), .Q (signal_7464) ) ;
    buf_clk cell_4934 ( .C (clk), .D (signal_7479), .Q (signal_7480) ) ;
    buf_clk cell_4950 ( .C (clk), .D (signal_7495), .Q (signal_7496) ) ;
    buf_clk cell_4966 ( .C (clk), .D (signal_7511), .Q (signal_7512) ) ;
    buf_clk cell_4982 ( .C (clk), .D (signal_7527), .Q (signal_7528) ) ;
    buf_clk cell_4998 ( .C (clk), .D (signal_7543), .Q (signal_7544) ) ;
    buf_clk cell_5014 ( .C (clk), .D (signal_7559), .Q (signal_7560) ) ;
    buf_clk cell_5030 ( .C (clk), .D (signal_7575), .Q (signal_7576) ) ;
    buf_clk cell_5046 ( .C (clk), .D (signal_7591), .Q (signal_7592) ) ;
    buf_clk cell_5062 ( .C (clk), .D (signal_7607), .Q (signal_7608) ) ;
    buf_clk cell_5078 ( .C (clk), .D (signal_7623), .Q (signal_7624) ) ;
    buf_clk cell_5094 ( .C (clk), .D (signal_7639), .Q (signal_7640) ) ;
    buf_clk cell_5110 ( .C (clk), .D (signal_7655), .Q (signal_7656) ) ;
    buf_clk cell_5126 ( .C (clk), .D (signal_7671), .Q (signal_7672) ) ;
    buf_clk cell_5142 ( .C (clk), .D (signal_7687), .Q (signal_7688) ) ;
    buf_clk cell_5158 ( .C (clk), .D (signal_7703), .Q (signal_7704) ) ;
    buf_clk cell_5174 ( .C (clk), .D (signal_7719), .Q (signal_7720) ) ;
    buf_clk cell_5190 ( .C (clk), .D (signal_7735), .Q (signal_7736) ) ;
    buf_clk cell_5206 ( .C (clk), .D (signal_7751), .Q (signal_7752) ) ;
    buf_clk cell_5222 ( .C (clk), .D (signal_7767), .Q (signal_7768) ) ;
    buf_clk cell_5238 ( .C (clk), .D (signal_7783), .Q (signal_7784) ) ;
    buf_clk cell_5254 ( .C (clk), .D (signal_7799), .Q (signal_7800) ) ;
    buf_clk cell_5270 ( .C (clk), .D (signal_7815), .Q (signal_7816) ) ;
    buf_clk cell_5286 ( .C (clk), .D (signal_7831), .Q (signal_7832) ) ;
    buf_clk cell_5302 ( .C (clk), .D (signal_7847), .Q (signal_7848) ) ;
    buf_clk cell_5318 ( .C (clk), .D (signal_7863), .Q (signal_7864) ) ;
    buf_clk cell_5334 ( .C (clk), .D (signal_7879), .Q (signal_7880) ) ;
    buf_clk cell_5350 ( .C (clk), .D (signal_7895), .Q (signal_7896) ) ;
    buf_clk cell_5366 ( .C (clk), .D (signal_7911), .Q (signal_7912) ) ;
    buf_clk cell_5382 ( .C (clk), .D (signal_7927), .Q (signal_7928) ) ;
    buf_clk cell_5398 ( .C (clk), .D (signal_7943), .Q (signal_7944) ) ;
    buf_clk cell_5414 ( .C (clk), .D (signal_7959), .Q (signal_7960) ) ;
    buf_clk cell_5430 ( .C (clk), .D (signal_7975), .Q (signal_7976) ) ;
    buf_clk cell_5446 ( .C (clk), .D (signal_7991), .Q (signal_7992) ) ;
    buf_clk cell_5462 ( .C (clk), .D (signal_8007), .Q (signal_8008) ) ;
    buf_clk cell_5478 ( .C (clk), .D (signal_8023), .Q (signal_8024) ) ;
    buf_clk cell_5494 ( .C (clk), .D (signal_8039), .Q (signal_8040) ) ;
    buf_clk cell_5510 ( .C (clk), .D (signal_8055), .Q (signal_8056) ) ;
    buf_clk cell_5526 ( .C (clk), .D (signal_8071), .Q (signal_8072) ) ;
    buf_clk cell_5542 ( .C (clk), .D (signal_8087), .Q (signal_8088) ) ;
    buf_clk cell_5558 ( .C (clk), .D (signal_8103), .Q (signal_8104) ) ;
    buf_clk cell_5574 ( .C (clk), .D (signal_8119), .Q (signal_8120) ) ;
    buf_clk cell_5590 ( .C (clk), .D (signal_8135), .Q (signal_8136) ) ;
    buf_clk cell_5606 ( .C (clk), .D (signal_8151), .Q (signal_8152) ) ;
    buf_clk cell_5622 ( .C (clk), .D (signal_8167), .Q (signal_8168) ) ;
    buf_clk cell_5638 ( .C (clk), .D (signal_8183), .Q (signal_8184) ) ;
    buf_clk cell_5654 ( .C (clk), .D (signal_8199), .Q (signal_8200) ) ;
    buf_clk cell_5670 ( .C (clk), .D (signal_8215), .Q (signal_8216) ) ;
    buf_clk cell_5686 ( .C (clk), .D (signal_8231), .Q (signal_8232) ) ;
    buf_clk cell_5702 ( .C (clk), .D (signal_8247), .Q (signal_8248) ) ;
    buf_clk cell_5718 ( .C (clk), .D (signal_8263), .Q (signal_8264) ) ;
    buf_clk cell_5734 ( .C (clk), .D (signal_8279), .Q (signal_8280) ) ;
    buf_clk cell_5750 ( .C (clk), .D (signal_8295), .Q (signal_8296) ) ;
    buf_clk cell_5766 ( .C (clk), .D (signal_8311), .Q (signal_8312) ) ;
    buf_clk cell_5782 ( .C (clk), .D (signal_8327), .Q (signal_8328) ) ;
    buf_clk cell_5798 ( .C (clk), .D (signal_8343), .Q (signal_8344) ) ;
    buf_clk cell_5814 ( .C (clk), .D (signal_8359), .Q (signal_8360) ) ;
    buf_clk cell_5830 ( .C (clk), .D (signal_8375), .Q (signal_8376) ) ;
    buf_clk cell_5846 ( .C (clk), .D (signal_8391), .Q (signal_8392) ) ;
    buf_clk cell_5862 ( .C (clk), .D (signal_8407), .Q (signal_8408) ) ;
    buf_clk cell_5878 ( .C (clk), .D (signal_8423), .Q (signal_8424) ) ;
    buf_clk cell_5894 ( .C (clk), .D (signal_8439), .Q (signal_8440) ) ;
    buf_clk cell_5910 ( .C (clk), .D (signal_8455), .Q (signal_8456) ) ;
    buf_clk cell_5926 ( .C (clk), .D (signal_8471), .Q (signal_8472) ) ;
    buf_clk cell_5942 ( .C (clk), .D (signal_8487), .Q (signal_8488) ) ;
    buf_clk cell_5958 ( .C (clk), .D (signal_8503), .Q (signal_8504) ) ;
    buf_clk cell_5974 ( .C (clk), .D (signal_8519), .Q (signal_8520) ) ;
    buf_clk cell_5990 ( .C (clk), .D (signal_8535), .Q (signal_8536) ) ;
    buf_clk cell_6006 ( .C (clk), .D (signal_8551), .Q (signal_8552) ) ;
    buf_clk cell_6022 ( .C (clk), .D (signal_8567), .Q (signal_8568) ) ;
    buf_clk cell_6038 ( .C (clk), .D (signal_8583), .Q (signal_8584) ) ;
    buf_clk cell_6054 ( .C (clk), .D (signal_8599), .Q (signal_8600) ) ;
    buf_clk cell_6070 ( .C (clk), .D (signal_8615), .Q (signal_8616) ) ;
    buf_clk cell_6086 ( .C (clk), .D (signal_8631), .Q (signal_8632) ) ;
    buf_clk cell_6102 ( .C (clk), .D (signal_8647), .Q (signal_8648) ) ;
    buf_clk cell_6118 ( .C (clk), .D (signal_8663), .Q (signal_8664) ) ;
    buf_clk cell_6134 ( .C (clk), .D (signal_8679), .Q (signal_8680) ) ;
    buf_clk cell_6150 ( .C (clk), .D (signal_8695), .Q (signal_8696) ) ;
    buf_clk cell_6166 ( .C (clk), .D (signal_8711), .Q (signal_8712) ) ;
    buf_clk cell_6182 ( .C (clk), .D (signal_8727), .Q (signal_8728) ) ;
    buf_clk cell_6198 ( .C (clk), .D (signal_8743), .Q (signal_8744) ) ;
    buf_clk cell_6214 ( .C (clk), .D (signal_8759), .Q (signal_8760) ) ;
    buf_clk cell_6230 ( .C (clk), .D (signal_8775), .Q (signal_8776) ) ;
    buf_clk cell_6246 ( .C (clk), .D (signal_8791), .Q (signal_8792) ) ;
    buf_clk cell_6262 ( .C (clk), .D (signal_8807), .Q (signal_8808) ) ;
    buf_clk cell_6278 ( .C (clk), .D (signal_8823), .Q (signal_8824) ) ;
    buf_clk cell_6294 ( .C (clk), .D (signal_8839), .Q (signal_8840) ) ;
    buf_clk cell_6310 ( .C (clk), .D (signal_8855), .Q (signal_8856) ) ;
    buf_clk cell_6326 ( .C (clk), .D (signal_8871), .Q (signal_8872) ) ;
    buf_clk cell_6342 ( .C (clk), .D (signal_8887), .Q (signal_8888) ) ;
    buf_clk cell_6358 ( .C (clk), .D (signal_8903), .Q (signal_8904) ) ;
    buf_clk cell_6374 ( .C (clk), .D (signal_8919), .Q (signal_8920) ) ;
    buf_clk cell_6390 ( .C (clk), .D (signal_8935), .Q (signal_8936) ) ;
    buf_clk cell_6406 ( .C (clk), .D (signal_8951), .Q (signal_8952) ) ;
    buf_clk cell_6422 ( .C (clk), .D (signal_8967), .Q (signal_8968) ) ;
    buf_clk cell_6438 ( .C (clk), .D (signal_8983), .Q (signal_8984) ) ;
    buf_clk cell_6454 ( .C (clk), .D (signal_8999), .Q (signal_9000) ) ;
    buf_clk cell_6470 ( .C (clk), .D (signal_9015), .Q (signal_9016) ) ;
    buf_clk cell_6486 ( .C (clk), .D (signal_9031), .Q (signal_9032) ) ;
    buf_clk cell_6502 ( .C (clk), .D (signal_9047), .Q (signal_9048) ) ;
    buf_clk cell_6518 ( .C (clk), .D (signal_9063), .Q (signal_9064) ) ;
    buf_clk cell_6534 ( .C (clk), .D (signal_9079), .Q (signal_9080) ) ;
    buf_clk cell_6550 ( .C (clk), .D (signal_9095), .Q (signal_9096) ) ;
    buf_clk cell_6566 ( .C (clk), .D (signal_9111), .Q (signal_9112) ) ;
    buf_clk cell_6582 ( .C (clk), .D (signal_9127), .Q (signal_9128) ) ;
    buf_clk cell_6598 ( .C (clk), .D (signal_9143), .Q (signal_9144) ) ;
    buf_clk cell_6614 ( .C (clk), .D (signal_9159), .Q (signal_9160) ) ;
    buf_clk cell_6630 ( .C (clk), .D (signal_9175), .Q (signal_9176) ) ;
    buf_clk cell_6646 ( .C (clk), .D (signal_9191), .Q (signal_9192) ) ;
    buf_clk cell_6662 ( .C (clk), .D (signal_9207), .Q (signal_9208) ) ;
    buf_clk cell_6678 ( .C (clk), .D (signal_9223), .Q (signal_9224) ) ;
    buf_clk cell_6694 ( .C (clk), .D (signal_9239), .Q (signal_9240) ) ;
    buf_clk cell_6710 ( .C (clk), .D (signal_9255), .Q (signal_9256) ) ;
    buf_clk cell_6726 ( .C (clk), .D (signal_9271), .Q (signal_9272) ) ;
    buf_clk cell_6742 ( .C (clk), .D (signal_9287), .Q (signal_9288) ) ;
    buf_clk cell_6758 ( .C (clk), .D (signal_9303), .Q (signal_9304) ) ;
    buf_clk cell_6774 ( .C (clk), .D (signal_9319), .Q (signal_9320) ) ;
    buf_clk cell_6790 ( .C (clk), .D (signal_9335), .Q (signal_9336) ) ;
    buf_clk cell_6806 ( .C (clk), .D (signal_9351), .Q (signal_9352) ) ;
    buf_clk cell_6822 ( .C (clk), .D (signal_9367), .Q (signal_9368) ) ;
    buf_clk cell_6838 ( .C (clk), .D (signal_9383), .Q (signal_9384) ) ;
    buf_clk cell_6854 ( .C (clk), .D (signal_9399), .Q (signal_9400) ) ;
    buf_clk cell_6870 ( .C (clk), .D (signal_9415), .Q (signal_9416) ) ;
    buf_clk cell_6886 ( .C (clk), .D (signal_9431), .Q (signal_9432) ) ;
    buf_clk cell_6902 ( .C (clk), .D (signal_9447), .Q (signal_9448) ) ;
    buf_clk cell_6918 ( .C (clk), .D (signal_9463), .Q (signal_9464) ) ;
    buf_clk cell_6934 ( .C (clk), .D (signal_9479), .Q (signal_9480) ) ;
    buf_clk cell_6950 ( .C (clk), .D (signal_9495), .Q (signal_9496) ) ;
    buf_clk cell_6966 ( .C (clk), .D (signal_9511), .Q (signal_9512) ) ;
    buf_clk cell_6982 ( .C (clk), .D (signal_9527), .Q (signal_9528) ) ;
    buf_clk cell_6998 ( .C (clk), .D (signal_9543), .Q (signal_9544) ) ;
    buf_clk cell_7014 ( .C (clk), .D (signal_9559), .Q (signal_9560) ) ;
    buf_clk cell_7030 ( .C (clk), .D (signal_9575), .Q (signal_9576) ) ;
    buf_clk cell_7046 ( .C (clk), .D (signal_9591), .Q (signal_9592) ) ;
    buf_clk cell_7062 ( .C (clk), .D (signal_9607), .Q (signal_9608) ) ;
    buf_clk cell_7078 ( .C (clk), .D (signal_9623), .Q (signal_9624) ) ;
    buf_clk cell_7094 ( .C (clk), .D (signal_9639), .Q (signal_9640) ) ;
    buf_clk cell_7110 ( .C (clk), .D (signal_9655), .Q (signal_9656) ) ;
    buf_clk cell_7126 ( .C (clk), .D (signal_9671), .Q (signal_9672) ) ;
    buf_clk cell_7142 ( .C (clk), .D (signal_9687), .Q (signal_9688) ) ;
    buf_clk cell_7158 ( .C (clk), .D (signal_9703), .Q (signal_9704) ) ;
    buf_clk cell_7174 ( .C (clk), .D (signal_9719), .Q (signal_9720) ) ;
    buf_clk cell_7190 ( .C (clk), .D (signal_9735), .Q (signal_9736) ) ;
    buf_clk cell_7206 ( .C (clk), .D (signal_9751), .Q (signal_9752) ) ;
    buf_clk cell_7222 ( .C (clk), .D (signal_9767), .Q (signal_9768) ) ;
    buf_clk cell_7238 ( .C (clk), .D (signal_9783), .Q (signal_9784) ) ;
    buf_clk cell_7254 ( .C (clk), .D (signal_9799), .Q (signal_9800) ) ;
    buf_clk cell_7270 ( .C (clk), .D (signal_9815), .Q (signal_9816) ) ;
    buf_clk cell_7286 ( .C (clk), .D (signal_9831), .Q (signal_9832) ) ;
    buf_clk cell_7302 ( .C (clk), .D (signal_9847), .Q (signal_9848) ) ;
    buf_clk cell_7318 ( .C (clk), .D (signal_9863), .Q (signal_9864) ) ;
    buf_clk cell_7334 ( .C (clk), .D (signal_9879), .Q (signal_9880) ) ;
    buf_clk cell_7350 ( .C (clk), .D (signal_9895), .Q (signal_9896) ) ;
    buf_clk cell_7366 ( .C (clk), .D (signal_9911), .Q (signal_9912) ) ;
    buf_clk cell_7382 ( .C (clk), .D (signal_9927), .Q (signal_9928) ) ;
    buf_clk cell_7398 ( .C (clk), .D (signal_9943), .Q (signal_9944) ) ;
    buf_clk cell_7414 ( .C (clk), .D (signal_9959), .Q (signal_9960) ) ;
    buf_clk cell_7430 ( .C (clk), .D (signal_9975), .Q (signal_9976) ) ;
    buf_clk cell_7446 ( .C (clk), .D (signal_9991), .Q (signal_9992) ) ;
    buf_clk cell_7462 ( .C (clk), .D (signal_10007), .Q (signal_10008) ) ;
    buf_clk cell_7478 ( .C (clk), .D (signal_10023), .Q (signal_10024) ) ;
    buf_clk cell_7494 ( .C (clk), .D (signal_10039), .Q (signal_10040) ) ;
    buf_clk cell_7510 ( .C (clk), .D (signal_10055), .Q (signal_10056) ) ;
    buf_clk cell_7526 ( .C (clk), .D (signal_10071), .Q (signal_10072) ) ;
    buf_clk cell_7542 ( .C (clk), .D (signal_10087), .Q (signal_10088) ) ;
    buf_clk cell_7558 ( .C (clk), .D (signal_10103), .Q (signal_10104) ) ;
    buf_clk cell_7574 ( .C (clk), .D (signal_10119), .Q (signal_10120) ) ;
    buf_clk cell_7590 ( .C (clk), .D (signal_10135), .Q (signal_10136) ) ;
    buf_clk cell_7606 ( .C (clk), .D (signal_10151), .Q (signal_10152) ) ;
    buf_clk cell_7622 ( .C (clk), .D (signal_10167), .Q (signal_10168) ) ;
    buf_clk cell_7638 ( .C (clk), .D (signal_10183), .Q (signal_10184) ) ;
    buf_clk cell_7654 ( .C (clk), .D (signal_10199), .Q (signal_10200) ) ;
    buf_clk cell_7670 ( .C (clk), .D (signal_10215), .Q (signal_10216) ) ;
    buf_clk cell_7686 ( .C (clk), .D (signal_10231), .Q (signal_10232) ) ;
    buf_clk cell_7702 ( .C (clk), .D (signal_10247), .Q (signal_10248) ) ;
    buf_clk cell_7718 ( .C (clk), .D (signal_10263), .Q (signal_10264) ) ;
    buf_clk cell_7734 ( .C (clk), .D (signal_10279), .Q (signal_10280) ) ;
    buf_clk cell_7750 ( .C (clk), .D (signal_10295), .Q (signal_10296) ) ;
    buf_clk cell_7766 ( .C (clk), .D (signal_10311), .Q (signal_10312) ) ;
    buf_clk cell_7782 ( .C (clk), .D (signal_10327), .Q (signal_10328) ) ;
    buf_clk cell_7798 ( .C (clk), .D (signal_10343), .Q (signal_10344) ) ;
    buf_clk cell_7814 ( .C (clk), .D (signal_10359), .Q (signal_10360) ) ;
    buf_clk cell_7830 ( .C (clk), .D (signal_10375), .Q (signal_10376) ) ;
    buf_clk cell_7846 ( .C (clk), .D (signal_10391), .Q (signal_10392) ) ;
    buf_clk cell_7862 ( .C (clk), .D (signal_10407), .Q (signal_10408) ) ;
    buf_clk cell_7878 ( .C (clk), .D (signal_10423), .Q (signal_10424) ) ;
    buf_clk cell_7894 ( .C (clk), .D (signal_10439), .Q (signal_10440) ) ;
    buf_clk cell_7910 ( .C (clk), .D (signal_10455), .Q (signal_10456) ) ;
    buf_clk cell_7926 ( .C (clk), .D (signal_10471), .Q (signal_10472) ) ;
    buf_clk cell_7942 ( .C (clk), .D (signal_10487), .Q (signal_10488) ) ;
    buf_clk cell_7958 ( .C (clk), .D (signal_10503), .Q (signal_10504) ) ;
    buf_clk cell_7974 ( .C (clk), .D (signal_10519), .Q (signal_10520) ) ;
    buf_clk cell_7990 ( .C (clk), .D (signal_10535), .Q (signal_10536) ) ;
    buf_clk cell_8006 ( .C (clk), .D (signal_10551), .Q (signal_10552) ) ;
    buf_clk cell_8022 ( .C (clk), .D (signal_10567), .Q (signal_10568) ) ;
    buf_clk cell_8038 ( .C (clk), .D (signal_10583), .Q (signal_10584) ) ;
    buf_clk cell_8054 ( .C (clk), .D (signal_10599), .Q (signal_10600) ) ;
    buf_clk cell_8070 ( .C (clk), .D (signal_10615), .Q (signal_10616) ) ;
    buf_clk cell_8086 ( .C (clk), .D (signal_10631), .Q (signal_10632) ) ;
    buf_clk cell_8102 ( .C (clk), .D (signal_10647), .Q (signal_10648) ) ;
    buf_clk cell_8118 ( .C (clk), .D (signal_10663), .Q (signal_10664) ) ;
    buf_clk cell_8134 ( .C (clk), .D (signal_10679), .Q (signal_10680) ) ;
    buf_clk cell_8150 ( .C (clk), .D (signal_10695), .Q (signal_10696) ) ;
    buf_clk cell_8166 ( .C (clk), .D (signal_10711), .Q (signal_10712) ) ;
    buf_clk cell_8182 ( .C (clk), .D (signal_10727), .Q (signal_10728) ) ;
    buf_clk cell_8198 ( .C (clk), .D (signal_10743), .Q (signal_10744) ) ;
    buf_clk cell_8214 ( .C (clk), .D (signal_10759), .Q (signal_10760) ) ;
    buf_clk cell_8230 ( .C (clk), .D (signal_10775), .Q (signal_10776) ) ;
    buf_clk cell_8246 ( .C (clk), .D (signal_10791), .Q (signal_10792) ) ;
    buf_clk cell_8262 ( .C (clk), .D (signal_10807), .Q (signal_10808) ) ;
    buf_clk cell_8278 ( .C (clk), .D (signal_10823), .Q (signal_10824) ) ;
    buf_clk cell_8294 ( .C (clk), .D (signal_10839), .Q (signal_10840) ) ;
    buf_clk cell_8310 ( .C (clk), .D (signal_10855), .Q (signal_10856) ) ;
    buf_clk cell_8326 ( .C (clk), .D (signal_10871), .Q (signal_10872) ) ;
    buf_clk cell_8342 ( .C (clk), .D (signal_10887), .Q (signal_10888) ) ;
    buf_clk cell_8358 ( .C (clk), .D (signal_10903), .Q (signal_10904) ) ;
    buf_clk cell_8374 ( .C (clk), .D (signal_10919), .Q (signal_10920) ) ;
    buf_clk cell_8390 ( .C (clk), .D (signal_10935), .Q (signal_10936) ) ;
    buf_clk cell_8406 ( .C (clk), .D (signal_10951), .Q (signal_10952) ) ;
    buf_clk cell_8422 ( .C (clk), .D (signal_10967), .Q (signal_10968) ) ;
    buf_clk cell_8438 ( .C (clk), .D (signal_10983), .Q (signal_10984) ) ;
    buf_clk cell_8454 ( .C (clk), .D (signal_10999), .Q (signal_11000) ) ;
    buf_clk cell_8470 ( .C (clk), .D (signal_11015), .Q (signal_11016) ) ;
    buf_clk cell_8486 ( .C (clk), .D (signal_11031), .Q (signal_11032) ) ;
    buf_clk cell_8502 ( .C (clk), .D (signal_11047), .Q (signal_11048) ) ;
    buf_clk cell_8518 ( .C (clk), .D (signal_11063), .Q (signal_11064) ) ;
    buf_clk cell_8534 ( .C (clk), .D (signal_11079), .Q (signal_11080) ) ;
    buf_clk cell_8550 ( .C (clk), .D (signal_11095), .Q (signal_11096) ) ;
    buf_clk cell_8566 ( .C (clk), .D (signal_11111), .Q (signal_11112) ) ;
    buf_clk cell_8582 ( .C (clk), .D (signal_11127), .Q (signal_11128) ) ;
    buf_clk cell_8598 ( .C (clk), .D (signal_11143), .Q (signal_11144) ) ;
    buf_clk cell_8614 ( .C (clk), .D (signal_11159), .Q (signal_11160) ) ;
    buf_clk cell_8630 ( .C (clk), .D (signal_11175), .Q (signal_11176) ) ;
    buf_clk cell_8646 ( .C (clk), .D (signal_11191), .Q (signal_11192) ) ;
    buf_clk cell_8662 ( .C (clk), .D (signal_11207), .Q (signal_11208) ) ;
    buf_clk cell_8678 ( .C (clk), .D (signal_11223), .Q (signal_11224) ) ;
    buf_clk cell_8694 ( .C (clk), .D (signal_11239), .Q (signal_11240) ) ;
    buf_clk cell_8710 ( .C (clk), .D (signal_11255), .Q (signal_11256) ) ;
    buf_clk cell_8726 ( .C (clk), .D (signal_11271), .Q (signal_11272) ) ;
    buf_clk cell_8742 ( .C (clk), .D (signal_11287), .Q (signal_11288) ) ;
    buf_clk cell_8758 ( .C (clk), .D (signal_11303), .Q (signal_11304) ) ;
    buf_clk cell_8774 ( .C (clk), .D (signal_11319), .Q (signal_11320) ) ;
    buf_clk cell_8790 ( .C (clk), .D (signal_11335), .Q (signal_11336) ) ;
    buf_clk cell_8806 ( .C (clk), .D (signal_11351), .Q (signal_11352) ) ;
    buf_clk cell_8822 ( .C (clk), .D (signal_11367), .Q (signal_11368) ) ;
    buf_clk cell_8838 ( .C (clk), .D (signal_11383), .Q (signal_11384) ) ;
    buf_clk cell_8854 ( .C (clk), .D (signal_11399), .Q (signal_11400) ) ;
    buf_clk cell_8870 ( .C (clk), .D (signal_11415), .Q (signal_11416) ) ;
    buf_clk cell_8886 ( .C (clk), .D (signal_11431), .Q (signal_11432) ) ;
    buf_clk cell_8902 ( .C (clk), .D (signal_11447), .Q (signal_11448) ) ;
    buf_clk cell_8918 ( .C (clk), .D (signal_11463), .Q (signal_11464) ) ;
    buf_clk cell_8934 ( .C (clk), .D (signal_11479), .Q (signal_11480) ) ;
    buf_clk cell_8950 ( .C (clk), .D (signal_11495), .Q (signal_11496) ) ;
    buf_clk cell_8966 ( .C (clk), .D (signal_11511), .Q (signal_11512) ) ;
    buf_clk cell_8982 ( .C (clk), .D (signal_11527), .Q (signal_11528) ) ;
    buf_clk cell_8998 ( .C (clk), .D (signal_11543), .Q (signal_11544) ) ;
    buf_clk cell_9014 ( .C (clk), .D (signal_11559), .Q (signal_11560) ) ;
    buf_clk cell_9030 ( .C (clk), .D (signal_11575), .Q (signal_11576) ) ;
    buf_clk cell_9046 ( .C (clk), .D (signal_11591), .Q (signal_11592) ) ;
    buf_clk cell_9062 ( .C (clk), .D (signal_11607), .Q (signal_11608) ) ;
    buf_clk cell_9078 ( .C (clk), .D (signal_11623), .Q (signal_11624) ) ;
    buf_clk cell_9094 ( .C (clk), .D (signal_11639), .Q (signal_11640) ) ;
    buf_clk cell_9110 ( .C (clk), .D (signal_11655), .Q (signal_11656) ) ;
    buf_clk cell_9126 ( .C (clk), .D (signal_11671), .Q (signal_11672) ) ;
    buf_clk cell_9142 ( .C (clk), .D (signal_11687), .Q (signal_11688) ) ;
    buf_clk cell_9158 ( .C (clk), .D (signal_11703), .Q (signal_11704) ) ;
    buf_clk cell_9174 ( .C (clk), .D (signal_11719), .Q (signal_11720) ) ;
    buf_clk cell_9190 ( .C (clk), .D (signal_11735), .Q (signal_11736) ) ;
    buf_clk cell_9206 ( .C (clk), .D (signal_11751), .Q (signal_11752) ) ;
    buf_clk cell_9222 ( .C (clk), .D (signal_11767), .Q (signal_11768) ) ;
    buf_clk cell_9238 ( .C (clk), .D (signal_11783), .Q (signal_11784) ) ;
    buf_clk cell_9254 ( .C (clk), .D (signal_11799), .Q (signal_11800) ) ;
    buf_clk cell_9270 ( .C (clk), .D (signal_11815), .Q (signal_11816) ) ;
    buf_clk cell_9286 ( .C (clk), .D (signal_11831), .Q (signal_11832) ) ;
    buf_clk cell_9302 ( .C (clk), .D (signal_11847), .Q (signal_11848) ) ;
    buf_clk cell_9318 ( .C (clk), .D (signal_11863), .Q (signal_11864) ) ;
    buf_clk cell_9334 ( .C (clk), .D (signal_11879), .Q (signal_11880) ) ;
    buf_clk cell_9350 ( .C (clk), .D (signal_11895), .Q (signal_11896) ) ;
    buf_clk cell_9366 ( .C (clk), .D (signal_11911), .Q (signal_11912) ) ;
    buf_clk cell_9382 ( .C (clk), .D (signal_11927), .Q (signal_11928) ) ;
    buf_clk cell_9398 ( .C (clk), .D (signal_11943), .Q (signal_11944) ) ;
    buf_clk cell_9414 ( .C (clk), .D (signal_11959), .Q (signal_11960) ) ;
    buf_clk cell_9430 ( .C (clk), .D (signal_11975), .Q (signal_11976) ) ;
    buf_clk cell_9446 ( .C (clk), .D (signal_11991), .Q (signal_11992) ) ;
    buf_clk cell_9462 ( .C (clk), .D (signal_12007), .Q (signal_12008) ) ;
    buf_clk cell_9478 ( .C (clk), .D (signal_12023), .Q (signal_12024) ) ;
    buf_clk cell_9494 ( .C (clk), .D (signal_12039), .Q (signal_12040) ) ;
    buf_clk cell_9510 ( .C (clk), .D (signal_12055), .Q (signal_12056) ) ;
    buf_clk cell_9526 ( .C (clk), .D (signal_12071), .Q (signal_12072) ) ;
    buf_clk cell_9542 ( .C (clk), .D (signal_12087), .Q (signal_12088) ) ;
    buf_clk cell_9558 ( .C (clk), .D (signal_12103), .Q (signal_12104) ) ;
    buf_clk cell_9574 ( .C (clk), .D (signal_12119), .Q (signal_12120) ) ;
    buf_clk cell_9590 ( .C (clk), .D (signal_12135), .Q (signal_12136) ) ;
    buf_clk cell_9606 ( .C (clk), .D (signal_12151), .Q (signal_12152) ) ;
    buf_clk cell_9622 ( .C (clk), .D (signal_12167), .Q (signal_12168) ) ;
    buf_clk cell_9638 ( .C (clk), .D (signal_12183), .Q (signal_12184) ) ;
    buf_clk cell_9654 ( .C (clk), .D (signal_12199), .Q (signal_12200) ) ;
    buf_clk cell_9670 ( .C (clk), .D (signal_12215), .Q (signal_12216) ) ;
    buf_clk cell_9686 ( .C (clk), .D (signal_12231), .Q (signal_12232) ) ;
    buf_clk cell_9702 ( .C (clk), .D (signal_12247), .Q (signal_12248) ) ;
    buf_clk cell_9718 ( .C (clk), .D (signal_12263), .Q (signal_12264) ) ;
    buf_clk cell_9734 ( .C (clk), .D (signal_12279), .Q (signal_12280) ) ;
    buf_clk cell_9750 ( .C (clk), .D (signal_12295), .Q (signal_12296) ) ;
    buf_clk cell_9766 ( .C (clk), .D (signal_12311), .Q (signal_12312) ) ;
    buf_clk cell_9782 ( .C (clk), .D (signal_12327), .Q (signal_12328) ) ;
    buf_clk cell_9798 ( .C (clk), .D (signal_12343), .Q (signal_12344) ) ;
    buf_clk cell_9814 ( .C (clk), .D (signal_12359), .Q (signal_12360) ) ;
    buf_clk cell_9830 ( .C (clk), .D (signal_12375), .Q (signal_12376) ) ;
    buf_clk cell_9846 ( .C (clk), .D (signal_12391), .Q (signal_12392) ) ;
    buf_clk cell_9862 ( .C (clk), .D (signal_12407), .Q (signal_12408) ) ;
    buf_clk cell_9878 ( .C (clk), .D (signal_12423), .Q (signal_12424) ) ;
    buf_clk cell_9894 ( .C (clk), .D (signal_12439), .Q (signal_12440) ) ;
    buf_clk cell_9910 ( .C (clk), .D (signal_12455), .Q (signal_12456) ) ;
    buf_clk cell_9926 ( .C (clk), .D (signal_12471), .Q (signal_12472) ) ;
    buf_clk cell_9942 ( .C (clk), .D (signal_12487), .Q (signal_12488) ) ;
    buf_clk cell_9958 ( .C (clk), .D (signal_12503), .Q (signal_12504) ) ;
    buf_clk cell_9974 ( .C (clk), .D (signal_12519), .Q (signal_12520) ) ;
    buf_clk cell_9990 ( .C (clk), .D (signal_12535), .Q (signal_12536) ) ;
    buf_clk cell_10006 ( .C (clk), .D (signal_12551), .Q (signal_12552) ) ;
    buf_clk cell_10022 ( .C (clk), .D (signal_12567), .Q (signal_12568) ) ;
    buf_clk cell_10038 ( .C (clk), .D (signal_12583), .Q (signal_12584) ) ;
    buf_clk cell_10054 ( .C (clk), .D (signal_12599), .Q (signal_12600) ) ;
    buf_clk cell_10070 ( .C (clk), .D (signal_12615), .Q (signal_12616) ) ;
    buf_clk cell_10086 ( .C (clk), .D (signal_12631), .Q (signal_12632) ) ;
    buf_clk cell_10102 ( .C (clk), .D (signal_12647), .Q (signal_12648) ) ;
    buf_clk cell_10118 ( .C (clk), .D (signal_12663), .Q (signal_12664) ) ;
    buf_clk cell_10134 ( .C (clk), .D (signal_12679), .Q (signal_12680) ) ;
    buf_clk cell_10150 ( .C (clk), .D (signal_12695), .Q (signal_12696) ) ;
    buf_clk cell_10166 ( .C (clk), .D (signal_12711), .Q (signal_12712) ) ;
    buf_clk cell_10182 ( .C (clk), .D (signal_12727), .Q (signal_12728) ) ;
    buf_clk cell_10198 ( .C (clk), .D (signal_12743), .Q (signal_12744) ) ;
    buf_clk cell_10214 ( .C (clk), .D (signal_12759), .Q (signal_12760) ) ;
    buf_clk cell_10230 ( .C (clk), .D (signal_12775), .Q (signal_12776) ) ;
    buf_clk cell_10246 ( .C (clk), .D (signal_12791), .Q (signal_12792) ) ;
    buf_clk cell_10262 ( .C (clk), .D (signal_12807), .Q (signal_12808) ) ;
    buf_clk cell_10278 ( .C (clk), .D (signal_12823), .Q (signal_12824) ) ;
    buf_clk cell_10294 ( .C (clk), .D (signal_12839), .Q (signal_12840) ) ;
    buf_clk cell_10310 ( .C (clk), .D (signal_12855), .Q (signal_12856) ) ;
    buf_clk cell_10326 ( .C (clk), .D (signal_12871), .Q (signal_12872) ) ;
    buf_clk cell_10342 ( .C (clk), .D (signal_12887), .Q (signal_12888) ) ;
    buf_clk cell_10358 ( .C (clk), .D (signal_12903), .Q (signal_12904) ) ;
    buf_clk cell_10374 ( .C (clk), .D (signal_12919), .Q (signal_12920) ) ;
    buf_clk cell_10390 ( .C (clk), .D (signal_12935), .Q (signal_12936) ) ;
    buf_clk cell_10406 ( .C (clk), .D (signal_12951), .Q (signal_12952) ) ;
    buf_clk cell_10422 ( .C (clk), .D (signal_12967), .Q (signal_12968) ) ;
    buf_clk cell_10438 ( .C (clk), .D (signal_12983), .Q (signal_12984) ) ;
    buf_clk cell_10454 ( .C (clk), .D (signal_12999), .Q (signal_13000) ) ;
    buf_clk cell_10470 ( .C (clk), .D (signal_13015), .Q (signal_13016) ) ;
    buf_clk cell_10486 ( .C (clk), .D (signal_13031), .Q (signal_13032) ) ;
    buf_clk cell_10502 ( .C (clk), .D (signal_13047), .Q (signal_13048) ) ;
    buf_clk cell_10518 ( .C (clk), .D (signal_13063), .Q (signal_13064) ) ;
    buf_clk cell_10534 ( .C (clk), .D (signal_13079), .Q (signal_13080) ) ;
    buf_clk cell_10550 ( .C (clk), .D (signal_13095), .Q (signal_13096) ) ;
    buf_clk cell_10566 ( .C (clk), .D (signal_13111), .Q (signal_13112) ) ;
    buf_clk cell_10582 ( .C (clk), .D (signal_13127), .Q (signal_13128) ) ;
    buf_clk cell_10598 ( .C (clk), .D (signal_13143), .Q (signal_13144) ) ;
    buf_clk cell_10614 ( .C (clk), .D (signal_13159), .Q (signal_13160) ) ;
    buf_clk cell_10630 ( .C (clk), .D (signal_13175), .Q (signal_13176) ) ;
    buf_clk cell_10646 ( .C (clk), .D (signal_13191), .Q (signal_13192) ) ;
    buf_clk cell_10662 ( .C (clk), .D (signal_13207), .Q (signal_13208) ) ;
    buf_clk cell_10678 ( .C (clk), .D (signal_13223), .Q (signal_13224) ) ;
    buf_clk cell_10694 ( .C (clk), .D (signal_13239), .Q (signal_13240) ) ;
    buf_clk cell_10710 ( .C (clk), .D (signal_13255), .Q (signal_13256) ) ;
    buf_clk cell_10726 ( .C (clk), .D (signal_13271), .Q (signal_13272) ) ;
    buf_clk cell_10742 ( .C (clk), .D (signal_13287), .Q (signal_13288) ) ;
    buf_clk cell_10758 ( .C (clk), .D (signal_13303), .Q (signal_13304) ) ;
    buf_clk cell_10774 ( .C (clk), .D (signal_13319), .Q (signal_13320) ) ;
    buf_clk cell_10790 ( .C (clk), .D (signal_13335), .Q (signal_13336) ) ;
    buf_clk cell_10806 ( .C (clk), .D (signal_13351), .Q (signal_13352) ) ;
    buf_clk cell_10822 ( .C (clk), .D (signal_13367), .Q (signal_13368) ) ;
    buf_clk cell_10838 ( .C (clk), .D (signal_13383), .Q (signal_13384) ) ;
    buf_clk cell_10854 ( .C (clk), .D (signal_13399), .Q (signal_13400) ) ;
    buf_clk cell_10870 ( .C (clk), .D (signal_13415), .Q (signal_13416) ) ;
    buf_clk cell_10886 ( .C (clk), .D (signal_13431), .Q (signal_13432) ) ;
    buf_clk cell_10902 ( .C (clk), .D (signal_13447), .Q (signal_13448) ) ;
    buf_clk cell_10918 ( .C (clk), .D (signal_13463), .Q (signal_13464) ) ;
    buf_clk cell_10934 ( .C (clk), .D (signal_13479), .Q (signal_13480) ) ;
    buf_clk cell_10950 ( .C (clk), .D (signal_13495), .Q (signal_13496) ) ;
    buf_clk cell_10966 ( .C (clk), .D (signal_13511), .Q (signal_13512) ) ;
    buf_clk cell_10982 ( .C (clk), .D (signal_13527), .Q (signal_13528) ) ;
    buf_clk cell_10998 ( .C (clk), .D (signal_13543), .Q (signal_13544) ) ;
    buf_clk cell_11014 ( .C (clk), .D (signal_13559), .Q (signal_13560) ) ;
    buf_clk cell_11030 ( .C (clk), .D (signal_13575), .Q (signal_13576) ) ;
    buf_clk cell_11046 ( .C (clk), .D (signal_13591), .Q (signal_13592) ) ;
    buf_clk cell_11062 ( .C (clk), .D (signal_13607), .Q (signal_13608) ) ;
    buf_clk cell_11078 ( .C (clk), .D (signal_13623), .Q (signal_13624) ) ;
    buf_clk cell_11094 ( .C (clk), .D (signal_13639), .Q (signal_13640) ) ;
    buf_clk cell_11110 ( .C (clk), .D (signal_13655), .Q (signal_13656) ) ;
    buf_clk cell_11126 ( .C (clk), .D (signal_13671), .Q (signal_13672) ) ;
    buf_clk cell_11142 ( .C (clk), .D (signal_13687), .Q (signal_13688) ) ;
    buf_clk cell_11158 ( .C (clk), .D (signal_13703), .Q (signal_13704) ) ;
    buf_clk cell_11174 ( .C (clk), .D (signal_13719), .Q (signal_13720) ) ;
    buf_clk cell_11190 ( .C (clk), .D (signal_13735), .Q (signal_13736) ) ;
    buf_clk cell_11206 ( .C (clk), .D (signal_13751), .Q (signal_13752) ) ;
    buf_clk cell_11222 ( .C (clk), .D (signal_13767), .Q (signal_13768) ) ;
    buf_clk cell_11238 ( .C (clk), .D (signal_13783), .Q (signal_13784) ) ;
    buf_clk cell_11254 ( .C (clk), .D (signal_13799), .Q (signal_13800) ) ;
    buf_clk cell_11270 ( .C (clk), .D (signal_13815), .Q (signal_13816) ) ;
    buf_clk cell_11286 ( .C (clk), .D (signal_13831), .Q (signal_13832) ) ;
    buf_clk cell_11302 ( .C (clk), .D (signal_13847), .Q (signal_13848) ) ;
    buf_clk cell_11318 ( .C (clk), .D (signal_13863), .Q (signal_13864) ) ;
    buf_clk cell_11334 ( .C (clk), .D (signal_13879), .Q (signal_13880) ) ;
    buf_clk cell_11350 ( .C (clk), .D (signal_13895), .Q (signal_13896) ) ;
    buf_clk cell_11366 ( .C (clk), .D (signal_13911), .Q (signal_13912) ) ;
    buf_clk cell_11382 ( .C (clk), .D (signal_13927), .Q (signal_13928) ) ;
    buf_clk cell_11398 ( .C (clk), .D (signal_13943), .Q (signal_13944) ) ;
    buf_clk cell_11414 ( .C (clk), .D (signal_13959), .Q (signal_13960) ) ;
    buf_clk cell_11430 ( .C (clk), .D (signal_13975), .Q (signal_13976) ) ;
    buf_clk cell_11446 ( .C (clk), .D (signal_13991), .Q (signal_13992) ) ;
    buf_clk cell_11462 ( .C (clk), .D (signal_14007), .Q (signal_14008) ) ;
    buf_clk cell_11478 ( .C (clk), .D (signal_14023), .Q (signal_14024) ) ;
    buf_clk cell_11494 ( .C (clk), .D (signal_14039), .Q (signal_14040) ) ;
    buf_clk cell_11510 ( .C (clk), .D (signal_14055), .Q (signal_14056) ) ;
    buf_clk cell_11526 ( .C (clk), .D (signal_14071), .Q (signal_14072) ) ;
    buf_clk cell_11542 ( .C (clk), .D (signal_14087), .Q (signal_14088) ) ;
    buf_clk cell_11558 ( .C (clk), .D (signal_14103), .Q (signal_14104) ) ;
    buf_clk cell_11574 ( .C (clk), .D (signal_14119), .Q (signal_14120) ) ;
    buf_clk cell_11590 ( .C (clk), .D (signal_14135), .Q (signal_14136) ) ;
    buf_clk cell_11606 ( .C (clk), .D (signal_14151), .Q (signal_14152) ) ;
    buf_clk cell_11622 ( .C (clk), .D (signal_14167), .Q (signal_14168) ) ;
    buf_clk cell_11638 ( .C (clk), .D (signal_14183), .Q (signal_14184) ) ;
    buf_clk cell_11654 ( .C (clk), .D (signal_14199), .Q (signal_14200) ) ;
    buf_clk cell_11670 ( .C (clk), .D (signal_14215), .Q (signal_14216) ) ;
    buf_clk cell_11686 ( .C (clk), .D (signal_14231), .Q (signal_14232) ) ;
    buf_clk cell_11702 ( .C (clk), .D (signal_14247), .Q (signal_14248) ) ;
    buf_clk cell_11718 ( .C (clk), .D (signal_14263), .Q (signal_14264) ) ;
    buf_clk cell_11734 ( .C (clk), .D (signal_14279), .Q (signal_14280) ) ;
    buf_clk cell_11750 ( .C (clk), .D (signal_14295), .Q (signal_14296) ) ;
    buf_clk cell_11766 ( .C (clk), .D (signal_14311), .Q (signal_14312) ) ;
    buf_clk cell_11782 ( .C (clk), .D (signal_14327), .Q (signal_14328) ) ;
    buf_clk cell_11798 ( .C (clk), .D (signal_14343), .Q (signal_14344) ) ;
    buf_clk cell_11814 ( .C (clk), .D (signal_14359), .Q (signal_14360) ) ;
    buf_clk cell_11830 ( .C (clk), .D (signal_14375), .Q (signal_14376) ) ;
    buf_clk cell_11846 ( .C (clk), .D (signal_14391), .Q (signal_14392) ) ;
    buf_clk cell_11862 ( .C (clk), .D (signal_14407), .Q (signal_14408) ) ;
    buf_clk cell_11878 ( .C (clk), .D (signal_14423), .Q (signal_14424) ) ;
    buf_clk cell_11894 ( .C (clk), .D (signal_14439), .Q (signal_14440) ) ;
    buf_clk cell_11910 ( .C (clk), .D (signal_14455), .Q (signal_14456) ) ;
    buf_clk cell_11926 ( .C (clk), .D (signal_14471), .Q (signal_14472) ) ;
    buf_clk cell_11942 ( .C (clk), .D (signal_14487), .Q (signal_14488) ) ;
    buf_clk cell_11958 ( .C (clk), .D (signal_14503), .Q (signal_14504) ) ;
    buf_clk cell_11974 ( .C (clk), .D (signal_14519), .Q (signal_14520) ) ;
    buf_clk cell_11990 ( .C (clk), .D (signal_14535), .Q (signal_14536) ) ;
    buf_clk cell_12006 ( .C (clk), .D (signal_14551), .Q (signal_14552) ) ;
    buf_clk cell_12022 ( .C (clk), .D (signal_14567), .Q (signal_14568) ) ;
    buf_clk cell_12038 ( .C (clk), .D (signal_14583), .Q (signal_14584) ) ;
    buf_clk cell_12054 ( .C (clk), .D (signal_14599), .Q (signal_14600) ) ;
    buf_clk cell_12070 ( .C (clk), .D (signal_14615), .Q (signal_14616) ) ;
    buf_clk cell_12086 ( .C (clk), .D (signal_14631), .Q (signal_14632) ) ;
    buf_clk cell_12102 ( .C (clk), .D (signal_14647), .Q (signal_14648) ) ;
    buf_clk cell_12118 ( .C (clk), .D (signal_14663), .Q (signal_14664) ) ;
    buf_clk cell_12134 ( .C (clk), .D (signal_14679), .Q (signal_14680) ) ;
    buf_clk cell_12150 ( .C (clk), .D (signal_14695), .Q (signal_14696) ) ;
    buf_clk cell_12166 ( .C (clk), .D (signal_14711), .Q (signal_14712) ) ;
    buf_clk cell_12182 ( .C (clk), .D (signal_14727), .Q (signal_14728) ) ;
    buf_clk cell_12198 ( .C (clk), .D (signal_14743), .Q (signal_14744) ) ;
    buf_clk cell_12214 ( .C (clk), .D (signal_14759), .Q (signal_14760) ) ;
    buf_clk cell_12230 ( .C (clk), .D (signal_14775), .Q (signal_14776) ) ;
    buf_clk cell_12246 ( .C (clk), .D (signal_14791), .Q (signal_14792) ) ;
    buf_clk cell_12262 ( .C (clk), .D (signal_14807), .Q (signal_14808) ) ;
    buf_clk cell_12278 ( .C (clk), .D (signal_14823), .Q (signal_14824) ) ;
    buf_clk cell_12294 ( .C (clk), .D (signal_14839), .Q (signal_14840) ) ;
    buf_clk cell_12310 ( .C (clk), .D (signal_14855), .Q (signal_14856) ) ;
    buf_clk cell_12326 ( .C (clk), .D (signal_14871), .Q (signal_14872) ) ;
    buf_clk cell_12342 ( .C (clk), .D (signal_14887), .Q (signal_14888) ) ;
    buf_clk cell_12358 ( .C (clk), .D (signal_14903), .Q (signal_14904) ) ;
    buf_clk cell_12374 ( .C (clk), .D (signal_14919), .Q (signal_14920) ) ;
    buf_clk cell_12390 ( .C (clk), .D (signal_14935), .Q (signal_14936) ) ;

    /* cells in depth 11 */
    buf_clk cell_2371 ( .C (clk), .D (signal_4916), .Q (signal_4917) ) ;
    buf_clk cell_2383 ( .C (clk), .D (signal_4928), .Q (signal_4929) ) ;
    buf_clk cell_2395 ( .C (clk), .D (signal_4940), .Q (signal_4941) ) ;
    buf_clk cell_2411 ( .C (clk), .D (signal_4956), .Q (signal_4957) ) ;
    buf_clk cell_2427 ( .C (clk), .D (signal_4972), .Q (signal_4973) ) ;
    buf_clk cell_2443 ( .C (clk), .D (signal_4988), .Q (signal_4989) ) ;
    buf_clk cell_2459 ( .C (clk), .D (signal_5004), .Q (signal_5005) ) ;
    buf_clk cell_2475 ( .C (clk), .D (signal_5020), .Q (signal_5021) ) ;
    buf_clk cell_2491 ( .C (clk), .D (signal_5036), .Q (signal_5037) ) ;
    buf_clk cell_2507 ( .C (clk), .D (signal_5052), .Q (signal_5053) ) ;
    buf_clk cell_2523 ( .C (clk), .D (signal_5068), .Q (signal_5069) ) ;
    buf_clk cell_2539 ( .C (clk), .D (signal_5084), .Q (signal_5085) ) ;
    buf_clk cell_2555 ( .C (clk), .D (signal_5100), .Q (signal_5101) ) ;
    buf_clk cell_2571 ( .C (clk), .D (signal_5116), .Q (signal_5117) ) ;
    buf_clk cell_2587 ( .C (clk), .D (signal_5132), .Q (signal_5133) ) ;
    buf_clk cell_2603 ( .C (clk), .D (signal_5148), .Q (signal_5149) ) ;
    buf_clk cell_2619 ( .C (clk), .D (signal_5164), .Q (signal_5165) ) ;
    buf_clk cell_2635 ( .C (clk), .D (signal_5180), .Q (signal_5181) ) ;
    buf_clk cell_2651 ( .C (clk), .D (signal_5196), .Q (signal_5197) ) ;
    buf_clk cell_2667 ( .C (clk), .D (signal_5212), .Q (signal_5213) ) ;
    buf_clk cell_2683 ( .C (clk), .D (signal_5228), .Q (signal_5229) ) ;
    buf_clk cell_2699 ( .C (clk), .D (signal_5244), .Q (signal_5245) ) ;
    buf_clk cell_2715 ( .C (clk), .D (signal_5260), .Q (signal_5261) ) ;
    buf_clk cell_2731 ( .C (clk), .D (signal_5276), .Q (signal_5277) ) ;
    buf_clk cell_2747 ( .C (clk), .D (signal_5292), .Q (signal_5293) ) ;
    buf_clk cell_2763 ( .C (clk), .D (signal_5308), .Q (signal_5309) ) ;
    buf_clk cell_2779 ( .C (clk), .D (signal_5324), .Q (signal_5325) ) ;
    buf_clk cell_2795 ( .C (clk), .D (signal_5340), .Q (signal_5341) ) ;
    buf_clk cell_2811 ( .C (clk), .D (signal_5356), .Q (signal_5357) ) ;
    buf_clk cell_2827 ( .C (clk), .D (signal_5372), .Q (signal_5373) ) ;
    buf_clk cell_2843 ( .C (clk), .D (signal_5388), .Q (signal_5389) ) ;
    buf_clk cell_2859 ( .C (clk), .D (signal_5404), .Q (signal_5405) ) ;
    buf_clk cell_2875 ( .C (clk), .D (signal_5420), .Q (signal_5421) ) ;
    buf_clk cell_2891 ( .C (clk), .D (signal_5436), .Q (signal_5437) ) ;
    buf_clk cell_2907 ( .C (clk), .D (signal_5452), .Q (signal_5453) ) ;
    buf_clk cell_2923 ( .C (clk), .D (signal_5468), .Q (signal_5469) ) ;
    buf_clk cell_2939 ( .C (clk), .D (signal_5484), .Q (signal_5485) ) ;
    buf_clk cell_2955 ( .C (clk), .D (signal_5500), .Q (signal_5501) ) ;
    buf_clk cell_2971 ( .C (clk), .D (signal_5516), .Q (signal_5517) ) ;
    buf_clk cell_2987 ( .C (clk), .D (signal_5532), .Q (signal_5533) ) ;
    buf_clk cell_3003 ( .C (clk), .D (signal_5548), .Q (signal_5549) ) ;
    buf_clk cell_3019 ( .C (clk), .D (signal_5564), .Q (signal_5565) ) ;
    buf_clk cell_3035 ( .C (clk), .D (signal_5580), .Q (signal_5581) ) ;
    buf_clk cell_3051 ( .C (clk), .D (signal_5596), .Q (signal_5597) ) ;
    buf_clk cell_3067 ( .C (clk), .D (signal_5612), .Q (signal_5613) ) ;
    buf_clk cell_3083 ( .C (clk), .D (signal_5628), .Q (signal_5629) ) ;
    buf_clk cell_3099 ( .C (clk), .D (signal_5644), .Q (signal_5645) ) ;
    buf_clk cell_3115 ( .C (clk), .D (signal_5660), .Q (signal_5661) ) ;
    buf_clk cell_3131 ( .C (clk), .D (signal_5676), .Q (signal_5677) ) ;
    buf_clk cell_3147 ( .C (clk), .D (signal_5692), .Q (signal_5693) ) ;
    buf_clk cell_3163 ( .C (clk), .D (signal_5708), .Q (signal_5709) ) ;
    buf_clk cell_3179 ( .C (clk), .D (signal_5724), .Q (signal_5725) ) ;
    buf_clk cell_3195 ( .C (clk), .D (signal_5740), .Q (signal_5741) ) ;
    buf_clk cell_3211 ( .C (clk), .D (signal_5756), .Q (signal_5757) ) ;
    buf_clk cell_3227 ( .C (clk), .D (signal_5772), .Q (signal_5773) ) ;
    buf_clk cell_3243 ( .C (clk), .D (signal_5788), .Q (signal_5789) ) ;
    buf_clk cell_3259 ( .C (clk), .D (signal_5804), .Q (signal_5805) ) ;
    buf_clk cell_3275 ( .C (clk), .D (signal_5820), .Q (signal_5821) ) ;
    buf_clk cell_3291 ( .C (clk), .D (signal_5836), .Q (signal_5837) ) ;
    buf_clk cell_3307 ( .C (clk), .D (signal_5852), .Q (signal_5853) ) ;
    buf_clk cell_3323 ( .C (clk), .D (signal_5868), .Q (signal_5869) ) ;
    buf_clk cell_3339 ( .C (clk), .D (signal_5884), .Q (signal_5885) ) ;
    buf_clk cell_3355 ( .C (clk), .D (signal_5900), .Q (signal_5901) ) ;
    buf_clk cell_3371 ( .C (clk), .D (signal_5916), .Q (signal_5917) ) ;
    buf_clk cell_3387 ( .C (clk), .D (signal_5932), .Q (signal_5933) ) ;
    buf_clk cell_3403 ( .C (clk), .D (signal_5948), .Q (signal_5949) ) ;
    buf_clk cell_3419 ( .C (clk), .D (signal_5964), .Q (signal_5965) ) ;
    buf_clk cell_3435 ( .C (clk), .D (signal_5980), .Q (signal_5981) ) ;
    buf_clk cell_3451 ( .C (clk), .D (signal_5996), .Q (signal_5997) ) ;
    buf_clk cell_3467 ( .C (clk), .D (signal_6012), .Q (signal_6013) ) ;
    buf_clk cell_3483 ( .C (clk), .D (signal_6028), .Q (signal_6029) ) ;
    buf_clk cell_3499 ( .C (clk), .D (signal_6044), .Q (signal_6045) ) ;
    buf_clk cell_3515 ( .C (clk), .D (signal_6060), .Q (signal_6061) ) ;
    buf_clk cell_3531 ( .C (clk), .D (signal_6076), .Q (signal_6077) ) ;
    buf_clk cell_3547 ( .C (clk), .D (signal_6092), .Q (signal_6093) ) ;
    buf_clk cell_3563 ( .C (clk), .D (signal_6108), .Q (signal_6109) ) ;
    buf_clk cell_3579 ( .C (clk), .D (signal_6124), .Q (signal_6125) ) ;
    buf_clk cell_3595 ( .C (clk), .D (signal_6140), .Q (signal_6141) ) ;
    buf_clk cell_3611 ( .C (clk), .D (signal_6156), .Q (signal_6157) ) ;
    buf_clk cell_3627 ( .C (clk), .D (signal_6172), .Q (signal_6173) ) ;
    buf_clk cell_3643 ( .C (clk), .D (signal_6188), .Q (signal_6189) ) ;
    buf_clk cell_3659 ( .C (clk), .D (signal_6204), .Q (signal_6205) ) ;
    buf_clk cell_3675 ( .C (clk), .D (signal_6220), .Q (signal_6221) ) ;
    buf_clk cell_3691 ( .C (clk), .D (signal_6236), .Q (signal_6237) ) ;
    buf_clk cell_3707 ( .C (clk), .D (signal_6252), .Q (signal_6253) ) ;
    buf_clk cell_3723 ( .C (clk), .D (signal_6268), .Q (signal_6269) ) ;
    buf_clk cell_3739 ( .C (clk), .D (signal_6284), .Q (signal_6285) ) ;
    buf_clk cell_3755 ( .C (clk), .D (signal_6300), .Q (signal_6301) ) ;
    buf_clk cell_3771 ( .C (clk), .D (signal_6316), .Q (signal_6317) ) ;
    buf_clk cell_3787 ( .C (clk), .D (signal_6332), .Q (signal_6333) ) ;
    buf_clk cell_3803 ( .C (clk), .D (signal_6348), .Q (signal_6349) ) ;
    buf_clk cell_3819 ( .C (clk), .D (signal_6364), .Q (signal_6365) ) ;
    buf_clk cell_3835 ( .C (clk), .D (signal_6380), .Q (signal_6381) ) ;
    buf_clk cell_3851 ( .C (clk), .D (signal_6396), .Q (signal_6397) ) ;
    buf_clk cell_3867 ( .C (clk), .D (signal_6412), .Q (signal_6413) ) ;
    buf_clk cell_3883 ( .C (clk), .D (signal_6428), .Q (signal_6429) ) ;
    buf_clk cell_3899 ( .C (clk), .D (signal_6444), .Q (signal_6445) ) ;
    buf_clk cell_3915 ( .C (clk), .D (signal_6460), .Q (signal_6461) ) ;
    buf_clk cell_3931 ( .C (clk), .D (signal_6476), .Q (signal_6477) ) ;
    buf_clk cell_3947 ( .C (clk), .D (signal_6492), .Q (signal_6493) ) ;
    buf_clk cell_3963 ( .C (clk), .D (signal_6508), .Q (signal_6509) ) ;
    buf_clk cell_3979 ( .C (clk), .D (signal_6524), .Q (signal_6525) ) ;
    buf_clk cell_3995 ( .C (clk), .D (signal_6540), .Q (signal_6541) ) ;
    buf_clk cell_4011 ( .C (clk), .D (signal_6556), .Q (signal_6557) ) ;
    buf_clk cell_4027 ( .C (clk), .D (signal_6572), .Q (signal_6573) ) ;
    buf_clk cell_4043 ( .C (clk), .D (signal_6588), .Q (signal_6589) ) ;
    buf_clk cell_4059 ( .C (clk), .D (signal_6604), .Q (signal_6605) ) ;
    buf_clk cell_4075 ( .C (clk), .D (signal_6620), .Q (signal_6621) ) ;
    buf_clk cell_4091 ( .C (clk), .D (signal_6636), .Q (signal_6637) ) ;
    buf_clk cell_4107 ( .C (clk), .D (signal_6652), .Q (signal_6653) ) ;
    buf_clk cell_4123 ( .C (clk), .D (signal_6668), .Q (signal_6669) ) ;
    buf_clk cell_4139 ( .C (clk), .D (signal_6684), .Q (signal_6685) ) ;
    buf_clk cell_4155 ( .C (clk), .D (signal_6700), .Q (signal_6701) ) ;
    buf_clk cell_4171 ( .C (clk), .D (signal_6716), .Q (signal_6717) ) ;
    buf_clk cell_4187 ( .C (clk), .D (signal_6732), .Q (signal_6733) ) ;
    buf_clk cell_4203 ( .C (clk), .D (signal_6748), .Q (signal_6749) ) ;
    buf_clk cell_4219 ( .C (clk), .D (signal_6764), .Q (signal_6765) ) ;
    buf_clk cell_4235 ( .C (clk), .D (signal_6780), .Q (signal_6781) ) ;
    buf_clk cell_4251 ( .C (clk), .D (signal_6796), .Q (signal_6797) ) ;
    buf_clk cell_4267 ( .C (clk), .D (signal_6812), .Q (signal_6813) ) ;
    buf_clk cell_4283 ( .C (clk), .D (signal_6828), .Q (signal_6829) ) ;
    buf_clk cell_4299 ( .C (clk), .D (signal_6844), .Q (signal_6845) ) ;
    buf_clk cell_4315 ( .C (clk), .D (signal_6860), .Q (signal_6861) ) ;
    buf_clk cell_4331 ( .C (clk), .D (signal_6876), .Q (signal_6877) ) ;
    buf_clk cell_4347 ( .C (clk), .D (signal_6892), .Q (signal_6893) ) ;
    buf_clk cell_4363 ( .C (clk), .D (signal_6908), .Q (signal_6909) ) ;
    buf_clk cell_4379 ( .C (clk), .D (signal_6924), .Q (signal_6925) ) ;
    buf_clk cell_4395 ( .C (clk), .D (signal_6940), .Q (signal_6941) ) ;
    buf_clk cell_4411 ( .C (clk), .D (signal_6956), .Q (signal_6957) ) ;
    buf_clk cell_4425 ( .C (clk), .D (signal_6970), .Q (signal_6971) ) ;
    buf_clk cell_4439 ( .C (clk), .D (signal_6984), .Q (signal_6985) ) ;
    buf_clk cell_4455 ( .C (clk), .D (signal_7000), .Q (signal_7001) ) ;
    buf_clk cell_4471 ( .C (clk), .D (signal_7016), .Q (signal_7017) ) ;
    buf_clk cell_4487 ( .C (clk), .D (signal_7032), .Q (signal_7033) ) ;
    buf_clk cell_4503 ( .C (clk), .D (signal_7048), .Q (signal_7049) ) ;
    buf_clk cell_4519 ( .C (clk), .D (signal_7064), .Q (signal_7065) ) ;
    buf_clk cell_4535 ( .C (clk), .D (signal_7080), .Q (signal_7081) ) ;
    buf_clk cell_4551 ( .C (clk), .D (signal_7096), .Q (signal_7097) ) ;
    buf_clk cell_4567 ( .C (clk), .D (signal_7112), .Q (signal_7113) ) ;
    buf_clk cell_4583 ( .C (clk), .D (signal_7128), .Q (signal_7129) ) ;
    buf_clk cell_4599 ( .C (clk), .D (signal_7144), .Q (signal_7145) ) ;
    buf_clk cell_4615 ( .C (clk), .D (signal_7160), .Q (signal_7161) ) ;
    buf_clk cell_4631 ( .C (clk), .D (signal_7176), .Q (signal_7177) ) ;
    buf_clk cell_4647 ( .C (clk), .D (signal_7192), .Q (signal_7193) ) ;
    buf_clk cell_4663 ( .C (clk), .D (signal_7208), .Q (signal_7209) ) ;
    buf_clk cell_4679 ( .C (clk), .D (signal_7224), .Q (signal_7225) ) ;
    buf_clk cell_4695 ( .C (clk), .D (signal_7240), .Q (signal_7241) ) ;
    buf_clk cell_4711 ( .C (clk), .D (signal_7256), .Q (signal_7257) ) ;
    buf_clk cell_4727 ( .C (clk), .D (signal_7272), .Q (signal_7273) ) ;
    buf_clk cell_4743 ( .C (clk), .D (signal_7288), .Q (signal_7289) ) ;
    buf_clk cell_4759 ( .C (clk), .D (signal_7304), .Q (signal_7305) ) ;
    buf_clk cell_4775 ( .C (clk), .D (signal_7320), .Q (signal_7321) ) ;
    buf_clk cell_4791 ( .C (clk), .D (signal_7336), .Q (signal_7337) ) ;
    buf_clk cell_4807 ( .C (clk), .D (signal_7352), .Q (signal_7353) ) ;
    buf_clk cell_4823 ( .C (clk), .D (signal_7368), .Q (signal_7369) ) ;
    buf_clk cell_4839 ( .C (clk), .D (signal_7384), .Q (signal_7385) ) ;
    buf_clk cell_4855 ( .C (clk), .D (signal_7400), .Q (signal_7401) ) ;
    buf_clk cell_4871 ( .C (clk), .D (signal_7416), .Q (signal_7417) ) ;
    buf_clk cell_4887 ( .C (clk), .D (signal_7432), .Q (signal_7433) ) ;
    buf_clk cell_4903 ( .C (clk), .D (signal_7448), .Q (signal_7449) ) ;
    buf_clk cell_4919 ( .C (clk), .D (signal_7464), .Q (signal_7465) ) ;
    buf_clk cell_4935 ( .C (clk), .D (signal_7480), .Q (signal_7481) ) ;
    buf_clk cell_4951 ( .C (clk), .D (signal_7496), .Q (signal_7497) ) ;
    buf_clk cell_4967 ( .C (clk), .D (signal_7512), .Q (signal_7513) ) ;
    buf_clk cell_4983 ( .C (clk), .D (signal_7528), .Q (signal_7529) ) ;
    buf_clk cell_4999 ( .C (clk), .D (signal_7544), .Q (signal_7545) ) ;
    buf_clk cell_5015 ( .C (clk), .D (signal_7560), .Q (signal_7561) ) ;
    buf_clk cell_5031 ( .C (clk), .D (signal_7576), .Q (signal_7577) ) ;
    buf_clk cell_5047 ( .C (clk), .D (signal_7592), .Q (signal_7593) ) ;
    buf_clk cell_5063 ( .C (clk), .D (signal_7608), .Q (signal_7609) ) ;
    buf_clk cell_5079 ( .C (clk), .D (signal_7624), .Q (signal_7625) ) ;
    buf_clk cell_5095 ( .C (clk), .D (signal_7640), .Q (signal_7641) ) ;
    buf_clk cell_5111 ( .C (clk), .D (signal_7656), .Q (signal_7657) ) ;
    buf_clk cell_5127 ( .C (clk), .D (signal_7672), .Q (signal_7673) ) ;
    buf_clk cell_5143 ( .C (clk), .D (signal_7688), .Q (signal_7689) ) ;
    buf_clk cell_5159 ( .C (clk), .D (signal_7704), .Q (signal_7705) ) ;
    buf_clk cell_5175 ( .C (clk), .D (signal_7720), .Q (signal_7721) ) ;
    buf_clk cell_5191 ( .C (clk), .D (signal_7736), .Q (signal_7737) ) ;
    buf_clk cell_5207 ( .C (clk), .D (signal_7752), .Q (signal_7753) ) ;
    buf_clk cell_5223 ( .C (clk), .D (signal_7768), .Q (signal_7769) ) ;
    buf_clk cell_5239 ( .C (clk), .D (signal_7784), .Q (signal_7785) ) ;
    buf_clk cell_5255 ( .C (clk), .D (signal_7800), .Q (signal_7801) ) ;
    buf_clk cell_5271 ( .C (clk), .D (signal_7816), .Q (signal_7817) ) ;
    buf_clk cell_5287 ( .C (clk), .D (signal_7832), .Q (signal_7833) ) ;
    buf_clk cell_5303 ( .C (clk), .D (signal_7848), .Q (signal_7849) ) ;
    buf_clk cell_5319 ( .C (clk), .D (signal_7864), .Q (signal_7865) ) ;
    buf_clk cell_5335 ( .C (clk), .D (signal_7880), .Q (signal_7881) ) ;
    buf_clk cell_5351 ( .C (clk), .D (signal_7896), .Q (signal_7897) ) ;
    buf_clk cell_5367 ( .C (clk), .D (signal_7912), .Q (signal_7913) ) ;
    buf_clk cell_5383 ( .C (clk), .D (signal_7928), .Q (signal_7929) ) ;
    buf_clk cell_5399 ( .C (clk), .D (signal_7944), .Q (signal_7945) ) ;
    buf_clk cell_5415 ( .C (clk), .D (signal_7960), .Q (signal_7961) ) ;
    buf_clk cell_5431 ( .C (clk), .D (signal_7976), .Q (signal_7977) ) ;
    buf_clk cell_5447 ( .C (clk), .D (signal_7992), .Q (signal_7993) ) ;
    buf_clk cell_5463 ( .C (clk), .D (signal_8008), .Q (signal_8009) ) ;
    buf_clk cell_5479 ( .C (clk), .D (signal_8024), .Q (signal_8025) ) ;
    buf_clk cell_5495 ( .C (clk), .D (signal_8040), .Q (signal_8041) ) ;
    buf_clk cell_5511 ( .C (clk), .D (signal_8056), .Q (signal_8057) ) ;
    buf_clk cell_5527 ( .C (clk), .D (signal_8072), .Q (signal_8073) ) ;
    buf_clk cell_5543 ( .C (clk), .D (signal_8088), .Q (signal_8089) ) ;
    buf_clk cell_5559 ( .C (clk), .D (signal_8104), .Q (signal_8105) ) ;
    buf_clk cell_5575 ( .C (clk), .D (signal_8120), .Q (signal_8121) ) ;
    buf_clk cell_5591 ( .C (clk), .D (signal_8136), .Q (signal_8137) ) ;
    buf_clk cell_5607 ( .C (clk), .D (signal_8152), .Q (signal_8153) ) ;
    buf_clk cell_5623 ( .C (clk), .D (signal_8168), .Q (signal_8169) ) ;
    buf_clk cell_5639 ( .C (clk), .D (signal_8184), .Q (signal_8185) ) ;
    buf_clk cell_5655 ( .C (clk), .D (signal_8200), .Q (signal_8201) ) ;
    buf_clk cell_5671 ( .C (clk), .D (signal_8216), .Q (signal_8217) ) ;
    buf_clk cell_5687 ( .C (clk), .D (signal_8232), .Q (signal_8233) ) ;
    buf_clk cell_5703 ( .C (clk), .D (signal_8248), .Q (signal_8249) ) ;
    buf_clk cell_5719 ( .C (clk), .D (signal_8264), .Q (signal_8265) ) ;
    buf_clk cell_5735 ( .C (clk), .D (signal_8280), .Q (signal_8281) ) ;
    buf_clk cell_5751 ( .C (clk), .D (signal_8296), .Q (signal_8297) ) ;
    buf_clk cell_5767 ( .C (clk), .D (signal_8312), .Q (signal_8313) ) ;
    buf_clk cell_5783 ( .C (clk), .D (signal_8328), .Q (signal_8329) ) ;
    buf_clk cell_5799 ( .C (clk), .D (signal_8344), .Q (signal_8345) ) ;
    buf_clk cell_5815 ( .C (clk), .D (signal_8360), .Q (signal_8361) ) ;
    buf_clk cell_5831 ( .C (clk), .D (signal_8376), .Q (signal_8377) ) ;
    buf_clk cell_5847 ( .C (clk), .D (signal_8392), .Q (signal_8393) ) ;
    buf_clk cell_5863 ( .C (clk), .D (signal_8408), .Q (signal_8409) ) ;
    buf_clk cell_5879 ( .C (clk), .D (signal_8424), .Q (signal_8425) ) ;
    buf_clk cell_5895 ( .C (clk), .D (signal_8440), .Q (signal_8441) ) ;
    buf_clk cell_5911 ( .C (clk), .D (signal_8456), .Q (signal_8457) ) ;
    buf_clk cell_5927 ( .C (clk), .D (signal_8472), .Q (signal_8473) ) ;
    buf_clk cell_5943 ( .C (clk), .D (signal_8488), .Q (signal_8489) ) ;
    buf_clk cell_5959 ( .C (clk), .D (signal_8504), .Q (signal_8505) ) ;
    buf_clk cell_5975 ( .C (clk), .D (signal_8520), .Q (signal_8521) ) ;
    buf_clk cell_5991 ( .C (clk), .D (signal_8536), .Q (signal_8537) ) ;
    buf_clk cell_6007 ( .C (clk), .D (signal_8552), .Q (signal_8553) ) ;
    buf_clk cell_6023 ( .C (clk), .D (signal_8568), .Q (signal_8569) ) ;
    buf_clk cell_6039 ( .C (clk), .D (signal_8584), .Q (signal_8585) ) ;
    buf_clk cell_6055 ( .C (clk), .D (signal_8600), .Q (signal_8601) ) ;
    buf_clk cell_6071 ( .C (clk), .D (signal_8616), .Q (signal_8617) ) ;
    buf_clk cell_6087 ( .C (clk), .D (signal_8632), .Q (signal_8633) ) ;
    buf_clk cell_6103 ( .C (clk), .D (signal_8648), .Q (signal_8649) ) ;
    buf_clk cell_6119 ( .C (clk), .D (signal_8664), .Q (signal_8665) ) ;
    buf_clk cell_6135 ( .C (clk), .D (signal_8680), .Q (signal_8681) ) ;
    buf_clk cell_6151 ( .C (clk), .D (signal_8696), .Q (signal_8697) ) ;
    buf_clk cell_6167 ( .C (clk), .D (signal_8712), .Q (signal_8713) ) ;
    buf_clk cell_6183 ( .C (clk), .D (signal_8728), .Q (signal_8729) ) ;
    buf_clk cell_6199 ( .C (clk), .D (signal_8744), .Q (signal_8745) ) ;
    buf_clk cell_6215 ( .C (clk), .D (signal_8760), .Q (signal_8761) ) ;
    buf_clk cell_6231 ( .C (clk), .D (signal_8776), .Q (signal_8777) ) ;
    buf_clk cell_6247 ( .C (clk), .D (signal_8792), .Q (signal_8793) ) ;
    buf_clk cell_6263 ( .C (clk), .D (signal_8808), .Q (signal_8809) ) ;
    buf_clk cell_6279 ( .C (clk), .D (signal_8824), .Q (signal_8825) ) ;
    buf_clk cell_6295 ( .C (clk), .D (signal_8840), .Q (signal_8841) ) ;
    buf_clk cell_6311 ( .C (clk), .D (signal_8856), .Q (signal_8857) ) ;
    buf_clk cell_6327 ( .C (clk), .D (signal_8872), .Q (signal_8873) ) ;
    buf_clk cell_6343 ( .C (clk), .D (signal_8888), .Q (signal_8889) ) ;
    buf_clk cell_6359 ( .C (clk), .D (signal_8904), .Q (signal_8905) ) ;
    buf_clk cell_6375 ( .C (clk), .D (signal_8920), .Q (signal_8921) ) ;
    buf_clk cell_6391 ( .C (clk), .D (signal_8936), .Q (signal_8937) ) ;
    buf_clk cell_6407 ( .C (clk), .D (signal_8952), .Q (signal_8953) ) ;
    buf_clk cell_6423 ( .C (clk), .D (signal_8968), .Q (signal_8969) ) ;
    buf_clk cell_6439 ( .C (clk), .D (signal_8984), .Q (signal_8985) ) ;
    buf_clk cell_6455 ( .C (clk), .D (signal_9000), .Q (signal_9001) ) ;
    buf_clk cell_6471 ( .C (clk), .D (signal_9016), .Q (signal_9017) ) ;
    buf_clk cell_6487 ( .C (clk), .D (signal_9032), .Q (signal_9033) ) ;
    buf_clk cell_6503 ( .C (clk), .D (signal_9048), .Q (signal_9049) ) ;
    buf_clk cell_6519 ( .C (clk), .D (signal_9064), .Q (signal_9065) ) ;
    buf_clk cell_6535 ( .C (clk), .D (signal_9080), .Q (signal_9081) ) ;
    buf_clk cell_6551 ( .C (clk), .D (signal_9096), .Q (signal_9097) ) ;
    buf_clk cell_6567 ( .C (clk), .D (signal_9112), .Q (signal_9113) ) ;
    buf_clk cell_6583 ( .C (clk), .D (signal_9128), .Q (signal_9129) ) ;
    buf_clk cell_6599 ( .C (clk), .D (signal_9144), .Q (signal_9145) ) ;
    buf_clk cell_6615 ( .C (clk), .D (signal_9160), .Q (signal_9161) ) ;
    buf_clk cell_6631 ( .C (clk), .D (signal_9176), .Q (signal_9177) ) ;
    buf_clk cell_6647 ( .C (clk), .D (signal_9192), .Q (signal_9193) ) ;
    buf_clk cell_6663 ( .C (clk), .D (signal_9208), .Q (signal_9209) ) ;
    buf_clk cell_6679 ( .C (clk), .D (signal_9224), .Q (signal_9225) ) ;
    buf_clk cell_6695 ( .C (clk), .D (signal_9240), .Q (signal_9241) ) ;
    buf_clk cell_6711 ( .C (clk), .D (signal_9256), .Q (signal_9257) ) ;
    buf_clk cell_6727 ( .C (clk), .D (signal_9272), .Q (signal_9273) ) ;
    buf_clk cell_6743 ( .C (clk), .D (signal_9288), .Q (signal_9289) ) ;
    buf_clk cell_6759 ( .C (clk), .D (signal_9304), .Q (signal_9305) ) ;
    buf_clk cell_6775 ( .C (clk), .D (signal_9320), .Q (signal_9321) ) ;
    buf_clk cell_6791 ( .C (clk), .D (signal_9336), .Q (signal_9337) ) ;
    buf_clk cell_6807 ( .C (clk), .D (signal_9352), .Q (signal_9353) ) ;
    buf_clk cell_6823 ( .C (clk), .D (signal_9368), .Q (signal_9369) ) ;
    buf_clk cell_6839 ( .C (clk), .D (signal_9384), .Q (signal_9385) ) ;
    buf_clk cell_6855 ( .C (clk), .D (signal_9400), .Q (signal_9401) ) ;
    buf_clk cell_6871 ( .C (clk), .D (signal_9416), .Q (signal_9417) ) ;
    buf_clk cell_6887 ( .C (clk), .D (signal_9432), .Q (signal_9433) ) ;
    buf_clk cell_6903 ( .C (clk), .D (signal_9448), .Q (signal_9449) ) ;
    buf_clk cell_6919 ( .C (clk), .D (signal_9464), .Q (signal_9465) ) ;
    buf_clk cell_6935 ( .C (clk), .D (signal_9480), .Q (signal_9481) ) ;
    buf_clk cell_6951 ( .C (clk), .D (signal_9496), .Q (signal_9497) ) ;
    buf_clk cell_6967 ( .C (clk), .D (signal_9512), .Q (signal_9513) ) ;
    buf_clk cell_6983 ( .C (clk), .D (signal_9528), .Q (signal_9529) ) ;
    buf_clk cell_6999 ( .C (clk), .D (signal_9544), .Q (signal_9545) ) ;
    buf_clk cell_7015 ( .C (clk), .D (signal_9560), .Q (signal_9561) ) ;
    buf_clk cell_7031 ( .C (clk), .D (signal_9576), .Q (signal_9577) ) ;
    buf_clk cell_7047 ( .C (clk), .D (signal_9592), .Q (signal_9593) ) ;
    buf_clk cell_7063 ( .C (clk), .D (signal_9608), .Q (signal_9609) ) ;
    buf_clk cell_7079 ( .C (clk), .D (signal_9624), .Q (signal_9625) ) ;
    buf_clk cell_7095 ( .C (clk), .D (signal_9640), .Q (signal_9641) ) ;
    buf_clk cell_7111 ( .C (clk), .D (signal_9656), .Q (signal_9657) ) ;
    buf_clk cell_7127 ( .C (clk), .D (signal_9672), .Q (signal_9673) ) ;
    buf_clk cell_7143 ( .C (clk), .D (signal_9688), .Q (signal_9689) ) ;
    buf_clk cell_7159 ( .C (clk), .D (signal_9704), .Q (signal_9705) ) ;
    buf_clk cell_7175 ( .C (clk), .D (signal_9720), .Q (signal_9721) ) ;
    buf_clk cell_7191 ( .C (clk), .D (signal_9736), .Q (signal_9737) ) ;
    buf_clk cell_7207 ( .C (clk), .D (signal_9752), .Q (signal_9753) ) ;
    buf_clk cell_7223 ( .C (clk), .D (signal_9768), .Q (signal_9769) ) ;
    buf_clk cell_7239 ( .C (clk), .D (signal_9784), .Q (signal_9785) ) ;
    buf_clk cell_7255 ( .C (clk), .D (signal_9800), .Q (signal_9801) ) ;
    buf_clk cell_7271 ( .C (clk), .D (signal_9816), .Q (signal_9817) ) ;
    buf_clk cell_7287 ( .C (clk), .D (signal_9832), .Q (signal_9833) ) ;
    buf_clk cell_7303 ( .C (clk), .D (signal_9848), .Q (signal_9849) ) ;
    buf_clk cell_7319 ( .C (clk), .D (signal_9864), .Q (signal_9865) ) ;
    buf_clk cell_7335 ( .C (clk), .D (signal_9880), .Q (signal_9881) ) ;
    buf_clk cell_7351 ( .C (clk), .D (signal_9896), .Q (signal_9897) ) ;
    buf_clk cell_7367 ( .C (clk), .D (signal_9912), .Q (signal_9913) ) ;
    buf_clk cell_7383 ( .C (clk), .D (signal_9928), .Q (signal_9929) ) ;
    buf_clk cell_7399 ( .C (clk), .D (signal_9944), .Q (signal_9945) ) ;
    buf_clk cell_7415 ( .C (clk), .D (signal_9960), .Q (signal_9961) ) ;
    buf_clk cell_7431 ( .C (clk), .D (signal_9976), .Q (signal_9977) ) ;
    buf_clk cell_7447 ( .C (clk), .D (signal_9992), .Q (signal_9993) ) ;
    buf_clk cell_7463 ( .C (clk), .D (signal_10008), .Q (signal_10009) ) ;
    buf_clk cell_7479 ( .C (clk), .D (signal_10024), .Q (signal_10025) ) ;
    buf_clk cell_7495 ( .C (clk), .D (signal_10040), .Q (signal_10041) ) ;
    buf_clk cell_7511 ( .C (clk), .D (signal_10056), .Q (signal_10057) ) ;
    buf_clk cell_7527 ( .C (clk), .D (signal_10072), .Q (signal_10073) ) ;
    buf_clk cell_7543 ( .C (clk), .D (signal_10088), .Q (signal_10089) ) ;
    buf_clk cell_7559 ( .C (clk), .D (signal_10104), .Q (signal_10105) ) ;
    buf_clk cell_7575 ( .C (clk), .D (signal_10120), .Q (signal_10121) ) ;
    buf_clk cell_7591 ( .C (clk), .D (signal_10136), .Q (signal_10137) ) ;
    buf_clk cell_7607 ( .C (clk), .D (signal_10152), .Q (signal_10153) ) ;
    buf_clk cell_7623 ( .C (clk), .D (signal_10168), .Q (signal_10169) ) ;
    buf_clk cell_7639 ( .C (clk), .D (signal_10184), .Q (signal_10185) ) ;
    buf_clk cell_7655 ( .C (clk), .D (signal_10200), .Q (signal_10201) ) ;
    buf_clk cell_7671 ( .C (clk), .D (signal_10216), .Q (signal_10217) ) ;
    buf_clk cell_7687 ( .C (clk), .D (signal_10232), .Q (signal_10233) ) ;
    buf_clk cell_7703 ( .C (clk), .D (signal_10248), .Q (signal_10249) ) ;
    buf_clk cell_7719 ( .C (clk), .D (signal_10264), .Q (signal_10265) ) ;
    buf_clk cell_7735 ( .C (clk), .D (signal_10280), .Q (signal_10281) ) ;
    buf_clk cell_7751 ( .C (clk), .D (signal_10296), .Q (signal_10297) ) ;
    buf_clk cell_7767 ( .C (clk), .D (signal_10312), .Q (signal_10313) ) ;
    buf_clk cell_7783 ( .C (clk), .D (signal_10328), .Q (signal_10329) ) ;
    buf_clk cell_7799 ( .C (clk), .D (signal_10344), .Q (signal_10345) ) ;
    buf_clk cell_7815 ( .C (clk), .D (signal_10360), .Q (signal_10361) ) ;
    buf_clk cell_7831 ( .C (clk), .D (signal_10376), .Q (signal_10377) ) ;
    buf_clk cell_7847 ( .C (clk), .D (signal_10392), .Q (signal_10393) ) ;
    buf_clk cell_7863 ( .C (clk), .D (signal_10408), .Q (signal_10409) ) ;
    buf_clk cell_7879 ( .C (clk), .D (signal_10424), .Q (signal_10425) ) ;
    buf_clk cell_7895 ( .C (clk), .D (signal_10440), .Q (signal_10441) ) ;
    buf_clk cell_7911 ( .C (clk), .D (signal_10456), .Q (signal_10457) ) ;
    buf_clk cell_7927 ( .C (clk), .D (signal_10472), .Q (signal_10473) ) ;
    buf_clk cell_7943 ( .C (clk), .D (signal_10488), .Q (signal_10489) ) ;
    buf_clk cell_7959 ( .C (clk), .D (signal_10504), .Q (signal_10505) ) ;
    buf_clk cell_7975 ( .C (clk), .D (signal_10520), .Q (signal_10521) ) ;
    buf_clk cell_7991 ( .C (clk), .D (signal_10536), .Q (signal_10537) ) ;
    buf_clk cell_8007 ( .C (clk), .D (signal_10552), .Q (signal_10553) ) ;
    buf_clk cell_8023 ( .C (clk), .D (signal_10568), .Q (signal_10569) ) ;
    buf_clk cell_8039 ( .C (clk), .D (signal_10584), .Q (signal_10585) ) ;
    buf_clk cell_8055 ( .C (clk), .D (signal_10600), .Q (signal_10601) ) ;
    buf_clk cell_8071 ( .C (clk), .D (signal_10616), .Q (signal_10617) ) ;
    buf_clk cell_8087 ( .C (clk), .D (signal_10632), .Q (signal_10633) ) ;
    buf_clk cell_8103 ( .C (clk), .D (signal_10648), .Q (signal_10649) ) ;
    buf_clk cell_8119 ( .C (clk), .D (signal_10664), .Q (signal_10665) ) ;
    buf_clk cell_8135 ( .C (clk), .D (signal_10680), .Q (signal_10681) ) ;
    buf_clk cell_8151 ( .C (clk), .D (signal_10696), .Q (signal_10697) ) ;
    buf_clk cell_8167 ( .C (clk), .D (signal_10712), .Q (signal_10713) ) ;
    buf_clk cell_8183 ( .C (clk), .D (signal_10728), .Q (signal_10729) ) ;
    buf_clk cell_8199 ( .C (clk), .D (signal_10744), .Q (signal_10745) ) ;
    buf_clk cell_8215 ( .C (clk), .D (signal_10760), .Q (signal_10761) ) ;
    buf_clk cell_8231 ( .C (clk), .D (signal_10776), .Q (signal_10777) ) ;
    buf_clk cell_8247 ( .C (clk), .D (signal_10792), .Q (signal_10793) ) ;
    buf_clk cell_8263 ( .C (clk), .D (signal_10808), .Q (signal_10809) ) ;
    buf_clk cell_8279 ( .C (clk), .D (signal_10824), .Q (signal_10825) ) ;
    buf_clk cell_8295 ( .C (clk), .D (signal_10840), .Q (signal_10841) ) ;
    buf_clk cell_8311 ( .C (clk), .D (signal_10856), .Q (signal_10857) ) ;
    buf_clk cell_8327 ( .C (clk), .D (signal_10872), .Q (signal_10873) ) ;
    buf_clk cell_8343 ( .C (clk), .D (signal_10888), .Q (signal_10889) ) ;
    buf_clk cell_8359 ( .C (clk), .D (signal_10904), .Q (signal_10905) ) ;
    buf_clk cell_8375 ( .C (clk), .D (signal_10920), .Q (signal_10921) ) ;
    buf_clk cell_8391 ( .C (clk), .D (signal_10936), .Q (signal_10937) ) ;
    buf_clk cell_8407 ( .C (clk), .D (signal_10952), .Q (signal_10953) ) ;
    buf_clk cell_8423 ( .C (clk), .D (signal_10968), .Q (signal_10969) ) ;
    buf_clk cell_8439 ( .C (clk), .D (signal_10984), .Q (signal_10985) ) ;
    buf_clk cell_8455 ( .C (clk), .D (signal_11000), .Q (signal_11001) ) ;
    buf_clk cell_8471 ( .C (clk), .D (signal_11016), .Q (signal_11017) ) ;
    buf_clk cell_8487 ( .C (clk), .D (signal_11032), .Q (signal_11033) ) ;
    buf_clk cell_8503 ( .C (clk), .D (signal_11048), .Q (signal_11049) ) ;
    buf_clk cell_8519 ( .C (clk), .D (signal_11064), .Q (signal_11065) ) ;
    buf_clk cell_8535 ( .C (clk), .D (signal_11080), .Q (signal_11081) ) ;
    buf_clk cell_8551 ( .C (clk), .D (signal_11096), .Q (signal_11097) ) ;
    buf_clk cell_8567 ( .C (clk), .D (signal_11112), .Q (signal_11113) ) ;
    buf_clk cell_8583 ( .C (clk), .D (signal_11128), .Q (signal_11129) ) ;
    buf_clk cell_8599 ( .C (clk), .D (signal_11144), .Q (signal_11145) ) ;
    buf_clk cell_8615 ( .C (clk), .D (signal_11160), .Q (signal_11161) ) ;
    buf_clk cell_8631 ( .C (clk), .D (signal_11176), .Q (signal_11177) ) ;
    buf_clk cell_8647 ( .C (clk), .D (signal_11192), .Q (signal_11193) ) ;
    buf_clk cell_8663 ( .C (clk), .D (signal_11208), .Q (signal_11209) ) ;
    buf_clk cell_8679 ( .C (clk), .D (signal_11224), .Q (signal_11225) ) ;
    buf_clk cell_8695 ( .C (clk), .D (signal_11240), .Q (signal_11241) ) ;
    buf_clk cell_8711 ( .C (clk), .D (signal_11256), .Q (signal_11257) ) ;
    buf_clk cell_8727 ( .C (clk), .D (signal_11272), .Q (signal_11273) ) ;
    buf_clk cell_8743 ( .C (clk), .D (signal_11288), .Q (signal_11289) ) ;
    buf_clk cell_8759 ( .C (clk), .D (signal_11304), .Q (signal_11305) ) ;
    buf_clk cell_8775 ( .C (clk), .D (signal_11320), .Q (signal_11321) ) ;
    buf_clk cell_8791 ( .C (clk), .D (signal_11336), .Q (signal_11337) ) ;
    buf_clk cell_8807 ( .C (clk), .D (signal_11352), .Q (signal_11353) ) ;
    buf_clk cell_8823 ( .C (clk), .D (signal_11368), .Q (signal_11369) ) ;
    buf_clk cell_8839 ( .C (clk), .D (signal_11384), .Q (signal_11385) ) ;
    buf_clk cell_8855 ( .C (clk), .D (signal_11400), .Q (signal_11401) ) ;
    buf_clk cell_8871 ( .C (clk), .D (signal_11416), .Q (signal_11417) ) ;
    buf_clk cell_8887 ( .C (clk), .D (signal_11432), .Q (signal_11433) ) ;
    buf_clk cell_8903 ( .C (clk), .D (signal_11448), .Q (signal_11449) ) ;
    buf_clk cell_8919 ( .C (clk), .D (signal_11464), .Q (signal_11465) ) ;
    buf_clk cell_8935 ( .C (clk), .D (signal_11480), .Q (signal_11481) ) ;
    buf_clk cell_8951 ( .C (clk), .D (signal_11496), .Q (signal_11497) ) ;
    buf_clk cell_8967 ( .C (clk), .D (signal_11512), .Q (signal_11513) ) ;
    buf_clk cell_8983 ( .C (clk), .D (signal_11528), .Q (signal_11529) ) ;
    buf_clk cell_8999 ( .C (clk), .D (signal_11544), .Q (signal_11545) ) ;
    buf_clk cell_9015 ( .C (clk), .D (signal_11560), .Q (signal_11561) ) ;
    buf_clk cell_9031 ( .C (clk), .D (signal_11576), .Q (signal_11577) ) ;
    buf_clk cell_9047 ( .C (clk), .D (signal_11592), .Q (signal_11593) ) ;
    buf_clk cell_9063 ( .C (clk), .D (signal_11608), .Q (signal_11609) ) ;
    buf_clk cell_9079 ( .C (clk), .D (signal_11624), .Q (signal_11625) ) ;
    buf_clk cell_9095 ( .C (clk), .D (signal_11640), .Q (signal_11641) ) ;
    buf_clk cell_9111 ( .C (clk), .D (signal_11656), .Q (signal_11657) ) ;
    buf_clk cell_9127 ( .C (clk), .D (signal_11672), .Q (signal_11673) ) ;
    buf_clk cell_9143 ( .C (clk), .D (signal_11688), .Q (signal_11689) ) ;
    buf_clk cell_9159 ( .C (clk), .D (signal_11704), .Q (signal_11705) ) ;
    buf_clk cell_9175 ( .C (clk), .D (signal_11720), .Q (signal_11721) ) ;
    buf_clk cell_9191 ( .C (clk), .D (signal_11736), .Q (signal_11737) ) ;
    buf_clk cell_9207 ( .C (clk), .D (signal_11752), .Q (signal_11753) ) ;
    buf_clk cell_9223 ( .C (clk), .D (signal_11768), .Q (signal_11769) ) ;
    buf_clk cell_9239 ( .C (clk), .D (signal_11784), .Q (signal_11785) ) ;
    buf_clk cell_9255 ( .C (clk), .D (signal_11800), .Q (signal_11801) ) ;
    buf_clk cell_9271 ( .C (clk), .D (signal_11816), .Q (signal_11817) ) ;
    buf_clk cell_9287 ( .C (clk), .D (signal_11832), .Q (signal_11833) ) ;
    buf_clk cell_9303 ( .C (clk), .D (signal_11848), .Q (signal_11849) ) ;
    buf_clk cell_9319 ( .C (clk), .D (signal_11864), .Q (signal_11865) ) ;
    buf_clk cell_9335 ( .C (clk), .D (signal_11880), .Q (signal_11881) ) ;
    buf_clk cell_9351 ( .C (clk), .D (signal_11896), .Q (signal_11897) ) ;
    buf_clk cell_9367 ( .C (clk), .D (signal_11912), .Q (signal_11913) ) ;
    buf_clk cell_9383 ( .C (clk), .D (signal_11928), .Q (signal_11929) ) ;
    buf_clk cell_9399 ( .C (clk), .D (signal_11944), .Q (signal_11945) ) ;
    buf_clk cell_9415 ( .C (clk), .D (signal_11960), .Q (signal_11961) ) ;
    buf_clk cell_9431 ( .C (clk), .D (signal_11976), .Q (signal_11977) ) ;
    buf_clk cell_9447 ( .C (clk), .D (signal_11992), .Q (signal_11993) ) ;
    buf_clk cell_9463 ( .C (clk), .D (signal_12008), .Q (signal_12009) ) ;
    buf_clk cell_9479 ( .C (clk), .D (signal_12024), .Q (signal_12025) ) ;
    buf_clk cell_9495 ( .C (clk), .D (signal_12040), .Q (signal_12041) ) ;
    buf_clk cell_9511 ( .C (clk), .D (signal_12056), .Q (signal_12057) ) ;
    buf_clk cell_9527 ( .C (clk), .D (signal_12072), .Q (signal_12073) ) ;
    buf_clk cell_9543 ( .C (clk), .D (signal_12088), .Q (signal_12089) ) ;
    buf_clk cell_9559 ( .C (clk), .D (signal_12104), .Q (signal_12105) ) ;
    buf_clk cell_9575 ( .C (clk), .D (signal_12120), .Q (signal_12121) ) ;
    buf_clk cell_9591 ( .C (clk), .D (signal_12136), .Q (signal_12137) ) ;
    buf_clk cell_9607 ( .C (clk), .D (signal_12152), .Q (signal_12153) ) ;
    buf_clk cell_9623 ( .C (clk), .D (signal_12168), .Q (signal_12169) ) ;
    buf_clk cell_9639 ( .C (clk), .D (signal_12184), .Q (signal_12185) ) ;
    buf_clk cell_9655 ( .C (clk), .D (signal_12200), .Q (signal_12201) ) ;
    buf_clk cell_9671 ( .C (clk), .D (signal_12216), .Q (signal_12217) ) ;
    buf_clk cell_9687 ( .C (clk), .D (signal_12232), .Q (signal_12233) ) ;
    buf_clk cell_9703 ( .C (clk), .D (signal_12248), .Q (signal_12249) ) ;
    buf_clk cell_9719 ( .C (clk), .D (signal_12264), .Q (signal_12265) ) ;
    buf_clk cell_9735 ( .C (clk), .D (signal_12280), .Q (signal_12281) ) ;
    buf_clk cell_9751 ( .C (clk), .D (signal_12296), .Q (signal_12297) ) ;
    buf_clk cell_9767 ( .C (clk), .D (signal_12312), .Q (signal_12313) ) ;
    buf_clk cell_9783 ( .C (clk), .D (signal_12328), .Q (signal_12329) ) ;
    buf_clk cell_9799 ( .C (clk), .D (signal_12344), .Q (signal_12345) ) ;
    buf_clk cell_9815 ( .C (clk), .D (signal_12360), .Q (signal_12361) ) ;
    buf_clk cell_9831 ( .C (clk), .D (signal_12376), .Q (signal_12377) ) ;
    buf_clk cell_9847 ( .C (clk), .D (signal_12392), .Q (signal_12393) ) ;
    buf_clk cell_9863 ( .C (clk), .D (signal_12408), .Q (signal_12409) ) ;
    buf_clk cell_9879 ( .C (clk), .D (signal_12424), .Q (signal_12425) ) ;
    buf_clk cell_9895 ( .C (clk), .D (signal_12440), .Q (signal_12441) ) ;
    buf_clk cell_9911 ( .C (clk), .D (signal_12456), .Q (signal_12457) ) ;
    buf_clk cell_9927 ( .C (clk), .D (signal_12472), .Q (signal_12473) ) ;
    buf_clk cell_9943 ( .C (clk), .D (signal_12488), .Q (signal_12489) ) ;
    buf_clk cell_9959 ( .C (clk), .D (signal_12504), .Q (signal_12505) ) ;
    buf_clk cell_9975 ( .C (clk), .D (signal_12520), .Q (signal_12521) ) ;
    buf_clk cell_9991 ( .C (clk), .D (signal_12536), .Q (signal_12537) ) ;
    buf_clk cell_10007 ( .C (clk), .D (signal_12552), .Q (signal_12553) ) ;
    buf_clk cell_10023 ( .C (clk), .D (signal_12568), .Q (signal_12569) ) ;
    buf_clk cell_10039 ( .C (clk), .D (signal_12584), .Q (signal_12585) ) ;
    buf_clk cell_10055 ( .C (clk), .D (signal_12600), .Q (signal_12601) ) ;
    buf_clk cell_10071 ( .C (clk), .D (signal_12616), .Q (signal_12617) ) ;
    buf_clk cell_10087 ( .C (clk), .D (signal_12632), .Q (signal_12633) ) ;
    buf_clk cell_10103 ( .C (clk), .D (signal_12648), .Q (signal_12649) ) ;
    buf_clk cell_10119 ( .C (clk), .D (signal_12664), .Q (signal_12665) ) ;
    buf_clk cell_10135 ( .C (clk), .D (signal_12680), .Q (signal_12681) ) ;
    buf_clk cell_10151 ( .C (clk), .D (signal_12696), .Q (signal_12697) ) ;
    buf_clk cell_10167 ( .C (clk), .D (signal_12712), .Q (signal_12713) ) ;
    buf_clk cell_10183 ( .C (clk), .D (signal_12728), .Q (signal_12729) ) ;
    buf_clk cell_10199 ( .C (clk), .D (signal_12744), .Q (signal_12745) ) ;
    buf_clk cell_10215 ( .C (clk), .D (signal_12760), .Q (signal_12761) ) ;
    buf_clk cell_10231 ( .C (clk), .D (signal_12776), .Q (signal_12777) ) ;
    buf_clk cell_10247 ( .C (clk), .D (signal_12792), .Q (signal_12793) ) ;
    buf_clk cell_10263 ( .C (clk), .D (signal_12808), .Q (signal_12809) ) ;
    buf_clk cell_10279 ( .C (clk), .D (signal_12824), .Q (signal_12825) ) ;
    buf_clk cell_10295 ( .C (clk), .D (signal_12840), .Q (signal_12841) ) ;
    buf_clk cell_10311 ( .C (clk), .D (signal_12856), .Q (signal_12857) ) ;
    buf_clk cell_10327 ( .C (clk), .D (signal_12872), .Q (signal_12873) ) ;
    buf_clk cell_10343 ( .C (clk), .D (signal_12888), .Q (signal_12889) ) ;
    buf_clk cell_10359 ( .C (clk), .D (signal_12904), .Q (signal_12905) ) ;
    buf_clk cell_10375 ( .C (clk), .D (signal_12920), .Q (signal_12921) ) ;
    buf_clk cell_10391 ( .C (clk), .D (signal_12936), .Q (signal_12937) ) ;
    buf_clk cell_10407 ( .C (clk), .D (signal_12952), .Q (signal_12953) ) ;
    buf_clk cell_10423 ( .C (clk), .D (signal_12968), .Q (signal_12969) ) ;
    buf_clk cell_10439 ( .C (clk), .D (signal_12984), .Q (signal_12985) ) ;
    buf_clk cell_10455 ( .C (clk), .D (signal_13000), .Q (signal_13001) ) ;
    buf_clk cell_10471 ( .C (clk), .D (signal_13016), .Q (signal_13017) ) ;
    buf_clk cell_10487 ( .C (clk), .D (signal_13032), .Q (signal_13033) ) ;
    buf_clk cell_10503 ( .C (clk), .D (signal_13048), .Q (signal_13049) ) ;
    buf_clk cell_10519 ( .C (clk), .D (signal_13064), .Q (signal_13065) ) ;
    buf_clk cell_10535 ( .C (clk), .D (signal_13080), .Q (signal_13081) ) ;
    buf_clk cell_10551 ( .C (clk), .D (signal_13096), .Q (signal_13097) ) ;
    buf_clk cell_10567 ( .C (clk), .D (signal_13112), .Q (signal_13113) ) ;
    buf_clk cell_10583 ( .C (clk), .D (signal_13128), .Q (signal_13129) ) ;
    buf_clk cell_10599 ( .C (clk), .D (signal_13144), .Q (signal_13145) ) ;
    buf_clk cell_10615 ( .C (clk), .D (signal_13160), .Q (signal_13161) ) ;
    buf_clk cell_10631 ( .C (clk), .D (signal_13176), .Q (signal_13177) ) ;
    buf_clk cell_10647 ( .C (clk), .D (signal_13192), .Q (signal_13193) ) ;
    buf_clk cell_10663 ( .C (clk), .D (signal_13208), .Q (signal_13209) ) ;
    buf_clk cell_10679 ( .C (clk), .D (signal_13224), .Q (signal_13225) ) ;
    buf_clk cell_10695 ( .C (clk), .D (signal_13240), .Q (signal_13241) ) ;
    buf_clk cell_10711 ( .C (clk), .D (signal_13256), .Q (signal_13257) ) ;
    buf_clk cell_10727 ( .C (clk), .D (signal_13272), .Q (signal_13273) ) ;
    buf_clk cell_10743 ( .C (clk), .D (signal_13288), .Q (signal_13289) ) ;
    buf_clk cell_10759 ( .C (clk), .D (signal_13304), .Q (signal_13305) ) ;
    buf_clk cell_10775 ( .C (clk), .D (signal_13320), .Q (signal_13321) ) ;
    buf_clk cell_10791 ( .C (clk), .D (signal_13336), .Q (signal_13337) ) ;
    buf_clk cell_10807 ( .C (clk), .D (signal_13352), .Q (signal_13353) ) ;
    buf_clk cell_10823 ( .C (clk), .D (signal_13368), .Q (signal_13369) ) ;
    buf_clk cell_10839 ( .C (clk), .D (signal_13384), .Q (signal_13385) ) ;
    buf_clk cell_10855 ( .C (clk), .D (signal_13400), .Q (signal_13401) ) ;
    buf_clk cell_10871 ( .C (clk), .D (signal_13416), .Q (signal_13417) ) ;
    buf_clk cell_10887 ( .C (clk), .D (signal_13432), .Q (signal_13433) ) ;
    buf_clk cell_10903 ( .C (clk), .D (signal_13448), .Q (signal_13449) ) ;
    buf_clk cell_10919 ( .C (clk), .D (signal_13464), .Q (signal_13465) ) ;
    buf_clk cell_10935 ( .C (clk), .D (signal_13480), .Q (signal_13481) ) ;
    buf_clk cell_10951 ( .C (clk), .D (signal_13496), .Q (signal_13497) ) ;
    buf_clk cell_10967 ( .C (clk), .D (signal_13512), .Q (signal_13513) ) ;
    buf_clk cell_10983 ( .C (clk), .D (signal_13528), .Q (signal_13529) ) ;
    buf_clk cell_10999 ( .C (clk), .D (signal_13544), .Q (signal_13545) ) ;
    buf_clk cell_11015 ( .C (clk), .D (signal_13560), .Q (signal_13561) ) ;
    buf_clk cell_11031 ( .C (clk), .D (signal_13576), .Q (signal_13577) ) ;
    buf_clk cell_11047 ( .C (clk), .D (signal_13592), .Q (signal_13593) ) ;
    buf_clk cell_11063 ( .C (clk), .D (signal_13608), .Q (signal_13609) ) ;
    buf_clk cell_11079 ( .C (clk), .D (signal_13624), .Q (signal_13625) ) ;
    buf_clk cell_11095 ( .C (clk), .D (signal_13640), .Q (signal_13641) ) ;
    buf_clk cell_11111 ( .C (clk), .D (signal_13656), .Q (signal_13657) ) ;
    buf_clk cell_11127 ( .C (clk), .D (signal_13672), .Q (signal_13673) ) ;
    buf_clk cell_11143 ( .C (clk), .D (signal_13688), .Q (signal_13689) ) ;
    buf_clk cell_11159 ( .C (clk), .D (signal_13704), .Q (signal_13705) ) ;
    buf_clk cell_11175 ( .C (clk), .D (signal_13720), .Q (signal_13721) ) ;
    buf_clk cell_11191 ( .C (clk), .D (signal_13736), .Q (signal_13737) ) ;
    buf_clk cell_11207 ( .C (clk), .D (signal_13752), .Q (signal_13753) ) ;
    buf_clk cell_11223 ( .C (clk), .D (signal_13768), .Q (signal_13769) ) ;
    buf_clk cell_11239 ( .C (clk), .D (signal_13784), .Q (signal_13785) ) ;
    buf_clk cell_11255 ( .C (clk), .D (signal_13800), .Q (signal_13801) ) ;
    buf_clk cell_11271 ( .C (clk), .D (signal_13816), .Q (signal_13817) ) ;
    buf_clk cell_11287 ( .C (clk), .D (signal_13832), .Q (signal_13833) ) ;
    buf_clk cell_11303 ( .C (clk), .D (signal_13848), .Q (signal_13849) ) ;
    buf_clk cell_11319 ( .C (clk), .D (signal_13864), .Q (signal_13865) ) ;
    buf_clk cell_11335 ( .C (clk), .D (signal_13880), .Q (signal_13881) ) ;
    buf_clk cell_11351 ( .C (clk), .D (signal_13896), .Q (signal_13897) ) ;
    buf_clk cell_11367 ( .C (clk), .D (signal_13912), .Q (signal_13913) ) ;
    buf_clk cell_11383 ( .C (clk), .D (signal_13928), .Q (signal_13929) ) ;
    buf_clk cell_11399 ( .C (clk), .D (signal_13944), .Q (signal_13945) ) ;
    buf_clk cell_11415 ( .C (clk), .D (signal_13960), .Q (signal_13961) ) ;
    buf_clk cell_11431 ( .C (clk), .D (signal_13976), .Q (signal_13977) ) ;
    buf_clk cell_11447 ( .C (clk), .D (signal_13992), .Q (signal_13993) ) ;
    buf_clk cell_11463 ( .C (clk), .D (signal_14008), .Q (signal_14009) ) ;
    buf_clk cell_11479 ( .C (clk), .D (signal_14024), .Q (signal_14025) ) ;
    buf_clk cell_11495 ( .C (clk), .D (signal_14040), .Q (signal_14041) ) ;
    buf_clk cell_11511 ( .C (clk), .D (signal_14056), .Q (signal_14057) ) ;
    buf_clk cell_11527 ( .C (clk), .D (signal_14072), .Q (signal_14073) ) ;
    buf_clk cell_11543 ( .C (clk), .D (signal_14088), .Q (signal_14089) ) ;
    buf_clk cell_11559 ( .C (clk), .D (signal_14104), .Q (signal_14105) ) ;
    buf_clk cell_11575 ( .C (clk), .D (signal_14120), .Q (signal_14121) ) ;
    buf_clk cell_11591 ( .C (clk), .D (signal_14136), .Q (signal_14137) ) ;
    buf_clk cell_11607 ( .C (clk), .D (signal_14152), .Q (signal_14153) ) ;
    buf_clk cell_11623 ( .C (clk), .D (signal_14168), .Q (signal_14169) ) ;
    buf_clk cell_11639 ( .C (clk), .D (signal_14184), .Q (signal_14185) ) ;
    buf_clk cell_11655 ( .C (clk), .D (signal_14200), .Q (signal_14201) ) ;
    buf_clk cell_11671 ( .C (clk), .D (signal_14216), .Q (signal_14217) ) ;
    buf_clk cell_11687 ( .C (clk), .D (signal_14232), .Q (signal_14233) ) ;
    buf_clk cell_11703 ( .C (clk), .D (signal_14248), .Q (signal_14249) ) ;
    buf_clk cell_11719 ( .C (clk), .D (signal_14264), .Q (signal_14265) ) ;
    buf_clk cell_11735 ( .C (clk), .D (signal_14280), .Q (signal_14281) ) ;
    buf_clk cell_11751 ( .C (clk), .D (signal_14296), .Q (signal_14297) ) ;
    buf_clk cell_11767 ( .C (clk), .D (signal_14312), .Q (signal_14313) ) ;
    buf_clk cell_11783 ( .C (clk), .D (signal_14328), .Q (signal_14329) ) ;
    buf_clk cell_11799 ( .C (clk), .D (signal_14344), .Q (signal_14345) ) ;
    buf_clk cell_11815 ( .C (clk), .D (signal_14360), .Q (signal_14361) ) ;
    buf_clk cell_11831 ( .C (clk), .D (signal_14376), .Q (signal_14377) ) ;
    buf_clk cell_11847 ( .C (clk), .D (signal_14392), .Q (signal_14393) ) ;
    buf_clk cell_11863 ( .C (clk), .D (signal_14408), .Q (signal_14409) ) ;
    buf_clk cell_11879 ( .C (clk), .D (signal_14424), .Q (signal_14425) ) ;
    buf_clk cell_11895 ( .C (clk), .D (signal_14440), .Q (signal_14441) ) ;
    buf_clk cell_11911 ( .C (clk), .D (signal_14456), .Q (signal_14457) ) ;
    buf_clk cell_11927 ( .C (clk), .D (signal_14472), .Q (signal_14473) ) ;
    buf_clk cell_11943 ( .C (clk), .D (signal_14488), .Q (signal_14489) ) ;
    buf_clk cell_11959 ( .C (clk), .D (signal_14504), .Q (signal_14505) ) ;
    buf_clk cell_11975 ( .C (clk), .D (signal_14520), .Q (signal_14521) ) ;
    buf_clk cell_11991 ( .C (clk), .D (signal_14536), .Q (signal_14537) ) ;
    buf_clk cell_12007 ( .C (clk), .D (signal_14552), .Q (signal_14553) ) ;
    buf_clk cell_12023 ( .C (clk), .D (signal_14568), .Q (signal_14569) ) ;
    buf_clk cell_12039 ( .C (clk), .D (signal_14584), .Q (signal_14585) ) ;
    buf_clk cell_12055 ( .C (clk), .D (signal_14600), .Q (signal_14601) ) ;
    buf_clk cell_12071 ( .C (clk), .D (signal_14616), .Q (signal_14617) ) ;
    buf_clk cell_12087 ( .C (clk), .D (signal_14632), .Q (signal_14633) ) ;
    buf_clk cell_12103 ( .C (clk), .D (signal_14648), .Q (signal_14649) ) ;
    buf_clk cell_12119 ( .C (clk), .D (signal_14664), .Q (signal_14665) ) ;
    buf_clk cell_12135 ( .C (clk), .D (signal_14680), .Q (signal_14681) ) ;
    buf_clk cell_12151 ( .C (clk), .D (signal_14696), .Q (signal_14697) ) ;
    buf_clk cell_12167 ( .C (clk), .D (signal_14712), .Q (signal_14713) ) ;
    buf_clk cell_12183 ( .C (clk), .D (signal_14728), .Q (signal_14729) ) ;
    buf_clk cell_12199 ( .C (clk), .D (signal_14744), .Q (signal_14745) ) ;
    buf_clk cell_12215 ( .C (clk), .D (signal_14760), .Q (signal_14761) ) ;
    buf_clk cell_12231 ( .C (clk), .D (signal_14776), .Q (signal_14777) ) ;
    buf_clk cell_12247 ( .C (clk), .D (signal_14792), .Q (signal_14793) ) ;
    buf_clk cell_12263 ( .C (clk), .D (signal_14808), .Q (signal_14809) ) ;
    buf_clk cell_12279 ( .C (clk), .D (signal_14824), .Q (signal_14825) ) ;
    buf_clk cell_12295 ( .C (clk), .D (signal_14840), .Q (signal_14841) ) ;
    buf_clk cell_12311 ( .C (clk), .D (signal_14856), .Q (signal_14857) ) ;
    buf_clk cell_12327 ( .C (clk), .D (signal_14872), .Q (signal_14873) ) ;
    buf_clk cell_12343 ( .C (clk), .D (signal_14888), .Q (signal_14889) ) ;
    buf_clk cell_12359 ( .C (clk), .D (signal_14904), .Q (signal_14905) ) ;
    buf_clk cell_12375 ( .C (clk), .D (signal_14920), .Q (signal_14921) ) ;
    buf_clk cell_12391 ( .C (clk), .D (signal_14936), .Q (signal_14937) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2089 ( .s ({signal_4906, signal_4896}), .b ({signal_3957, signal_2294}), .a ({signal_3956, signal_2293}), .clk (clk), .r (Fresh[375]), .c ({signal_4124, signal_2357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2090 ( .s ({signal_4906, signal_4896}), .b ({signal_3959, signal_2296}), .a ({signal_3958, signal_2295}), .clk (clk), .r (Fresh[376]), .c ({signal_4125, signal_2358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2091 ( .s ({signal_4906, signal_4896}), .b ({signal_3961, signal_2298}), .a ({signal_3960, signal_2297}), .clk (clk), .r (Fresh[377]), .c ({signal_4126, signal_2359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2092 ( .s ({signal_4906, signal_4896}), .b ({signal_3963, signal_2300}), .a ({signal_3962, signal_2299}), .clk (clk), .r (Fresh[378]), .c ({signal_4127, signal_2360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2093 ( .s ({signal_4906, signal_4896}), .b ({signal_3965, signal_2302}), .a ({signal_3964, signal_2301}), .clk (clk), .r (Fresh[379]), .c ({signal_4128, signal_2361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2094 ( .s ({signal_4906, signal_4896}), .b ({signal_3967, signal_2304}), .a ({signal_3966, signal_2303}), .clk (clk), .r (Fresh[380]), .c ({signal_4129, signal_2362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2095 ( .s ({signal_4906, signal_4896}), .b ({signal_3969, signal_2306}), .a ({signal_3968, signal_2305}), .clk (clk), .r (Fresh[381]), .c ({signal_4130, signal_2363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2096 ( .s ({signal_4906, signal_4896}), .b ({signal_3971, signal_2308}), .a ({signal_3970, signal_2307}), .clk (clk), .r (Fresh[382]), .c ({signal_4131, signal_2364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2097 ( .s ({signal_4906, signal_4896}), .b ({signal_3973, signal_2310}), .a ({signal_3972, signal_2309}), .clk (clk), .r (Fresh[383]), .c ({signal_4132, signal_2365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2098 ( .s ({signal_4906, signal_4896}), .b ({signal_3975, signal_2312}), .a ({signal_3974, signal_2311}), .clk (clk), .r (Fresh[384]), .c ({signal_4133, signal_2366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2099 ( .s ({signal_4906, signal_4896}), .b ({signal_3977, signal_2314}), .a ({signal_3976, signal_2313}), .clk (clk), .r (Fresh[385]), .c ({signal_4134, signal_2367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2100 ( .s ({signal_4906, signal_4896}), .b ({signal_3979, signal_2316}), .a ({signal_3978, signal_2315}), .clk (clk), .r (Fresh[386]), .c ({signal_4135, signal_2368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2101 ( .s ({signal_4906, signal_4896}), .b ({signal_3981, signal_2318}), .a ({signal_3980, signal_2317}), .clk (clk), .r (Fresh[387]), .c ({signal_4136, signal_2369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2102 ( .s ({signal_4906, signal_4896}), .b ({signal_3983, signal_2320}), .a ({signal_3982, signal_2319}), .clk (clk), .r (Fresh[388]), .c ({signal_4137, signal_2370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2103 ( .s ({signal_4906, signal_4896}), .b ({signal_3985, signal_2322}), .a ({signal_3984, signal_2321}), .clk (clk), .r (Fresh[389]), .c ({signal_4138, signal_2371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2104 ( .s ({signal_4906, signal_4896}), .b ({signal_3987, signal_2324}), .a ({signal_3986, signal_2323}), .clk (clk), .r (Fresh[390]), .c ({signal_4139, signal_2372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2105 ( .s ({signal_4906, signal_4896}), .b ({signal_3989, signal_2326}), .a ({signal_3988, signal_2325}), .clk (clk), .r (Fresh[391]), .c ({signal_4140, signal_2373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2106 ( .s ({signal_4906, signal_4896}), .b ({signal_3991, signal_2328}), .a ({signal_3990, signal_2327}), .clk (clk), .r (Fresh[392]), .c ({signal_4141, signal_2374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2107 ( .s ({signal_4906, signal_4896}), .b ({signal_3993, signal_2330}), .a ({signal_3992, signal_2329}), .clk (clk), .r (Fresh[393]), .c ({signal_4142, signal_2375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2108 ( .s ({signal_4906, signal_4896}), .b ({signal_3995, signal_2332}), .a ({signal_3994, signal_2331}), .clk (clk), .r (Fresh[394]), .c ({signal_4143, signal_2376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2109 ( .s ({signal_4906, signal_4896}), .b ({signal_3997, signal_2334}), .a ({signal_3996, signal_2333}), .clk (clk), .r (Fresh[395]), .c ({signal_4144, signal_2377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2110 ( .s ({signal_4906, signal_4896}), .b ({signal_3999, signal_2336}), .a ({signal_3998, signal_2335}), .clk (clk), .r (Fresh[396]), .c ({signal_4145, signal_2378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2111 ( .s ({signal_4906, signal_4896}), .b ({signal_4001, signal_2338}), .a ({signal_4000, signal_2337}), .clk (clk), .r (Fresh[397]), .c ({signal_4146, signal_2379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2112 ( .s ({signal_4906, signal_4896}), .b ({signal_4003, signal_2340}), .a ({signal_4002, signal_2339}), .clk (clk), .r (Fresh[398]), .c ({signal_4147, signal_2380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2113 ( .s ({signal_4906, signal_4896}), .b ({signal_4005, signal_2342}), .a ({signal_4004, signal_2341}), .clk (clk), .r (Fresh[399]), .c ({signal_4148, signal_2381}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2114 ( .s ({signal_4906, signal_4896}), .b ({signal_4007, signal_2344}), .a ({signal_4006, signal_2343}), .clk (clk), .r (Fresh[400]), .c ({signal_4149, signal_2382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2115 ( .s ({signal_4906, signal_4896}), .b ({signal_4009, signal_2346}), .a ({signal_4008, signal_2345}), .clk (clk), .r (Fresh[401]), .c ({signal_4150, signal_2383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2116 ( .s ({signal_4906, signal_4896}), .b ({signal_4011, signal_2348}), .a ({signal_4010, signal_2347}), .clk (clk), .r (Fresh[402]), .c ({signal_4151, signal_2384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2117 ( .s ({signal_4906, signal_4896}), .b ({signal_4013, signal_2350}), .a ({signal_4012, signal_2349}), .clk (clk), .r (Fresh[403]), .c ({signal_4152, signal_2385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2118 ( .s ({signal_4906, signal_4896}), .b ({signal_4015, signal_2352}), .a ({signal_4014, signal_2351}), .clk (clk), .r (Fresh[404]), .c ({signal_4153, signal_2386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2119 ( .s ({signal_4906, signal_4896}), .b ({signal_4017, signal_2354}), .a ({signal_4016, signal_2353}), .clk (clk), .r (Fresh[405]), .c ({signal_4154, signal_2387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2120 ( .s ({signal_4906, signal_4896}), .b ({signal_4019, signal_2356}), .a ({signal_4018, signal_2355}), .clk (clk), .r (Fresh[406]), .c ({signal_4155, signal_2388}) ) ;
    buf_clk cell_2372 ( .C (clk), .D (signal_4917), .Q (signal_4918) ) ;
    buf_clk cell_2384 ( .C (clk), .D (signal_4929), .Q (signal_4930) ) ;
    buf_clk cell_2396 ( .C (clk), .D (signal_4941), .Q (signal_4942) ) ;
    buf_clk cell_2412 ( .C (clk), .D (signal_4957), .Q (signal_4958) ) ;
    buf_clk cell_2428 ( .C (clk), .D (signal_4973), .Q (signal_4974) ) ;
    buf_clk cell_2444 ( .C (clk), .D (signal_4989), .Q (signal_4990) ) ;
    buf_clk cell_2460 ( .C (clk), .D (signal_5005), .Q (signal_5006) ) ;
    buf_clk cell_2476 ( .C (clk), .D (signal_5021), .Q (signal_5022) ) ;
    buf_clk cell_2492 ( .C (clk), .D (signal_5037), .Q (signal_5038) ) ;
    buf_clk cell_2508 ( .C (clk), .D (signal_5053), .Q (signal_5054) ) ;
    buf_clk cell_2524 ( .C (clk), .D (signal_5069), .Q (signal_5070) ) ;
    buf_clk cell_2540 ( .C (clk), .D (signal_5085), .Q (signal_5086) ) ;
    buf_clk cell_2556 ( .C (clk), .D (signal_5101), .Q (signal_5102) ) ;
    buf_clk cell_2572 ( .C (clk), .D (signal_5117), .Q (signal_5118) ) ;
    buf_clk cell_2588 ( .C (clk), .D (signal_5133), .Q (signal_5134) ) ;
    buf_clk cell_2604 ( .C (clk), .D (signal_5149), .Q (signal_5150) ) ;
    buf_clk cell_2620 ( .C (clk), .D (signal_5165), .Q (signal_5166) ) ;
    buf_clk cell_2636 ( .C (clk), .D (signal_5181), .Q (signal_5182) ) ;
    buf_clk cell_2652 ( .C (clk), .D (signal_5197), .Q (signal_5198) ) ;
    buf_clk cell_2668 ( .C (clk), .D (signal_5213), .Q (signal_5214) ) ;
    buf_clk cell_2684 ( .C (clk), .D (signal_5229), .Q (signal_5230) ) ;
    buf_clk cell_2700 ( .C (clk), .D (signal_5245), .Q (signal_5246) ) ;
    buf_clk cell_2716 ( .C (clk), .D (signal_5261), .Q (signal_5262) ) ;
    buf_clk cell_2732 ( .C (clk), .D (signal_5277), .Q (signal_5278) ) ;
    buf_clk cell_2748 ( .C (clk), .D (signal_5293), .Q (signal_5294) ) ;
    buf_clk cell_2764 ( .C (clk), .D (signal_5309), .Q (signal_5310) ) ;
    buf_clk cell_2780 ( .C (clk), .D (signal_5325), .Q (signal_5326) ) ;
    buf_clk cell_2796 ( .C (clk), .D (signal_5341), .Q (signal_5342) ) ;
    buf_clk cell_2812 ( .C (clk), .D (signal_5357), .Q (signal_5358) ) ;
    buf_clk cell_2828 ( .C (clk), .D (signal_5373), .Q (signal_5374) ) ;
    buf_clk cell_2844 ( .C (clk), .D (signal_5389), .Q (signal_5390) ) ;
    buf_clk cell_2860 ( .C (clk), .D (signal_5405), .Q (signal_5406) ) ;
    buf_clk cell_2876 ( .C (clk), .D (signal_5421), .Q (signal_5422) ) ;
    buf_clk cell_2892 ( .C (clk), .D (signal_5437), .Q (signal_5438) ) ;
    buf_clk cell_2908 ( .C (clk), .D (signal_5453), .Q (signal_5454) ) ;
    buf_clk cell_2924 ( .C (clk), .D (signal_5469), .Q (signal_5470) ) ;
    buf_clk cell_2940 ( .C (clk), .D (signal_5485), .Q (signal_5486) ) ;
    buf_clk cell_2956 ( .C (clk), .D (signal_5501), .Q (signal_5502) ) ;
    buf_clk cell_2972 ( .C (clk), .D (signal_5517), .Q (signal_5518) ) ;
    buf_clk cell_2988 ( .C (clk), .D (signal_5533), .Q (signal_5534) ) ;
    buf_clk cell_3004 ( .C (clk), .D (signal_5549), .Q (signal_5550) ) ;
    buf_clk cell_3020 ( .C (clk), .D (signal_5565), .Q (signal_5566) ) ;
    buf_clk cell_3036 ( .C (clk), .D (signal_5581), .Q (signal_5582) ) ;
    buf_clk cell_3052 ( .C (clk), .D (signal_5597), .Q (signal_5598) ) ;
    buf_clk cell_3068 ( .C (clk), .D (signal_5613), .Q (signal_5614) ) ;
    buf_clk cell_3084 ( .C (clk), .D (signal_5629), .Q (signal_5630) ) ;
    buf_clk cell_3100 ( .C (clk), .D (signal_5645), .Q (signal_5646) ) ;
    buf_clk cell_3116 ( .C (clk), .D (signal_5661), .Q (signal_5662) ) ;
    buf_clk cell_3132 ( .C (clk), .D (signal_5677), .Q (signal_5678) ) ;
    buf_clk cell_3148 ( .C (clk), .D (signal_5693), .Q (signal_5694) ) ;
    buf_clk cell_3164 ( .C (clk), .D (signal_5709), .Q (signal_5710) ) ;
    buf_clk cell_3180 ( .C (clk), .D (signal_5725), .Q (signal_5726) ) ;
    buf_clk cell_3196 ( .C (clk), .D (signal_5741), .Q (signal_5742) ) ;
    buf_clk cell_3212 ( .C (clk), .D (signal_5757), .Q (signal_5758) ) ;
    buf_clk cell_3228 ( .C (clk), .D (signal_5773), .Q (signal_5774) ) ;
    buf_clk cell_3244 ( .C (clk), .D (signal_5789), .Q (signal_5790) ) ;
    buf_clk cell_3260 ( .C (clk), .D (signal_5805), .Q (signal_5806) ) ;
    buf_clk cell_3276 ( .C (clk), .D (signal_5821), .Q (signal_5822) ) ;
    buf_clk cell_3292 ( .C (clk), .D (signal_5837), .Q (signal_5838) ) ;
    buf_clk cell_3308 ( .C (clk), .D (signal_5853), .Q (signal_5854) ) ;
    buf_clk cell_3324 ( .C (clk), .D (signal_5869), .Q (signal_5870) ) ;
    buf_clk cell_3340 ( .C (clk), .D (signal_5885), .Q (signal_5886) ) ;
    buf_clk cell_3356 ( .C (clk), .D (signal_5901), .Q (signal_5902) ) ;
    buf_clk cell_3372 ( .C (clk), .D (signal_5917), .Q (signal_5918) ) ;
    buf_clk cell_3388 ( .C (clk), .D (signal_5933), .Q (signal_5934) ) ;
    buf_clk cell_3404 ( .C (clk), .D (signal_5949), .Q (signal_5950) ) ;
    buf_clk cell_3420 ( .C (clk), .D (signal_5965), .Q (signal_5966) ) ;
    buf_clk cell_3436 ( .C (clk), .D (signal_5981), .Q (signal_5982) ) ;
    buf_clk cell_3452 ( .C (clk), .D (signal_5997), .Q (signal_5998) ) ;
    buf_clk cell_3468 ( .C (clk), .D (signal_6013), .Q (signal_6014) ) ;
    buf_clk cell_3484 ( .C (clk), .D (signal_6029), .Q (signal_6030) ) ;
    buf_clk cell_3500 ( .C (clk), .D (signal_6045), .Q (signal_6046) ) ;
    buf_clk cell_3516 ( .C (clk), .D (signal_6061), .Q (signal_6062) ) ;
    buf_clk cell_3532 ( .C (clk), .D (signal_6077), .Q (signal_6078) ) ;
    buf_clk cell_3548 ( .C (clk), .D (signal_6093), .Q (signal_6094) ) ;
    buf_clk cell_3564 ( .C (clk), .D (signal_6109), .Q (signal_6110) ) ;
    buf_clk cell_3580 ( .C (clk), .D (signal_6125), .Q (signal_6126) ) ;
    buf_clk cell_3596 ( .C (clk), .D (signal_6141), .Q (signal_6142) ) ;
    buf_clk cell_3612 ( .C (clk), .D (signal_6157), .Q (signal_6158) ) ;
    buf_clk cell_3628 ( .C (clk), .D (signal_6173), .Q (signal_6174) ) ;
    buf_clk cell_3644 ( .C (clk), .D (signal_6189), .Q (signal_6190) ) ;
    buf_clk cell_3660 ( .C (clk), .D (signal_6205), .Q (signal_6206) ) ;
    buf_clk cell_3676 ( .C (clk), .D (signal_6221), .Q (signal_6222) ) ;
    buf_clk cell_3692 ( .C (clk), .D (signal_6237), .Q (signal_6238) ) ;
    buf_clk cell_3708 ( .C (clk), .D (signal_6253), .Q (signal_6254) ) ;
    buf_clk cell_3724 ( .C (clk), .D (signal_6269), .Q (signal_6270) ) ;
    buf_clk cell_3740 ( .C (clk), .D (signal_6285), .Q (signal_6286) ) ;
    buf_clk cell_3756 ( .C (clk), .D (signal_6301), .Q (signal_6302) ) ;
    buf_clk cell_3772 ( .C (clk), .D (signal_6317), .Q (signal_6318) ) ;
    buf_clk cell_3788 ( .C (clk), .D (signal_6333), .Q (signal_6334) ) ;
    buf_clk cell_3804 ( .C (clk), .D (signal_6349), .Q (signal_6350) ) ;
    buf_clk cell_3820 ( .C (clk), .D (signal_6365), .Q (signal_6366) ) ;
    buf_clk cell_3836 ( .C (clk), .D (signal_6381), .Q (signal_6382) ) ;
    buf_clk cell_3852 ( .C (clk), .D (signal_6397), .Q (signal_6398) ) ;
    buf_clk cell_3868 ( .C (clk), .D (signal_6413), .Q (signal_6414) ) ;
    buf_clk cell_3884 ( .C (clk), .D (signal_6429), .Q (signal_6430) ) ;
    buf_clk cell_3900 ( .C (clk), .D (signal_6445), .Q (signal_6446) ) ;
    buf_clk cell_3916 ( .C (clk), .D (signal_6461), .Q (signal_6462) ) ;
    buf_clk cell_3932 ( .C (clk), .D (signal_6477), .Q (signal_6478) ) ;
    buf_clk cell_3948 ( .C (clk), .D (signal_6493), .Q (signal_6494) ) ;
    buf_clk cell_3964 ( .C (clk), .D (signal_6509), .Q (signal_6510) ) ;
    buf_clk cell_3980 ( .C (clk), .D (signal_6525), .Q (signal_6526) ) ;
    buf_clk cell_3996 ( .C (clk), .D (signal_6541), .Q (signal_6542) ) ;
    buf_clk cell_4012 ( .C (clk), .D (signal_6557), .Q (signal_6558) ) ;
    buf_clk cell_4028 ( .C (clk), .D (signal_6573), .Q (signal_6574) ) ;
    buf_clk cell_4044 ( .C (clk), .D (signal_6589), .Q (signal_6590) ) ;
    buf_clk cell_4060 ( .C (clk), .D (signal_6605), .Q (signal_6606) ) ;
    buf_clk cell_4076 ( .C (clk), .D (signal_6621), .Q (signal_6622) ) ;
    buf_clk cell_4092 ( .C (clk), .D (signal_6637), .Q (signal_6638) ) ;
    buf_clk cell_4108 ( .C (clk), .D (signal_6653), .Q (signal_6654) ) ;
    buf_clk cell_4124 ( .C (clk), .D (signal_6669), .Q (signal_6670) ) ;
    buf_clk cell_4140 ( .C (clk), .D (signal_6685), .Q (signal_6686) ) ;
    buf_clk cell_4156 ( .C (clk), .D (signal_6701), .Q (signal_6702) ) ;
    buf_clk cell_4172 ( .C (clk), .D (signal_6717), .Q (signal_6718) ) ;
    buf_clk cell_4188 ( .C (clk), .D (signal_6733), .Q (signal_6734) ) ;
    buf_clk cell_4204 ( .C (clk), .D (signal_6749), .Q (signal_6750) ) ;
    buf_clk cell_4220 ( .C (clk), .D (signal_6765), .Q (signal_6766) ) ;
    buf_clk cell_4236 ( .C (clk), .D (signal_6781), .Q (signal_6782) ) ;
    buf_clk cell_4252 ( .C (clk), .D (signal_6797), .Q (signal_6798) ) ;
    buf_clk cell_4268 ( .C (clk), .D (signal_6813), .Q (signal_6814) ) ;
    buf_clk cell_4284 ( .C (clk), .D (signal_6829), .Q (signal_6830) ) ;
    buf_clk cell_4300 ( .C (clk), .D (signal_6845), .Q (signal_6846) ) ;
    buf_clk cell_4316 ( .C (clk), .D (signal_6861), .Q (signal_6862) ) ;
    buf_clk cell_4332 ( .C (clk), .D (signal_6877), .Q (signal_6878) ) ;
    buf_clk cell_4348 ( .C (clk), .D (signal_6893), .Q (signal_6894) ) ;
    buf_clk cell_4364 ( .C (clk), .D (signal_6909), .Q (signal_6910) ) ;
    buf_clk cell_4380 ( .C (clk), .D (signal_6925), .Q (signal_6926) ) ;
    buf_clk cell_4396 ( .C (clk), .D (signal_6941), .Q (signal_6942) ) ;
    buf_clk cell_4412 ( .C (clk), .D (signal_6957), .Q (signal_6958) ) ;
    buf_clk cell_4426 ( .C (clk), .D (signal_6971), .Q (signal_6972) ) ;
    buf_clk cell_4440 ( .C (clk), .D (signal_6985), .Q (signal_6986) ) ;
    buf_clk cell_4456 ( .C (clk), .D (signal_7001), .Q (signal_7002) ) ;
    buf_clk cell_4472 ( .C (clk), .D (signal_7017), .Q (signal_7018) ) ;
    buf_clk cell_4488 ( .C (clk), .D (signal_7033), .Q (signal_7034) ) ;
    buf_clk cell_4504 ( .C (clk), .D (signal_7049), .Q (signal_7050) ) ;
    buf_clk cell_4520 ( .C (clk), .D (signal_7065), .Q (signal_7066) ) ;
    buf_clk cell_4536 ( .C (clk), .D (signal_7081), .Q (signal_7082) ) ;
    buf_clk cell_4552 ( .C (clk), .D (signal_7097), .Q (signal_7098) ) ;
    buf_clk cell_4568 ( .C (clk), .D (signal_7113), .Q (signal_7114) ) ;
    buf_clk cell_4584 ( .C (clk), .D (signal_7129), .Q (signal_7130) ) ;
    buf_clk cell_4600 ( .C (clk), .D (signal_7145), .Q (signal_7146) ) ;
    buf_clk cell_4616 ( .C (clk), .D (signal_7161), .Q (signal_7162) ) ;
    buf_clk cell_4632 ( .C (clk), .D (signal_7177), .Q (signal_7178) ) ;
    buf_clk cell_4648 ( .C (clk), .D (signal_7193), .Q (signal_7194) ) ;
    buf_clk cell_4664 ( .C (clk), .D (signal_7209), .Q (signal_7210) ) ;
    buf_clk cell_4680 ( .C (clk), .D (signal_7225), .Q (signal_7226) ) ;
    buf_clk cell_4696 ( .C (clk), .D (signal_7241), .Q (signal_7242) ) ;
    buf_clk cell_4712 ( .C (clk), .D (signal_7257), .Q (signal_7258) ) ;
    buf_clk cell_4728 ( .C (clk), .D (signal_7273), .Q (signal_7274) ) ;
    buf_clk cell_4744 ( .C (clk), .D (signal_7289), .Q (signal_7290) ) ;
    buf_clk cell_4760 ( .C (clk), .D (signal_7305), .Q (signal_7306) ) ;
    buf_clk cell_4776 ( .C (clk), .D (signal_7321), .Q (signal_7322) ) ;
    buf_clk cell_4792 ( .C (clk), .D (signal_7337), .Q (signal_7338) ) ;
    buf_clk cell_4808 ( .C (clk), .D (signal_7353), .Q (signal_7354) ) ;
    buf_clk cell_4824 ( .C (clk), .D (signal_7369), .Q (signal_7370) ) ;
    buf_clk cell_4840 ( .C (clk), .D (signal_7385), .Q (signal_7386) ) ;
    buf_clk cell_4856 ( .C (clk), .D (signal_7401), .Q (signal_7402) ) ;
    buf_clk cell_4872 ( .C (clk), .D (signal_7417), .Q (signal_7418) ) ;
    buf_clk cell_4888 ( .C (clk), .D (signal_7433), .Q (signal_7434) ) ;
    buf_clk cell_4904 ( .C (clk), .D (signal_7449), .Q (signal_7450) ) ;
    buf_clk cell_4920 ( .C (clk), .D (signal_7465), .Q (signal_7466) ) ;
    buf_clk cell_4936 ( .C (clk), .D (signal_7481), .Q (signal_7482) ) ;
    buf_clk cell_4952 ( .C (clk), .D (signal_7497), .Q (signal_7498) ) ;
    buf_clk cell_4968 ( .C (clk), .D (signal_7513), .Q (signal_7514) ) ;
    buf_clk cell_4984 ( .C (clk), .D (signal_7529), .Q (signal_7530) ) ;
    buf_clk cell_5000 ( .C (clk), .D (signal_7545), .Q (signal_7546) ) ;
    buf_clk cell_5016 ( .C (clk), .D (signal_7561), .Q (signal_7562) ) ;
    buf_clk cell_5032 ( .C (clk), .D (signal_7577), .Q (signal_7578) ) ;
    buf_clk cell_5048 ( .C (clk), .D (signal_7593), .Q (signal_7594) ) ;
    buf_clk cell_5064 ( .C (clk), .D (signal_7609), .Q (signal_7610) ) ;
    buf_clk cell_5080 ( .C (clk), .D (signal_7625), .Q (signal_7626) ) ;
    buf_clk cell_5096 ( .C (clk), .D (signal_7641), .Q (signal_7642) ) ;
    buf_clk cell_5112 ( .C (clk), .D (signal_7657), .Q (signal_7658) ) ;
    buf_clk cell_5128 ( .C (clk), .D (signal_7673), .Q (signal_7674) ) ;
    buf_clk cell_5144 ( .C (clk), .D (signal_7689), .Q (signal_7690) ) ;
    buf_clk cell_5160 ( .C (clk), .D (signal_7705), .Q (signal_7706) ) ;
    buf_clk cell_5176 ( .C (clk), .D (signal_7721), .Q (signal_7722) ) ;
    buf_clk cell_5192 ( .C (clk), .D (signal_7737), .Q (signal_7738) ) ;
    buf_clk cell_5208 ( .C (clk), .D (signal_7753), .Q (signal_7754) ) ;
    buf_clk cell_5224 ( .C (clk), .D (signal_7769), .Q (signal_7770) ) ;
    buf_clk cell_5240 ( .C (clk), .D (signal_7785), .Q (signal_7786) ) ;
    buf_clk cell_5256 ( .C (clk), .D (signal_7801), .Q (signal_7802) ) ;
    buf_clk cell_5272 ( .C (clk), .D (signal_7817), .Q (signal_7818) ) ;
    buf_clk cell_5288 ( .C (clk), .D (signal_7833), .Q (signal_7834) ) ;
    buf_clk cell_5304 ( .C (clk), .D (signal_7849), .Q (signal_7850) ) ;
    buf_clk cell_5320 ( .C (clk), .D (signal_7865), .Q (signal_7866) ) ;
    buf_clk cell_5336 ( .C (clk), .D (signal_7881), .Q (signal_7882) ) ;
    buf_clk cell_5352 ( .C (clk), .D (signal_7897), .Q (signal_7898) ) ;
    buf_clk cell_5368 ( .C (clk), .D (signal_7913), .Q (signal_7914) ) ;
    buf_clk cell_5384 ( .C (clk), .D (signal_7929), .Q (signal_7930) ) ;
    buf_clk cell_5400 ( .C (clk), .D (signal_7945), .Q (signal_7946) ) ;
    buf_clk cell_5416 ( .C (clk), .D (signal_7961), .Q (signal_7962) ) ;
    buf_clk cell_5432 ( .C (clk), .D (signal_7977), .Q (signal_7978) ) ;
    buf_clk cell_5448 ( .C (clk), .D (signal_7993), .Q (signal_7994) ) ;
    buf_clk cell_5464 ( .C (clk), .D (signal_8009), .Q (signal_8010) ) ;
    buf_clk cell_5480 ( .C (clk), .D (signal_8025), .Q (signal_8026) ) ;
    buf_clk cell_5496 ( .C (clk), .D (signal_8041), .Q (signal_8042) ) ;
    buf_clk cell_5512 ( .C (clk), .D (signal_8057), .Q (signal_8058) ) ;
    buf_clk cell_5528 ( .C (clk), .D (signal_8073), .Q (signal_8074) ) ;
    buf_clk cell_5544 ( .C (clk), .D (signal_8089), .Q (signal_8090) ) ;
    buf_clk cell_5560 ( .C (clk), .D (signal_8105), .Q (signal_8106) ) ;
    buf_clk cell_5576 ( .C (clk), .D (signal_8121), .Q (signal_8122) ) ;
    buf_clk cell_5592 ( .C (clk), .D (signal_8137), .Q (signal_8138) ) ;
    buf_clk cell_5608 ( .C (clk), .D (signal_8153), .Q (signal_8154) ) ;
    buf_clk cell_5624 ( .C (clk), .D (signal_8169), .Q (signal_8170) ) ;
    buf_clk cell_5640 ( .C (clk), .D (signal_8185), .Q (signal_8186) ) ;
    buf_clk cell_5656 ( .C (clk), .D (signal_8201), .Q (signal_8202) ) ;
    buf_clk cell_5672 ( .C (clk), .D (signal_8217), .Q (signal_8218) ) ;
    buf_clk cell_5688 ( .C (clk), .D (signal_8233), .Q (signal_8234) ) ;
    buf_clk cell_5704 ( .C (clk), .D (signal_8249), .Q (signal_8250) ) ;
    buf_clk cell_5720 ( .C (clk), .D (signal_8265), .Q (signal_8266) ) ;
    buf_clk cell_5736 ( .C (clk), .D (signal_8281), .Q (signal_8282) ) ;
    buf_clk cell_5752 ( .C (clk), .D (signal_8297), .Q (signal_8298) ) ;
    buf_clk cell_5768 ( .C (clk), .D (signal_8313), .Q (signal_8314) ) ;
    buf_clk cell_5784 ( .C (clk), .D (signal_8329), .Q (signal_8330) ) ;
    buf_clk cell_5800 ( .C (clk), .D (signal_8345), .Q (signal_8346) ) ;
    buf_clk cell_5816 ( .C (clk), .D (signal_8361), .Q (signal_8362) ) ;
    buf_clk cell_5832 ( .C (clk), .D (signal_8377), .Q (signal_8378) ) ;
    buf_clk cell_5848 ( .C (clk), .D (signal_8393), .Q (signal_8394) ) ;
    buf_clk cell_5864 ( .C (clk), .D (signal_8409), .Q (signal_8410) ) ;
    buf_clk cell_5880 ( .C (clk), .D (signal_8425), .Q (signal_8426) ) ;
    buf_clk cell_5896 ( .C (clk), .D (signal_8441), .Q (signal_8442) ) ;
    buf_clk cell_5912 ( .C (clk), .D (signal_8457), .Q (signal_8458) ) ;
    buf_clk cell_5928 ( .C (clk), .D (signal_8473), .Q (signal_8474) ) ;
    buf_clk cell_5944 ( .C (clk), .D (signal_8489), .Q (signal_8490) ) ;
    buf_clk cell_5960 ( .C (clk), .D (signal_8505), .Q (signal_8506) ) ;
    buf_clk cell_5976 ( .C (clk), .D (signal_8521), .Q (signal_8522) ) ;
    buf_clk cell_5992 ( .C (clk), .D (signal_8537), .Q (signal_8538) ) ;
    buf_clk cell_6008 ( .C (clk), .D (signal_8553), .Q (signal_8554) ) ;
    buf_clk cell_6024 ( .C (clk), .D (signal_8569), .Q (signal_8570) ) ;
    buf_clk cell_6040 ( .C (clk), .D (signal_8585), .Q (signal_8586) ) ;
    buf_clk cell_6056 ( .C (clk), .D (signal_8601), .Q (signal_8602) ) ;
    buf_clk cell_6072 ( .C (clk), .D (signal_8617), .Q (signal_8618) ) ;
    buf_clk cell_6088 ( .C (clk), .D (signal_8633), .Q (signal_8634) ) ;
    buf_clk cell_6104 ( .C (clk), .D (signal_8649), .Q (signal_8650) ) ;
    buf_clk cell_6120 ( .C (clk), .D (signal_8665), .Q (signal_8666) ) ;
    buf_clk cell_6136 ( .C (clk), .D (signal_8681), .Q (signal_8682) ) ;
    buf_clk cell_6152 ( .C (clk), .D (signal_8697), .Q (signal_8698) ) ;
    buf_clk cell_6168 ( .C (clk), .D (signal_8713), .Q (signal_8714) ) ;
    buf_clk cell_6184 ( .C (clk), .D (signal_8729), .Q (signal_8730) ) ;
    buf_clk cell_6200 ( .C (clk), .D (signal_8745), .Q (signal_8746) ) ;
    buf_clk cell_6216 ( .C (clk), .D (signal_8761), .Q (signal_8762) ) ;
    buf_clk cell_6232 ( .C (clk), .D (signal_8777), .Q (signal_8778) ) ;
    buf_clk cell_6248 ( .C (clk), .D (signal_8793), .Q (signal_8794) ) ;
    buf_clk cell_6264 ( .C (clk), .D (signal_8809), .Q (signal_8810) ) ;
    buf_clk cell_6280 ( .C (clk), .D (signal_8825), .Q (signal_8826) ) ;
    buf_clk cell_6296 ( .C (clk), .D (signal_8841), .Q (signal_8842) ) ;
    buf_clk cell_6312 ( .C (clk), .D (signal_8857), .Q (signal_8858) ) ;
    buf_clk cell_6328 ( .C (clk), .D (signal_8873), .Q (signal_8874) ) ;
    buf_clk cell_6344 ( .C (clk), .D (signal_8889), .Q (signal_8890) ) ;
    buf_clk cell_6360 ( .C (clk), .D (signal_8905), .Q (signal_8906) ) ;
    buf_clk cell_6376 ( .C (clk), .D (signal_8921), .Q (signal_8922) ) ;
    buf_clk cell_6392 ( .C (clk), .D (signal_8937), .Q (signal_8938) ) ;
    buf_clk cell_6408 ( .C (clk), .D (signal_8953), .Q (signal_8954) ) ;
    buf_clk cell_6424 ( .C (clk), .D (signal_8969), .Q (signal_8970) ) ;
    buf_clk cell_6440 ( .C (clk), .D (signal_8985), .Q (signal_8986) ) ;
    buf_clk cell_6456 ( .C (clk), .D (signal_9001), .Q (signal_9002) ) ;
    buf_clk cell_6472 ( .C (clk), .D (signal_9017), .Q (signal_9018) ) ;
    buf_clk cell_6488 ( .C (clk), .D (signal_9033), .Q (signal_9034) ) ;
    buf_clk cell_6504 ( .C (clk), .D (signal_9049), .Q (signal_9050) ) ;
    buf_clk cell_6520 ( .C (clk), .D (signal_9065), .Q (signal_9066) ) ;
    buf_clk cell_6536 ( .C (clk), .D (signal_9081), .Q (signal_9082) ) ;
    buf_clk cell_6552 ( .C (clk), .D (signal_9097), .Q (signal_9098) ) ;
    buf_clk cell_6568 ( .C (clk), .D (signal_9113), .Q (signal_9114) ) ;
    buf_clk cell_6584 ( .C (clk), .D (signal_9129), .Q (signal_9130) ) ;
    buf_clk cell_6600 ( .C (clk), .D (signal_9145), .Q (signal_9146) ) ;
    buf_clk cell_6616 ( .C (clk), .D (signal_9161), .Q (signal_9162) ) ;
    buf_clk cell_6632 ( .C (clk), .D (signal_9177), .Q (signal_9178) ) ;
    buf_clk cell_6648 ( .C (clk), .D (signal_9193), .Q (signal_9194) ) ;
    buf_clk cell_6664 ( .C (clk), .D (signal_9209), .Q (signal_9210) ) ;
    buf_clk cell_6680 ( .C (clk), .D (signal_9225), .Q (signal_9226) ) ;
    buf_clk cell_6696 ( .C (clk), .D (signal_9241), .Q (signal_9242) ) ;
    buf_clk cell_6712 ( .C (clk), .D (signal_9257), .Q (signal_9258) ) ;
    buf_clk cell_6728 ( .C (clk), .D (signal_9273), .Q (signal_9274) ) ;
    buf_clk cell_6744 ( .C (clk), .D (signal_9289), .Q (signal_9290) ) ;
    buf_clk cell_6760 ( .C (clk), .D (signal_9305), .Q (signal_9306) ) ;
    buf_clk cell_6776 ( .C (clk), .D (signal_9321), .Q (signal_9322) ) ;
    buf_clk cell_6792 ( .C (clk), .D (signal_9337), .Q (signal_9338) ) ;
    buf_clk cell_6808 ( .C (clk), .D (signal_9353), .Q (signal_9354) ) ;
    buf_clk cell_6824 ( .C (clk), .D (signal_9369), .Q (signal_9370) ) ;
    buf_clk cell_6840 ( .C (clk), .D (signal_9385), .Q (signal_9386) ) ;
    buf_clk cell_6856 ( .C (clk), .D (signal_9401), .Q (signal_9402) ) ;
    buf_clk cell_6872 ( .C (clk), .D (signal_9417), .Q (signal_9418) ) ;
    buf_clk cell_6888 ( .C (clk), .D (signal_9433), .Q (signal_9434) ) ;
    buf_clk cell_6904 ( .C (clk), .D (signal_9449), .Q (signal_9450) ) ;
    buf_clk cell_6920 ( .C (clk), .D (signal_9465), .Q (signal_9466) ) ;
    buf_clk cell_6936 ( .C (clk), .D (signal_9481), .Q (signal_9482) ) ;
    buf_clk cell_6952 ( .C (clk), .D (signal_9497), .Q (signal_9498) ) ;
    buf_clk cell_6968 ( .C (clk), .D (signal_9513), .Q (signal_9514) ) ;
    buf_clk cell_6984 ( .C (clk), .D (signal_9529), .Q (signal_9530) ) ;
    buf_clk cell_7000 ( .C (clk), .D (signal_9545), .Q (signal_9546) ) ;
    buf_clk cell_7016 ( .C (clk), .D (signal_9561), .Q (signal_9562) ) ;
    buf_clk cell_7032 ( .C (clk), .D (signal_9577), .Q (signal_9578) ) ;
    buf_clk cell_7048 ( .C (clk), .D (signal_9593), .Q (signal_9594) ) ;
    buf_clk cell_7064 ( .C (clk), .D (signal_9609), .Q (signal_9610) ) ;
    buf_clk cell_7080 ( .C (clk), .D (signal_9625), .Q (signal_9626) ) ;
    buf_clk cell_7096 ( .C (clk), .D (signal_9641), .Q (signal_9642) ) ;
    buf_clk cell_7112 ( .C (clk), .D (signal_9657), .Q (signal_9658) ) ;
    buf_clk cell_7128 ( .C (clk), .D (signal_9673), .Q (signal_9674) ) ;
    buf_clk cell_7144 ( .C (clk), .D (signal_9689), .Q (signal_9690) ) ;
    buf_clk cell_7160 ( .C (clk), .D (signal_9705), .Q (signal_9706) ) ;
    buf_clk cell_7176 ( .C (clk), .D (signal_9721), .Q (signal_9722) ) ;
    buf_clk cell_7192 ( .C (clk), .D (signal_9737), .Q (signal_9738) ) ;
    buf_clk cell_7208 ( .C (clk), .D (signal_9753), .Q (signal_9754) ) ;
    buf_clk cell_7224 ( .C (clk), .D (signal_9769), .Q (signal_9770) ) ;
    buf_clk cell_7240 ( .C (clk), .D (signal_9785), .Q (signal_9786) ) ;
    buf_clk cell_7256 ( .C (clk), .D (signal_9801), .Q (signal_9802) ) ;
    buf_clk cell_7272 ( .C (clk), .D (signal_9817), .Q (signal_9818) ) ;
    buf_clk cell_7288 ( .C (clk), .D (signal_9833), .Q (signal_9834) ) ;
    buf_clk cell_7304 ( .C (clk), .D (signal_9849), .Q (signal_9850) ) ;
    buf_clk cell_7320 ( .C (clk), .D (signal_9865), .Q (signal_9866) ) ;
    buf_clk cell_7336 ( .C (clk), .D (signal_9881), .Q (signal_9882) ) ;
    buf_clk cell_7352 ( .C (clk), .D (signal_9897), .Q (signal_9898) ) ;
    buf_clk cell_7368 ( .C (clk), .D (signal_9913), .Q (signal_9914) ) ;
    buf_clk cell_7384 ( .C (clk), .D (signal_9929), .Q (signal_9930) ) ;
    buf_clk cell_7400 ( .C (clk), .D (signal_9945), .Q (signal_9946) ) ;
    buf_clk cell_7416 ( .C (clk), .D (signal_9961), .Q (signal_9962) ) ;
    buf_clk cell_7432 ( .C (clk), .D (signal_9977), .Q (signal_9978) ) ;
    buf_clk cell_7448 ( .C (clk), .D (signal_9993), .Q (signal_9994) ) ;
    buf_clk cell_7464 ( .C (clk), .D (signal_10009), .Q (signal_10010) ) ;
    buf_clk cell_7480 ( .C (clk), .D (signal_10025), .Q (signal_10026) ) ;
    buf_clk cell_7496 ( .C (clk), .D (signal_10041), .Q (signal_10042) ) ;
    buf_clk cell_7512 ( .C (clk), .D (signal_10057), .Q (signal_10058) ) ;
    buf_clk cell_7528 ( .C (clk), .D (signal_10073), .Q (signal_10074) ) ;
    buf_clk cell_7544 ( .C (clk), .D (signal_10089), .Q (signal_10090) ) ;
    buf_clk cell_7560 ( .C (clk), .D (signal_10105), .Q (signal_10106) ) ;
    buf_clk cell_7576 ( .C (clk), .D (signal_10121), .Q (signal_10122) ) ;
    buf_clk cell_7592 ( .C (clk), .D (signal_10137), .Q (signal_10138) ) ;
    buf_clk cell_7608 ( .C (clk), .D (signal_10153), .Q (signal_10154) ) ;
    buf_clk cell_7624 ( .C (clk), .D (signal_10169), .Q (signal_10170) ) ;
    buf_clk cell_7640 ( .C (clk), .D (signal_10185), .Q (signal_10186) ) ;
    buf_clk cell_7656 ( .C (clk), .D (signal_10201), .Q (signal_10202) ) ;
    buf_clk cell_7672 ( .C (clk), .D (signal_10217), .Q (signal_10218) ) ;
    buf_clk cell_7688 ( .C (clk), .D (signal_10233), .Q (signal_10234) ) ;
    buf_clk cell_7704 ( .C (clk), .D (signal_10249), .Q (signal_10250) ) ;
    buf_clk cell_7720 ( .C (clk), .D (signal_10265), .Q (signal_10266) ) ;
    buf_clk cell_7736 ( .C (clk), .D (signal_10281), .Q (signal_10282) ) ;
    buf_clk cell_7752 ( .C (clk), .D (signal_10297), .Q (signal_10298) ) ;
    buf_clk cell_7768 ( .C (clk), .D (signal_10313), .Q (signal_10314) ) ;
    buf_clk cell_7784 ( .C (clk), .D (signal_10329), .Q (signal_10330) ) ;
    buf_clk cell_7800 ( .C (clk), .D (signal_10345), .Q (signal_10346) ) ;
    buf_clk cell_7816 ( .C (clk), .D (signal_10361), .Q (signal_10362) ) ;
    buf_clk cell_7832 ( .C (clk), .D (signal_10377), .Q (signal_10378) ) ;
    buf_clk cell_7848 ( .C (clk), .D (signal_10393), .Q (signal_10394) ) ;
    buf_clk cell_7864 ( .C (clk), .D (signal_10409), .Q (signal_10410) ) ;
    buf_clk cell_7880 ( .C (clk), .D (signal_10425), .Q (signal_10426) ) ;
    buf_clk cell_7896 ( .C (clk), .D (signal_10441), .Q (signal_10442) ) ;
    buf_clk cell_7912 ( .C (clk), .D (signal_10457), .Q (signal_10458) ) ;
    buf_clk cell_7928 ( .C (clk), .D (signal_10473), .Q (signal_10474) ) ;
    buf_clk cell_7944 ( .C (clk), .D (signal_10489), .Q (signal_10490) ) ;
    buf_clk cell_7960 ( .C (clk), .D (signal_10505), .Q (signal_10506) ) ;
    buf_clk cell_7976 ( .C (clk), .D (signal_10521), .Q (signal_10522) ) ;
    buf_clk cell_7992 ( .C (clk), .D (signal_10537), .Q (signal_10538) ) ;
    buf_clk cell_8008 ( .C (clk), .D (signal_10553), .Q (signal_10554) ) ;
    buf_clk cell_8024 ( .C (clk), .D (signal_10569), .Q (signal_10570) ) ;
    buf_clk cell_8040 ( .C (clk), .D (signal_10585), .Q (signal_10586) ) ;
    buf_clk cell_8056 ( .C (clk), .D (signal_10601), .Q (signal_10602) ) ;
    buf_clk cell_8072 ( .C (clk), .D (signal_10617), .Q (signal_10618) ) ;
    buf_clk cell_8088 ( .C (clk), .D (signal_10633), .Q (signal_10634) ) ;
    buf_clk cell_8104 ( .C (clk), .D (signal_10649), .Q (signal_10650) ) ;
    buf_clk cell_8120 ( .C (clk), .D (signal_10665), .Q (signal_10666) ) ;
    buf_clk cell_8136 ( .C (clk), .D (signal_10681), .Q (signal_10682) ) ;
    buf_clk cell_8152 ( .C (clk), .D (signal_10697), .Q (signal_10698) ) ;
    buf_clk cell_8168 ( .C (clk), .D (signal_10713), .Q (signal_10714) ) ;
    buf_clk cell_8184 ( .C (clk), .D (signal_10729), .Q (signal_10730) ) ;
    buf_clk cell_8200 ( .C (clk), .D (signal_10745), .Q (signal_10746) ) ;
    buf_clk cell_8216 ( .C (clk), .D (signal_10761), .Q (signal_10762) ) ;
    buf_clk cell_8232 ( .C (clk), .D (signal_10777), .Q (signal_10778) ) ;
    buf_clk cell_8248 ( .C (clk), .D (signal_10793), .Q (signal_10794) ) ;
    buf_clk cell_8264 ( .C (clk), .D (signal_10809), .Q (signal_10810) ) ;
    buf_clk cell_8280 ( .C (clk), .D (signal_10825), .Q (signal_10826) ) ;
    buf_clk cell_8296 ( .C (clk), .D (signal_10841), .Q (signal_10842) ) ;
    buf_clk cell_8312 ( .C (clk), .D (signal_10857), .Q (signal_10858) ) ;
    buf_clk cell_8328 ( .C (clk), .D (signal_10873), .Q (signal_10874) ) ;
    buf_clk cell_8344 ( .C (clk), .D (signal_10889), .Q (signal_10890) ) ;
    buf_clk cell_8360 ( .C (clk), .D (signal_10905), .Q (signal_10906) ) ;
    buf_clk cell_8376 ( .C (clk), .D (signal_10921), .Q (signal_10922) ) ;
    buf_clk cell_8392 ( .C (clk), .D (signal_10937), .Q (signal_10938) ) ;
    buf_clk cell_8408 ( .C (clk), .D (signal_10953), .Q (signal_10954) ) ;
    buf_clk cell_8424 ( .C (clk), .D (signal_10969), .Q (signal_10970) ) ;
    buf_clk cell_8440 ( .C (clk), .D (signal_10985), .Q (signal_10986) ) ;
    buf_clk cell_8456 ( .C (clk), .D (signal_11001), .Q (signal_11002) ) ;
    buf_clk cell_8472 ( .C (clk), .D (signal_11017), .Q (signal_11018) ) ;
    buf_clk cell_8488 ( .C (clk), .D (signal_11033), .Q (signal_11034) ) ;
    buf_clk cell_8504 ( .C (clk), .D (signal_11049), .Q (signal_11050) ) ;
    buf_clk cell_8520 ( .C (clk), .D (signal_11065), .Q (signal_11066) ) ;
    buf_clk cell_8536 ( .C (clk), .D (signal_11081), .Q (signal_11082) ) ;
    buf_clk cell_8552 ( .C (clk), .D (signal_11097), .Q (signal_11098) ) ;
    buf_clk cell_8568 ( .C (clk), .D (signal_11113), .Q (signal_11114) ) ;
    buf_clk cell_8584 ( .C (clk), .D (signal_11129), .Q (signal_11130) ) ;
    buf_clk cell_8600 ( .C (clk), .D (signal_11145), .Q (signal_11146) ) ;
    buf_clk cell_8616 ( .C (clk), .D (signal_11161), .Q (signal_11162) ) ;
    buf_clk cell_8632 ( .C (clk), .D (signal_11177), .Q (signal_11178) ) ;
    buf_clk cell_8648 ( .C (clk), .D (signal_11193), .Q (signal_11194) ) ;
    buf_clk cell_8664 ( .C (clk), .D (signal_11209), .Q (signal_11210) ) ;
    buf_clk cell_8680 ( .C (clk), .D (signal_11225), .Q (signal_11226) ) ;
    buf_clk cell_8696 ( .C (clk), .D (signal_11241), .Q (signal_11242) ) ;
    buf_clk cell_8712 ( .C (clk), .D (signal_11257), .Q (signal_11258) ) ;
    buf_clk cell_8728 ( .C (clk), .D (signal_11273), .Q (signal_11274) ) ;
    buf_clk cell_8744 ( .C (clk), .D (signal_11289), .Q (signal_11290) ) ;
    buf_clk cell_8760 ( .C (clk), .D (signal_11305), .Q (signal_11306) ) ;
    buf_clk cell_8776 ( .C (clk), .D (signal_11321), .Q (signal_11322) ) ;
    buf_clk cell_8792 ( .C (clk), .D (signal_11337), .Q (signal_11338) ) ;
    buf_clk cell_8808 ( .C (clk), .D (signal_11353), .Q (signal_11354) ) ;
    buf_clk cell_8824 ( .C (clk), .D (signal_11369), .Q (signal_11370) ) ;
    buf_clk cell_8840 ( .C (clk), .D (signal_11385), .Q (signal_11386) ) ;
    buf_clk cell_8856 ( .C (clk), .D (signal_11401), .Q (signal_11402) ) ;
    buf_clk cell_8872 ( .C (clk), .D (signal_11417), .Q (signal_11418) ) ;
    buf_clk cell_8888 ( .C (clk), .D (signal_11433), .Q (signal_11434) ) ;
    buf_clk cell_8904 ( .C (clk), .D (signal_11449), .Q (signal_11450) ) ;
    buf_clk cell_8920 ( .C (clk), .D (signal_11465), .Q (signal_11466) ) ;
    buf_clk cell_8936 ( .C (clk), .D (signal_11481), .Q (signal_11482) ) ;
    buf_clk cell_8952 ( .C (clk), .D (signal_11497), .Q (signal_11498) ) ;
    buf_clk cell_8968 ( .C (clk), .D (signal_11513), .Q (signal_11514) ) ;
    buf_clk cell_8984 ( .C (clk), .D (signal_11529), .Q (signal_11530) ) ;
    buf_clk cell_9000 ( .C (clk), .D (signal_11545), .Q (signal_11546) ) ;
    buf_clk cell_9016 ( .C (clk), .D (signal_11561), .Q (signal_11562) ) ;
    buf_clk cell_9032 ( .C (clk), .D (signal_11577), .Q (signal_11578) ) ;
    buf_clk cell_9048 ( .C (clk), .D (signal_11593), .Q (signal_11594) ) ;
    buf_clk cell_9064 ( .C (clk), .D (signal_11609), .Q (signal_11610) ) ;
    buf_clk cell_9080 ( .C (clk), .D (signal_11625), .Q (signal_11626) ) ;
    buf_clk cell_9096 ( .C (clk), .D (signal_11641), .Q (signal_11642) ) ;
    buf_clk cell_9112 ( .C (clk), .D (signal_11657), .Q (signal_11658) ) ;
    buf_clk cell_9128 ( .C (clk), .D (signal_11673), .Q (signal_11674) ) ;
    buf_clk cell_9144 ( .C (clk), .D (signal_11689), .Q (signal_11690) ) ;
    buf_clk cell_9160 ( .C (clk), .D (signal_11705), .Q (signal_11706) ) ;
    buf_clk cell_9176 ( .C (clk), .D (signal_11721), .Q (signal_11722) ) ;
    buf_clk cell_9192 ( .C (clk), .D (signal_11737), .Q (signal_11738) ) ;
    buf_clk cell_9208 ( .C (clk), .D (signal_11753), .Q (signal_11754) ) ;
    buf_clk cell_9224 ( .C (clk), .D (signal_11769), .Q (signal_11770) ) ;
    buf_clk cell_9240 ( .C (clk), .D (signal_11785), .Q (signal_11786) ) ;
    buf_clk cell_9256 ( .C (clk), .D (signal_11801), .Q (signal_11802) ) ;
    buf_clk cell_9272 ( .C (clk), .D (signal_11817), .Q (signal_11818) ) ;
    buf_clk cell_9288 ( .C (clk), .D (signal_11833), .Q (signal_11834) ) ;
    buf_clk cell_9304 ( .C (clk), .D (signal_11849), .Q (signal_11850) ) ;
    buf_clk cell_9320 ( .C (clk), .D (signal_11865), .Q (signal_11866) ) ;
    buf_clk cell_9336 ( .C (clk), .D (signal_11881), .Q (signal_11882) ) ;
    buf_clk cell_9352 ( .C (clk), .D (signal_11897), .Q (signal_11898) ) ;
    buf_clk cell_9368 ( .C (clk), .D (signal_11913), .Q (signal_11914) ) ;
    buf_clk cell_9384 ( .C (clk), .D (signal_11929), .Q (signal_11930) ) ;
    buf_clk cell_9400 ( .C (clk), .D (signal_11945), .Q (signal_11946) ) ;
    buf_clk cell_9416 ( .C (clk), .D (signal_11961), .Q (signal_11962) ) ;
    buf_clk cell_9432 ( .C (clk), .D (signal_11977), .Q (signal_11978) ) ;
    buf_clk cell_9448 ( .C (clk), .D (signal_11993), .Q (signal_11994) ) ;
    buf_clk cell_9464 ( .C (clk), .D (signal_12009), .Q (signal_12010) ) ;
    buf_clk cell_9480 ( .C (clk), .D (signal_12025), .Q (signal_12026) ) ;
    buf_clk cell_9496 ( .C (clk), .D (signal_12041), .Q (signal_12042) ) ;
    buf_clk cell_9512 ( .C (clk), .D (signal_12057), .Q (signal_12058) ) ;
    buf_clk cell_9528 ( .C (clk), .D (signal_12073), .Q (signal_12074) ) ;
    buf_clk cell_9544 ( .C (clk), .D (signal_12089), .Q (signal_12090) ) ;
    buf_clk cell_9560 ( .C (clk), .D (signal_12105), .Q (signal_12106) ) ;
    buf_clk cell_9576 ( .C (clk), .D (signal_12121), .Q (signal_12122) ) ;
    buf_clk cell_9592 ( .C (clk), .D (signal_12137), .Q (signal_12138) ) ;
    buf_clk cell_9608 ( .C (clk), .D (signal_12153), .Q (signal_12154) ) ;
    buf_clk cell_9624 ( .C (clk), .D (signal_12169), .Q (signal_12170) ) ;
    buf_clk cell_9640 ( .C (clk), .D (signal_12185), .Q (signal_12186) ) ;
    buf_clk cell_9656 ( .C (clk), .D (signal_12201), .Q (signal_12202) ) ;
    buf_clk cell_9672 ( .C (clk), .D (signal_12217), .Q (signal_12218) ) ;
    buf_clk cell_9688 ( .C (clk), .D (signal_12233), .Q (signal_12234) ) ;
    buf_clk cell_9704 ( .C (clk), .D (signal_12249), .Q (signal_12250) ) ;
    buf_clk cell_9720 ( .C (clk), .D (signal_12265), .Q (signal_12266) ) ;
    buf_clk cell_9736 ( .C (clk), .D (signal_12281), .Q (signal_12282) ) ;
    buf_clk cell_9752 ( .C (clk), .D (signal_12297), .Q (signal_12298) ) ;
    buf_clk cell_9768 ( .C (clk), .D (signal_12313), .Q (signal_12314) ) ;
    buf_clk cell_9784 ( .C (clk), .D (signal_12329), .Q (signal_12330) ) ;
    buf_clk cell_9800 ( .C (clk), .D (signal_12345), .Q (signal_12346) ) ;
    buf_clk cell_9816 ( .C (clk), .D (signal_12361), .Q (signal_12362) ) ;
    buf_clk cell_9832 ( .C (clk), .D (signal_12377), .Q (signal_12378) ) ;
    buf_clk cell_9848 ( .C (clk), .D (signal_12393), .Q (signal_12394) ) ;
    buf_clk cell_9864 ( .C (clk), .D (signal_12409), .Q (signal_12410) ) ;
    buf_clk cell_9880 ( .C (clk), .D (signal_12425), .Q (signal_12426) ) ;
    buf_clk cell_9896 ( .C (clk), .D (signal_12441), .Q (signal_12442) ) ;
    buf_clk cell_9912 ( .C (clk), .D (signal_12457), .Q (signal_12458) ) ;
    buf_clk cell_9928 ( .C (clk), .D (signal_12473), .Q (signal_12474) ) ;
    buf_clk cell_9944 ( .C (clk), .D (signal_12489), .Q (signal_12490) ) ;
    buf_clk cell_9960 ( .C (clk), .D (signal_12505), .Q (signal_12506) ) ;
    buf_clk cell_9976 ( .C (clk), .D (signal_12521), .Q (signal_12522) ) ;
    buf_clk cell_9992 ( .C (clk), .D (signal_12537), .Q (signal_12538) ) ;
    buf_clk cell_10008 ( .C (clk), .D (signal_12553), .Q (signal_12554) ) ;
    buf_clk cell_10024 ( .C (clk), .D (signal_12569), .Q (signal_12570) ) ;
    buf_clk cell_10040 ( .C (clk), .D (signal_12585), .Q (signal_12586) ) ;
    buf_clk cell_10056 ( .C (clk), .D (signal_12601), .Q (signal_12602) ) ;
    buf_clk cell_10072 ( .C (clk), .D (signal_12617), .Q (signal_12618) ) ;
    buf_clk cell_10088 ( .C (clk), .D (signal_12633), .Q (signal_12634) ) ;
    buf_clk cell_10104 ( .C (clk), .D (signal_12649), .Q (signal_12650) ) ;
    buf_clk cell_10120 ( .C (clk), .D (signal_12665), .Q (signal_12666) ) ;
    buf_clk cell_10136 ( .C (clk), .D (signal_12681), .Q (signal_12682) ) ;
    buf_clk cell_10152 ( .C (clk), .D (signal_12697), .Q (signal_12698) ) ;
    buf_clk cell_10168 ( .C (clk), .D (signal_12713), .Q (signal_12714) ) ;
    buf_clk cell_10184 ( .C (clk), .D (signal_12729), .Q (signal_12730) ) ;
    buf_clk cell_10200 ( .C (clk), .D (signal_12745), .Q (signal_12746) ) ;
    buf_clk cell_10216 ( .C (clk), .D (signal_12761), .Q (signal_12762) ) ;
    buf_clk cell_10232 ( .C (clk), .D (signal_12777), .Q (signal_12778) ) ;
    buf_clk cell_10248 ( .C (clk), .D (signal_12793), .Q (signal_12794) ) ;
    buf_clk cell_10264 ( .C (clk), .D (signal_12809), .Q (signal_12810) ) ;
    buf_clk cell_10280 ( .C (clk), .D (signal_12825), .Q (signal_12826) ) ;
    buf_clk cell_10296 ( .C (clk), .D (signal_12841), .Q (signal_12842) ) ;
    buf_clk cell_10312 ( .C (clk), .D (signal_12857), .Q (signal_12858) ) ;
    buf_clk cell_10328 ( .C (clk), .D (signal_12873), .Q (signal_12874) ) ;
    buf_clk cell_10344 ( .C (clk), .D (signal_12889), .Q (signal_12890) ) ;
    buf_clk cell_10360 ( .C (clk), .D (signal_12905), .Q (signal_12906) ) ;
    buf_clk cell_10376 ( .C (clk), .D (signal_12921), .Q (signal_12922) ) ;
    buf_clk cell_10392 ( .C (clk), .D (signal_12937), .Q (signal_12938) ) ;
    buf_clk cell_10408 ( .C (clk), .D (signal_12953), .Q (signal_12954) ) ;
    buf_clk cell_10424 ( .C (clk), .D (signal_12969), .Q (signal_12970) ) ;
    buf_clk cell_10440 ( .C (clk), .D (signal_12985), .Q (signal_12986) ) ;
    buf_clk cell_10456 ( .C (clk), .D (signal_13001), .Q (signal_13002) ) ;
    buf_clk cell_10472 ( .C (clk), .D (signal_13017), .Q (signal_13018) ) ;
    buf_clk cell_10488 ( .C (clk), .D (signal_13033), .Q (signal_13034) ) ;
    buf_clk cell_10504 ( .C (clk), .D (signal_13049), .Q (signal_13050) ) ;
    buf_clk cell_10520 ( .C (clk), .D (signal_13065), .Q (signal_13066) ) ;
    buf_clk cell_10536 ( .C (clk), .D (signal_13081), .Q (signal_13082) ) ;
    buf_clk cell_10552 ( .C (clk), .D (signal_13097), .Q (signal_13098) ) ;
    buf_clk cell_10568 ( .C (clk), .D (signal_13113), .Q (signal_13114) ) ;
    buf_clk cell_10584 ( .C (clk), .D (signal_13129), .Q (signal_13130) ) ;
    buf_clk cell_10600 ( .C (clk), .D (signal_13145), .Q (signal_13146) ) ;
    buf_clk cell_10616 ( .C (clk), .D (signal_13161), .Q (signal_13162) ) ;
    buf_clk cell_10632 ( .C (clk), .D (signal_13177), .Q (signal_13178) ) ;
    buf_clk cell_10648 ( .C (clk), .D (signal_13193), .Q (signal_13194) ) ;
    buf_clk cell_10664 ( .C (clk), .D (signal_13209), .Q (signal_13210) ) ;
    buf_clk cell_10680 ( .C (clk), .D (signal_13225), .Q (signal_13226) ) ;
    buf_clk cell_10696 ( .C (clk), .D (signal_13241), .Q (signal_13242) ) ;
    buf_clk cell_10712 ( .C (clk), .D (signal_13257), .Q (signal_13258) ) ;
    buf_clk cell_10728 ( .C (clk), .D (signal_13273), .Q (signal_13274) ) ;
    buf_clk cell_10744 ( .C (clk), .D (signal_13289), .Q (signal_13290) ) ;
    buf_clk cell_10760 ( .C (clk), .D (signal_13305), .Q (signal_13306) ) ;
    buf_clk cell_10776 ( .C (clk), .D (signal_13321), .Q (signal_13322) ) ;
    buf_clk cell_10792 ( .C (clk), .D (signal_13337), .Q (signal_13338) ) ;
    buf_clk cell_10808 ( .C (clk), .D (signal_13353), .Q (signal_13354) ) ;
    buf_clk cell_10824 ( .C (clk), .D (signal_13369), .Q (signal_13370) ) ;
    buf_clk cell_10840 ( .C (clk), .D (signal_13385), .Q (signal_13386) ) ;
    buf_clk cell_10856 ( .C (clk), .D (signal_13401), .Q (signal_13402) ) ;
    buf_clk cell_10872 ( .C (clk), .D (signal_13417), .Q (signal_13418) ) ;
    buf_clk cell_10888 ( .C (clk), .D (signal_13433), .Q (signal_13434) ) ;
    buf_clk cell_10904 ( .C (clk), .D (signal_13449), .Q (signal_13450) ) ;
    buf_clk cell_10920 ( .C (clk), .D (signal_13465), .Q (signal_13466) ) ;
    buf_clk cell_10936 ( .C (clk), .D (signal_13481), .Q (signal_13482) ) ;
    buf_clk cell_10952 ( .C (clk), .D (signal_13497), .Q (signal_13498) ) ;
    buf_clk cell_10968 ( .C (clk), .D (signal_13513), .Q (signal_13514) ) ;
    buf_clk cell_10984 ( .C (clk), .D (signal_13529), .Q (signal_13530) ) ;
    buf_clk cell_11000 ( .C (clk), .D (signal_13545), .Q (signal_13546) ) ;
    buf_clk cell_11016 ( .C (clk), .D (signal_13561), .Q (signal_13562) ) ;
    buf_clk cell_11032 ( .C (clk), .D (signal_13577), .Q (signal_13578) ) ;
    buf_clk cell_11048 ( .C (clk), .D (signal_13593), .Q (signal_13594) ) ;
    buf_clk cell_11064 ( .C (clk), .D (signal_13609), .Q (signal_13610) ) ;
    buf_clk cell_11080 ( .C (clk), .D (signal_13625), .Q (signal_13626) ) ;
    buf_clk cell_11096 ( .C (clk), .D (signal_13641), .Q (signal_13642) ) ;
    buf_clk cell_11112 ( .C (clk), .D (signal_13657), .Q (signal_13658) ) ;
    buf_clk cell_11128 ( .C (clk), .D (signal_13673), .Q (signal_13674) ) ;
    buf_clk cell_11144 ( .C (clk), .D (signal_13689), .Q (signal_13690) ) ;
    buf_clk cell_11160 ( .C (clk), .D (signal_13705), .Q (signal_13706) ) ;
    buf_clk cell_11176 ( .C (clk), .D (signal_13721), .Q (signal_13722) ) ;
    buf_clk cell_11192 ( .C (clk), .D (signal_13737), .Q (signal_13738) ) ;
    buf_clk cell_11208 ( .C (clk), .D (signal_13753), .Q (signal_13754) ) ;
    buf_clk cell_11224 ( .C (clk), .D (signal_13769), .Q (signal_13770) ) ;
    buf_clk cell_11240 ( .C (clk), .D (signal_13785), .Q (signal_13786) ) ;
    buf_clk cell_11256 ( .C (clk), .D (signal_13801), .Q (signal_13802) ) ;
    buf_clk cell_11272 ( .C (clk), .D (signal_13817), .Q (signal_13818) ) ;
    buf_clk cell_11288 ( .C (clk), .D (signal_13833), .Q (signal_13834) ) ;
    buf_clk cell_11304 ( .C (clk), .D (signal_13849), .Q (signal_13850) ) ;
    buf_clk cell_11320 ( .C (clk), .D (signal_13865), .Q (signal_13866) ) ;
    buf_clk cell_11336 ( .C (clk), .D (signal_13881), .Q (signal_13882) ) ;
    buf_clk cell_11352 ( .C (clk), .D (signal_13897), .Q (signal_13898) ) ;
    buf_clk cell_11368 ( .C (clk), .D (signal_13913), .Q (signal_13914) ) ;
    buf_clk cell_11384 ( .C (clk), .D (signal_13929), .Q (signal_13930) ) ;
    buf_clk cell_11400 ( .C (clk), .D (signal_13945), .Q (signal_13946) ) ;
    buf_clk cell_11416 ( .C (clk), .D (signal_13961), .Q (signal_13962) ) ;
    buf_clk cell_11432 ( .C (clk), .D (signal_13977), .Q (signal_13978) ) ;
    buf_clk cell_11448 ( .C (clk), .D (signal_13993), .Q (signal_13994) ) ;
    buf_clk cell_11464 ( .C (clk), .D (signal_14009), .Q (signal_14010) ) ;
    buf_clk cell_11480 ( .C (clk), .D (signal_14025), .Q (signal_14026) ) ;
    buf_clk cell_11496 ( .C (clk), .D (signal_14041), .Q (signal_14042) ) ;
    buf_clk cell_11512 ( .C (clk), .D (signal_14057), .Q (signal_14058) ) ;
    buf_clk cell_11528 ( .C (clk), .D (signal_14073), .Q (signal_14074) ) ;
    buf_clk cell_11544 ( .C (clk), .D (signal_14089), .Q (signal_14090) ) ;
    buf_clk cell_11560 ( .C (clk), .D (signal_14105), .Q (signal_14106) ) ;
    buf_clk cell_11576 ( .C (clk), .D (signal_14121), .Q (signal_14122) ) ;
    buf_clk cell_11592 ( .C (clk), .D (signal_14137), .Q (signal_14138) ) ;
    buf_clk cell_11608 ( .C (clk), .D (signal_14153), .Q (signal_14154) ) ;
    buf_clk cell_11624 ( .C (clk), .D (signal_14169), .Q (signal_14170) ) ;
    buf_clk cell_11640 ( .C (clk), .D (signal_14185), .Q (signal_14186) ) ;
    buf_clk cell_11656 ( .C (clk), .D (signal_14201), .Q (signal_14202) ) ;
    buf_clk cell_11672 ( .C (clk), .D (signal_14217), .Q (signal_14218) ) ;
    buf_clk cell_11688 ( .C (clk), .D (signal_14233), .Q (signal_14234) ) ;
    buf_clk cell_11704 ( .C (clk), .D (signal_14249), .Q (signal_14250) ) ;
    buf_clk cell_11720 ( .C (clk), .D (signal_14265), .Q (signal_14266) ) ;
    buf_clk cell_11736 ( .C (clk), .D (signal_14281), .Q (signal_14282) ) ;
    buf_clk cell_11752 ( .C (clk), .D (signal_14297), .Q (signal_14298) ) ;
    buf_clk cell_11768 ( .C (clk), .D (signal_14313), .Q (signal_14314) ) ;
    buf_clk cell_11784 ( .C (clk), .D (signal_14329), .Q (signal_14330) ) ;
    buf_clk cell_11800 ( .C (clk), .D (signal_14345), .Q (signal_14346) ) ;
    buf_clk cell_11816 ( .C (clk), .D (signal_14361), .Q (signal_14362) ) ;
    buf_clk cell_11832 ( .C (clk), .D (signal_14377), .Q (signal_14378) ) ;
    buf_clk cell_11848 ( .C (clk), .D (signal_14393), .Q (signal_14394) ) ;
    buf_clk cell_11864 ( .C (clk), .D (signal_14409), .Q (signal_14410) ) ;
    buf_clk cell_11880 ( .C (clk), .D (signal_14425), .Q (signal_14426) ) ;
    buf_clk cell_11896 ( .C (clk), .D (signal_14441), .Q (signal_14442) ) ;
    buf_clk cell_11912 ( .C (clk), .D (signal_14457), .Q (signal_14458) ) ;
    buf_clk cell_11928 ( .C (clk), .D (signal_14473), .Q (signal_14474) ) ;
    buf_clk cell_11944 ( .C (clk), .D (signal_14489), .Q (signal_14490) ) ;
    buf_clk cell_11960 ( .C (clk), .D (signal_14505), .Q (signal_14506) ) ;
    buf_clk cell_11976 ( .C (clk), .D (signal_14521), .Q (signal_14522) ) ;
    buf_clk cell_11992 ( .C (clk), .D (signal_14537), .Q (signal_14538) ) ;
    buf_clk cell_12008 ( .C (clk), .D (signal_14553), .Q (signal_14554) ) ;
    buf_clk cell_12024 ( .C (clk), .D (signal_14569), .Q (signal_14570) ) ;
    buf_clk cell_12040 ( .C (clk), .D (signal_14585), .Q (signal_14586) ) ;
    buf_clk cell_12056 ( .C (clk), .D (signal_14601), .Q (signal_14602) ) ;
    buf_clk cell_12072 ( .C (clk), .D (signal_14617), .Q (signal_14618) ) ;
    buf_clk cell_12088 ( .C (clk), .D (signal_14633), .Q (signal_14634) ) ;
    buf_clk cell_12104 ( .C (clk), .D (signal_14649), .Q (signal_14650) ) ;
    buf_clk cell_12120 ( .C (clk), .D (signal_14665), .Q (signal_14666) ) ;
    buf_clk cell_12136 ( .C (clk), .D (signal_14681), .Q (signal_14682) ) ;
    buf_clk cell_12152 ( .C (clk), .D (signal_14697), .Q (signal_14698) ) ;
    buf_clk cell_12168 ( .C (clk), .D (signal_14713), .Q (signal_14714) ) ;
    buf_clk cell_12184 ( .C (clk), .D (signal_14729), .Q (signal_14730) ) ;
    buf_clk cell_12200 ( .C (clk), .D (signal_14745), .Q (signal_14746) ) ;
    buf_clk cell_12216 ( .C (clk), .D (signal_14761), .Q (signal_14762) ) ;
    buf_clk cell_12232 ( .C (clk), .D (signal_14777), .Q (signal_14778) ) ;
    buf_clk cell_12248 ( .C (clk), .D (signal_14793), .Q (signal_14794) ) ;
    buf_clk cell_12264 ( .C (clk), .D (signal_14809), .Q (signal_14810) ) ;
    buf_clk cell_12280 ( .C (clk), .D (signal_14825), .Q (signal_14826) ) ;
    buf_clk cell_12296 ( .C (clk), .D (signal_14841), .Q (signal_14842) ) ;
    buf_clk cell_12312 ( .C (clk), .D (signal_14857), .Q (signal_14858) ) ;
    buf_clk cell_12328 ( .C (clk), .D (signal_14873), .Q (signal_14874) ) ;
    buf_clk cell_12344 ( .C (clk), .D (signal_14889), .Q (signal_14890) ) ;
    buf_clk cell_12360 ( .C (clk), .D (signal_14905), .Q (signal_14906) ) ;
    buf_clk cell_12376 ( .C (clk), .D (signal_14921), .Q (signal_14922) ) ;
    buf_clk cell_12392 ( .C (clk), .D (signal_14937), .Q (signal_14938) ) ;

    /* cells in depth 13 */
    buf_clk cell_2397 ( .C (clk), .D (signal_4942), .Q (signal_4943) ) ;
    buf_clk cell_2413 ( .C (clk), .D (signal_4958), .Q (signal_4959) ) ;
    buf_clk cell_2429 ( .C (clk), .D (signal_4974), .Q (signal_4975) ) ;
    buf_clk cell_2445 ( .C (clk), .D (signal_4990), .Q (signal_4991) ) ;
    buf_clk cell_2461 ( .C (clk), .D (signal_5006), .Q (signal_5007) ) ;
    buf_clk cell_2477 ( .C (clk), .D (signal_5022), .Q (signal_5023) ) ;
    buf_clk cell_2493 ( .C (clk), .D (signal_5038), .Q (signal_5039) ) ;
    buf_clk cell_2509 ( .C (clk), .D (signal_5054), .Q (signal_5055) ) ;
    buf_clk cell_2525 ( .C (clk), .D (signal_5070), .Q (signal_5071) ) ;
    buf_clk cell_2541 ( .C (clk), .D (signal_5086), .Q (signal_5087) ) ;
    buf_clk cell_2557 ( .C (clk), .D (signal_5102), .Q (signal_5103) ) ;
    buf_clk cell_2573 ( .C (clk), .D (signal_5118), .Q (signal_5119) ) ;
    buf_clk cell_2589 ( .C (clk), .D (signal_5134), .Q (signal_5135) ) ;
    buf_clk cell_2605 ( .C (clk), .D (signal_5150), .Q (signal_5151) ) ;
    buf_clk cell_2621 ( .C (clk), .D (signal_5166), .Q (signal_5167) ) ;
    buf_clk cell_2637 ( .C (clk), .D (signal_5182), .Q (signal_5183) ) ;
    buf_clk cell_2653 ( .C (clk), .D (signal_5198), .Q (signal_5199) ) ;
    buf_clk cell_2669 ( .C (clk), .D (signal_5214), .Q (signal_5215) ) ;
    buf_clk cell_2685 ( .C (clk), .D (signal_5230), .Q (signal_5231) ) ;
    buf_clk cell_2701 ( .C (clk), .D (signal_5246), .Q (signal_5247) ) ;
    buf_clk cell_2717 ( .C (clk), .D (signal_5262), .Q (signal_5263) ) ;
    buf_clk cell_2733 ( .C (clk), .D (signal_5278), .Q (signal_5279) ) ;
    buf_clk cell_2749 ( .C (clk), .D (signal_5294), .Q (signal_5295) ) ;
    buf_clk cell_2765 ( .C (clk), .D (signal_5310), .Q (signal_5311) ) ;
    buf_clk cell_2781 ( .C (clk), .D (signal_5326), .Q (signal_5327) ) ;
    buf_clk cell_2797 ( .C (clk), .D (signal_5342), .Q (signal_5343) ) ;
    buf_clk cell_2813 ( .C (clk), .D (signal_5358), .Q (signal_5359) ) ;
    buf_clk cell_2829 ( .C (clk), .D (signal_5374), .Q (signal_5375) ) ;
    buf_clk cell_2845 ( .C (clk), .D (signal_5390), .Q (signal_5391) ) ;
    buf_clk cell_2861 ( .C (clk), .D (signal_5406), .Q (signal_5407) ) ;
    buf_clk cell_2877 ( .C (clk), .D (signal_5422), .Q (signal_5423) ) ;
    buf_clk cell_2893 ( .C (clk), .D (signal_5438), .Q (signal_5439) ) ;
    buf_clk cell_2909 ( .C (clk), .D (signal_5454), .Q (signal_5455) ) ;
    buf_clk cell_2925 ( .C (clk), .D (signal_5470), .Q (signal_5471) ) ;
    buf_clk cell_2941 ( .C (clk), .D (signal_5486), .Q (signal_5487) ) ;
    buf_clk cell_2957 ( .C (clk), .D (signal_5502), .Q (signal_5503) ) ;
    buf_clk cell_2973 ( .C (clk), .D (signal_5518), .Q (signal_5519) ) ;
    buf_clk cell_2989 ( .C (clk), .D (signal_5534), .Q (signal_5535) ) ;
    buf_clk cell_3005 ( .C (clk), .D (signal_5550), .Q (signal_5551) ) ;
    buf_clk cell_3021 ( .C (clk), .D (signal_5566), .Q (signal_5567) ) ;
    buf_clk cell_3037 ( .C (clk), .D (signal_5582), .Q (signal_5583) ) ;
    buf_clk cell_3053 ( .C (clk), .D (signal_5598), .Q (signal_5599) ) ;
    buf_clk cell_3069 ( .C (clk), .D (signal_5614), .Q (signal_5615) ) ;
    buf_clk cell_3085 ( .C (clk), .D (signal_5630), .Q (signal_5631) ) ;
    buf_clk cell_3101 ( .C (clk), .D (signal_5646), .Q (signal_5647) ) ;
    buf_clk cell_3117 ( .C (clk), .D (signal_5662), .Q (signal_5663) ) ;
    buf_clk cell_3133 ( .C (clk), .D (signal_5678), .Q (signal_5679) ) ;
    buf_clk cell_3149 ( .C (clk), .D (signal_5694), .Q (signal_5695) ) ;
    buf_clk cell_3165 ( .C (clk), .D (signal_5710), .Q (signal_5711) ) ;
    buf_clk cell_3181 ( .C (clk), .D (signal_5726), .Q (signal_5727) ) ;
    buf_clk cell_3197 ( .C (clk), .D (signal_5742), .Q (signal_5743) ) ;
    buf_clk cell_3213 ( .C (clk), .D (signal_5758), .Q (signal_5759) ) ;
    buf_clk cell_3229 ( .C (clk), .D (signal_5774), .Q (signal_5775) ) ;
    buf_clk cell_3245 ( .C (clk), .D (signal_5790), .Q (signal_5791) ) ;
    buf_clk cell_3261 ( .C (clk), .D (signal_5806), .Q (signal_5807) ) ;
    buf_clk cell_3277 ( .C (clk), .D (signal_5822), .Q (signal_5823) ) ;
    buf_clk cell_3293 ( .C (clk), .D (signal_5838), .Q (signal_5839) ) ;
    buf_clk cell_3309 ( .C (clk), .D (signal_5854), .Q (signal_5855) ) ;
    buf_clk cell_3325 ( .C (clk), .D (signal_5870), .Q (signal_5871) ) ;
    buf_clk cell_3341 ( .C (clk), .D (signal_5886), .Q (signal_5887) ) ;
    buf_clk cell_3357 ( .C (clk), .D (signal_5902), .Q (signal_5903) ) ;
    buf_clk cell_3373 ( .C (clk), .D (signal_5918), .Q (signal_5919) ) ;
    buf_clk cell_3389 ( .C (clk), .D (signal_5934), .Q (signal_5935) ) ;
    buf_clk cell_3405 ( .C (clk), .D (signal_5950), .Q (signal_5951) ) ;
    buf_clk cell_3421 ( .C (clk), .D (signal_5966), .Q (signal_5967) ) ;
    buf_clk cell_3437 ( .C (clk), .D (signal_5982), .Q (signal_5983) ) ;
    buf_clk cell_3453 ( .C (clk), .D (signal_5998), .Q (signal_5999) ) ;
    buf_clk cell_3469 ( .C (clk), .D (signal_6014), .Q (signal_6015) ) ;
    buf_clk cell_3485 ( .C (clk), .D (signal_6030), .Q (signal_6031) ) ;
    buf_clk cell_3501 ( .C (clk), .D (signal_6046), .Q (signal_6047) ) ;
    buf_clk cell_3517 ( .C (clk), .D (signal_6062), .Q (signal_6063) ) ;
    buf_clk cell_3533 ( .C (clk), .D (signal_6078), .Q (signal_6079) ) ;
    buf_clk cell_3549 ( .C (clk), .D (signal_6094), .Q (signal_6095) ) ;
    buf_clk cell_3565 ( .C (clk), .D (signal_6110), .Q (signal_6111) ) ;
    buf_clk cell_3581 ( .C (clk), .D (signal_6126), .Q (signal_6127) ) ;
    buf_clk cell_3597 ( .C (clk), .D (signal_6142), .Q (signal_6143) ) ;
    buf_clk cell_3613 ( .C (clk), .D (signal_6158), .Q (signal_6159) ) ;
    buf_clk cell_3629 ( .C (clk), .D (signal_6174), .Q (signal_6175) ) ;
    buf_clk cell_3645 ( .C (clk), .D (signal_6190), .Q (signal_6191) ) ;
    buf_clk cell_3661 ( .C (clk), .D (signal_6206), .Q (signal_6207) ) ;
    buf_clk cell_3677 ( .C (clk), .D (signal_6222), .Q (signal_6223) ) ;
    buf_clk cell_3693 ( .C (clk), .D (signal_6238), .Q (signal_6239) ) ;
    buf_clk cell_3709 ( .C (clk), .D (signal_6254), .Q (signal_6255) ) ;
    buf_clk cell_3725 ( .C (clk), .D (signal_6270), .Q (signal_6271) ) ;
    buf_clk cell_3741 ( .C (clk), .D (signal_6286), .Q (signal_6287) ) ;
    buf_clk cell_3757 ( .C (clk), .D (signal_6302), .Q (signal_6303) ) ;
    buf_clk cell_3773 ( .C (clk), .D (signal_6318), .Q (signal_6319) ) ;
    buf_clk cell_3789 ( .C (clk), .D (signal_6334), .Q (signal_6335) ) ;
    buf_clk cell_3805 ( .C (clk), .D (signal_6350), .Q (signal_6351) ) ;
    buf_clk cell_3821 ( .C (clk), .D (signal_6366), .Q (signal_6367) ) ;
    buf_clk cell_3837 ( .C (clk), .D (signal_6382), .Q (signal_6383) ) ;
    buf_clk cell_3853 ( .C (clk), .D (signal_6398), .Q (signal_6399) ) ;
    buf_clk cell_3869 ( .C (clk), .D (signal_6414), .Q (signal_6415) ) ;
    buf_clk cell_3885 ( .C (clk), .D (signal_6430), .Q (signal_6431) ) ;
    buf_clk cell_3901 ( .C (clk), .D (signal_6446), .Q (signal_6447) ) ;
    buf_clk cell_3917 ( .C (clk), .D (signal_6462), .Q (signal_6463) ) ;
    buf_clk cell_3933 ( .C (clk), .D (signal_6478), .Q (signal_6479) ) ;
    buf_clk cell_3949 ( .C (clk), .D (signal_6494), .Q (signal_6495) ) ;
    buf_clk cell_3965 ( .C (clk), .D (signal_6510), .Q (signal_6511) ) ;
    buf_clk cell_3981 ( .C (clk), .D (signal_6526), .Q (signal_6527) ) ;
    buf_clk cell_3997 ( .C (clk), .D (signal_6542), .Q (signal_6543) ) ;
    buf_clk cell_4013 ( .C (clk), .D (signal_6558), .Q (signal_6559) ) ;
    buf_clk cell_4029 ( .C (clk), .D (signal_6574), .Q (signal_6575) ) ;
    buf_clk cell_4045 ( .C (clk), .D (signal_6590), .Q (signal_6591) ) ;
    buf_clk cell_4061 ( .C (clk), .D (signal_6606), .Q (signal_6607) ) ;
    buf_clk cell_4077 ( .C (clk), .D (signal_6622), .Q (signal_6623) ) ;
    buf_clk cell_4093 ( .C (clk), .D (signal_6638), .Q (signal_6639) ) ;
    buf_clk cell_4109 ( .C (clk), .D (signal_6654), .Q (signal_6655) ) ;
    buf_clk cell_4125 ( .C (clk), .D (signal_6670), .Q (signal_6671) ) ;
    buf_clk cell_4141 ( .C (clk), .D (signal_6686), .Q (signal_6687) ) ;
    buf_clk cell_4157 ( .C (clk), .D (signal_6702), .Q (signal_6703) ) ;
    buf_clk cell_4173 ( .C (clk), .D (signal_6718), .Q (signal_6719) ) ;
    buf_clk cell_4189 ( .C (clk), .D (signal_6734), .Q (signal_6735) ) ;
    buf_clk cell_4205 ( .C (clk), .D (signal_6750), .Q (signal_6751) ) ;
    buf_clk cell_4221 ( .C (clk), .D (signal_6766), .Q (signal_6767) ) ;
    buf_clk cell_4237 ( .C (clk), .D (signal_6782), .Q (signal_6783) ) ;
    buf_clk cell_4253 ( .C (clk), .D (signal_6798), .Q (signal_6799) ) ;
    buf_clk cell_4269 ( .C (clk), .D (signal_6814), .Q (signal_6815) ) ;
    buf_clk cell_4285 ( .C (clk), .D (signal_6830), .Q (signal_6831) ) ;
    buf_clk cell_4301 ( .C (clk), .D (signal_6846), .Q (signal_6847) ) ;
    buf_clk cell_4317 ( .C (clk), .D (signal_6862), .Q (signal_6863) ) ;
    buf_clk cell_4333 ( .C (clk), .D (signal_6878), .Q (signal_6879) ) ;
    buf_clk cell_4349 ( .C (clk), .D (signal_6894), .Q (signal_6895) ) ;
    buf_clk cell_4365 ( .C (clk), .D (signal_6910), .Q (signal_6911) ) ;
    buf_clk cell_4381 ( .C (clk), .D (signal_6926), .Q (signal_6927) ) ;
    buf_clk cell_4397 ( .C (clk), .D (signal_6942), .Q (signal_6943) ) ;
    buf_clk cell_4413 ( .C (clk), .D (signal_6958), .Q (signal_6959) ) ;
    buf_clk cell_4427 ( .C (clk), .D (signal_6972), .Q (signal_6973) ) ;
    buf_clk cell_4441 ( .C (clk), .D (signal_6986), .Q (signal_6987) ) ;
    buf_clk cell_4457 ( .C (clk), .D (signal_7002), .Q (signal_7003) ) ;
    buf_clk cell_4473 ( .C (clk), .D (signal_7018), .Q (signal_7019) ) ;
    buf_clk cell_4489 ( .C (clk), .D (signal_7034), .Q (signal_7035) ) ;
    buf_clk cell_4505 ( .C (clk), .D (signal_7050), .Q (signal_7051) ) ;
    buf_clk cell_4521 ( .C (clk), .D (signal_7066), .Q (signal_7067) ) ;
    buf_clk cell_4537 ( .C (clk), .D (signal_7082), .Q (signal_7083) ) ;
    buf_clk cell_4553 ( .C (clk), .D (signal_7098), .Q (signal_7099) ) ;
    buf_clk cell_4569 ( .C (clk), .D (signal_7114), .Q (signal_7115) ) ;
    buf_clk cell_4585 ( .C (clk), .D (signal_7130), .Q (signal_7131) ) ;
    buf_clk cell_4601 ( .C (clk), .D (signal_7146), .Q (signal_7147) ) ;
    buf_clk cell_4617 ( .C (clk), .D (signal_7162), .Q (signal_7163) ) ;
    buf_clk cell_4633 ( .C (clk), .D (signal_7178), .Q (signal_7179) ) ;
    buf_clk cell_4649 ( .C (clk), .D (signal_7194), .Q (signal_7195) ) ;
    buf_clk cell_4665 ( .C (clk), .D (signal_7210), .Q (signal_7211) ) ;
    buf_clk cell_4681 ( .C (clk), .D (signal_7226), .Q (signal_7227) ) ;
    buf_clk cell_4697 ( .C (clk), .D (signal_7242), .Q (signal_7243) ) ;
    buf_clk cell_4713 ( .C (clk), .D (signal_7258), .Q (signal_7259) ) ;
    buf_clk cell_4729 ( .C (clk), .D (signal_7274), .Q (signal_7275) ) ;
    buf_clk cell_4745 ( .C (clk), .D (signal_7290), .Q (signal_7291) ) ;
    buf_clk cell_4761 ( .C (clk), .D (signal_7306), .Q (signal_7307) ) ;
    buf_clk cell_4777 ( .C (clk), .D (signal_7322), .Q (signal_7323) ) ;
    buf_clk cell_4793 ( .C (clk), .D (signal_7338), .Q (signal_7339) ) ;
    buf_clk cell_4809 ( .C (clk), .D (signal_7354), .Q (signal_7355) ) ;
    buf_clk cell_4825 ( .C (clk), .D (signal_7370), .Q (signal_7371) ) ;
    buf_clk cell_4841 ( .C (clk), .D (signal_7386), .Q (signal_7387) ) ;
    buf_clk cell_4857 ( .C (clk), .D (signal_7402), .Q (signal_7403) ) ;
    buf_clk cell_4873 ( .C (clk), .D (signal_7418), .Q (signal_7419) ) ;
    buf_clk cell_4889 ( .C (clk), .D (signal_7434), .Q (signal_7435) ) ;
    buf_clk cell_4905 ( .C (clk), .D (signal_7450), .Q (signal_7451) ) ;
    buf_clk cell_4921 ( .C (clk), .D (signal_7466), .Q (signal_7467) ) ;
    buf_clk cell_4937 ( .C (clk), .D (signal_7482), .Q (signal_7483) ) ;
    buf_clk cell_4953 ( .C (clk), .D (signal_7498), .Q (signal_7499) ) ;
    buf_clk cell_4969 ( .C (clk), .D (signal_7514), .Q (signal_7515) ) ;
    buf_clk cell_4985 ( .C (clk), .D (signal_7530), .Q (signal_7531) ) ;
    buf_clk cell_5001 ( .C (clk), .D (signal_7546), .Q (signal_7547) ) ;
    buf_clk cell_5017 ( .C (clk), .D (signal_7562), .Q (signal_7563) ) ;
    buf_clk cell_5033 ( .C (clk), .D (signal_7578), .Q (signal_7579) ) ;
    buf_clk cell_5049 ( .C (clk), .D (signal_7594), .Q (signal_7595) ) ;
    buf_clk cell_5065 ( .C (clk), .D (signal_7610), .Q (signal_7611) ) ;
    buf_clk cell_5081 ( .C (clk), .D (signal_7626), .Q (signal_7627) ) ;
    buf_clk cell_5097 ( .C (clk), .D (signal_7642), .Q (signal_7643) ) ;
    buf_clk cell_5113 ( .C (clk), .D (signal_7658), .Q (signal_7659) ) ;
    buf_clk cell_5129 ( .C (clk), .D (signal_7674), .Q (signal_7675) ) ;
    buf_clk cell_5145 ( .C (clk), .D (signal_7690), .Q (signal_7691) ) ;
    buf_clk cell_5161 ( .C (clk), .D (signal_7706), .Q (signal_7707) ) ;
    buf_clk cell_5177 ( .C (clk), .D (signal_7722), .Q (signal_7723) ) ;
    buf_clk cell_5193 ( .C (clk), .D (signal_7738), .Q (signal_7739) ) ;
    buf_clk cell_5209 ( .C (clk), .D (signal_7754), .Q (signal_7755) ) ;
    buf_clk cell_5225 ( .C (clk), .D (signal_7770), .Q (signal_7771) ) ;
    buf_clk cell_5241 ( .C (clk), .D (signal_7786), .Q (signal_7787) ) ;
    buf_clk cell_5257 ( .C (clk), .D (signal_7802), .Q (signal_7803) ) ;
    buf_clk cell_5273 ( .C (clk), .D (signal_7818), .Q (signal_7819) ) ;
    buf_clk cell_5289 ( .C (clk), .D (signal_7834), .Q (signal_7835) ) ;
    buf_clk cell_5305 ( .C (clk), .D (signal_7850), .Q (signal_7851) ) ;
    buf_clk cell_5321 ( .C (clk), .D (signal_7866), .Q (signal_7867) ) ;
    buf_clk cell_5337 ( .C (clk), .D (signal_7882), .Q (signal_7883) ) ;
    buf_clk cell_5353 ( .C (clk), .D (signal_7898), .Q (signal_7899) ) ;
    buf_clk cell_5369 ( .C (clk), .D (signal_7914), .Q (signal_7915) ) ;
    buf_clk cell_5385 ( .C (clk), .D (signal_7930), .Q (signal_7931) ) ;
    buf_clk cell_5401 ( .C (clk), .D (signal_7946), .Q (signal_7947) ) ;
    buf_clk cell_5417 ( .C (clk), .D (signal_7962), .Q (signal_7963) ) ;
    buf_clk cell_5433 ( .C (clk), .D (signal_7978), .Q (signal_7979) ) ;
    buf_clk cell_5449 ( .C (clk), .D (signal_7994), .Q (signal_7995) ) ;
    buf_clk cell_5465 ( .C (clk), .D (signal_8010), .Q (signal_8011) ) ;
    buf_clk cell_5481 ( .C (clk), .D (signal_8026), .Q (signal_8027) ) ;
    buf_clk cell_5497 ( .C (clk), .D (signal_8042), .Q (signal_8043) ) ;
    buf_clk cell_5513 ( .C (clk), .D (signal_8058), .Q (signal_8059) ) ;
    buf_clk cell_5529 ( .C (clk), .D (signal_8074), .Q (signal_8075) ) ;
    buf_clk cell_5545 ( .C (clk), .D (signal_8090), .Q (signal_8091) ) ;
    buf_clk cell_5561 ( .C (clk), .D (signal_8106), .Q (signal_8107) ) ;
    buf_clk cell_5577 ( .C (clk), .D (signal_8122), .Q (signal_8123) ) ;
    buf_clk cell_5593 ( .C (clk), .D (signal_8138), .Q (signal_8139) ) ;
    buf_clk cell_5609 ( .C (clk), .D (signal_8154), .Q (signal_8155) ) ;
    buf_clk cell_5625 ( .C (clk), .D (signal_8170), .Q (signal_8171) ) ;
    buf_clk cell_5641 ( .C (clk), .D (signal_8186), .Q (signal_8187) ) ;
    buf_clk cell_5657 ( .C (clk), .D (signal_8202), .Q (signal_8203) ) ;
    buf_clk cell_5673 ( .C (clk), .D (signal_8218), .Q (signal_8219) ) ;
    buf_clk cell_5689 ( .C (clk), .D (signal_8234), .Q (signal_8235) ) ;
    buf_clk cell_5705 ( .C (clk), .D (signal_8250), .Q (signal_8251) ) ;
    buf_clk cell_5721 ( .C (clk), .D (signal_8266), .Q (signal_8267) ) ;
    buf_clk cell_5737 ( .C (clk), .D (signal_8282), .Q (signal_8283) ) ;
    buf_clk cell_5753 ( .C (clk), .D (signal_8298), .Q (signal_8299) ) ;
    buf_clk cell_5769 ( .C (clk), .D (signal_8314), .Q (signal_8315) ) ;
    buf_clk cell_5785 ( .C (clk), .D (signal_8330), .Q (signal_8331) ) ;
    buf_clk cell_5801 ( .C (clk), .D (signal_8346), .Q (signal_8347) ) ;
    buf_clk cell_5817 ( .C (clk), .D (signal_8362), .Q (signal_8363) ) ;
    buf_clk cell_5833 ( .C (clk), .D (signal_8378), .Q (signal_8379) ) ;
    buf_clk cell_5849 ( .C (clk), .D (signal_8394), .Q (signal_8395) ) ;
    buf_clk cell_5865 ( .C (clk), .D (signal_8410), .Q (signal_8411) ) ;
    buf_clk cell_5881 ( .C (clk), .D (signal_8426), .Q (signal_8427) ) ;
    buf_clk cell_5897 ( .C (clk), .D (signal_8442), .Q (signal_8443) ) ;
    buf_clk cell_5913 ( .C (clk), .D (signal_8458), .Q (signal_8459) ) ;
    buf_clk cell_5929 ( .C (clk), .D (signal_8474), .Q (signal_8475) ) ;
    buf_clk cell_5945 ( .C (clk), .D (signal_8490), .Q (signal_8491) ) ;
    buf_clk cell_5961 ( .C (clk), .D (signal_8506), .Q (signal_8507) ) ;
    buf_clk cell_5977 ( .C (clk), .D (signal_8522), .Q (signal_8523) ) ;
    buf_clk cell_5993 ( .C (clk), .D (signal_8538), .Q (signal_8539) ) ;
    buf_clk cell_6009 ( .C (clk), .D (signal_8554), .Q (signal_8555) ) ;
    buf_clk cell_6025 ( .C (clk), .D (signal_8570), .Q (signal_8571) ) ;
    buf_clk cell_6041 ( .C (clk), .D (signal_8586), .Q (signal_8587) ) ;
    buf_clk cell_6057 ( .C (clk), .D (signal_8602), .Q (signal_8603) ) ;
    buf_clk cell_6073 ( .C (clk), .D (signal_8618), .Q (signal_8619) ) ;
    buf_clk cell_6089 ( .C (clk), .D (signal_8634), .Q (signal_8635) ) ;
    buf_clk cell_6105 ( .C (clk), .D (signal_8650), .Q (signal_8651) ) ;
    buf_clk cell_6121 ( .C (clk), .D (signal_8666), .Q (signal_8667) ) ;
    buf_clk cell_6137 ( .C (clk), .D (signal_8682), .Q (signal_8683) ) ;
    buf_clk cell_6153 ( .C (clk), .D (signal_8698), .Q (signal_8699) ) ;
    buf_clk cell_6169 ( .C (clk), .D (signal_8714), .Q (signal_8715) ) ;
    buf_clk cell_6185 ( .C (clk), .D (signal_8730), .Q (signal_8731) ) ;
    buf_clk cell_6201 ( .C (clk), .D (signal_8746), .Q (signal_8747) ) ;
    buf_clk cell_6217 ( .C (clk), .D (signal_8762), .Q (signal_8763) ) ;
    buf_clk cell_6233 ( .C (clk), .D (signal_8778), .Q (signal_8779) ) ;
    buf_clk cell_6249 ( .C (clk), .D (signal_8794), .Q (signal_8795) ) ;
    buf_clk cell_6265 ( .C (clk), .D (signal_8810), .Q (signal_8811) ) ;
    buf_clk cell_6281 ( .C (clk), .D (signal_8826), .Q (signal_8827) ) ;
    buf_clk cell_6297 ( .C (clk), .D (signal_8842), .Q (signal_8843) ) ;
    buf_clk cell_6313 ( .C (clk), .D (signal_8858), .Q (signal_8859) ) ;
    buf_clk cell_6329 ( .C (clk), .D (signal_8874), .Q (signal_8875) ) ;
    buf_clk cell_6345 ( .C (clk), .D (signal_8890), .Q (signal_8891) ) ;
    buf_clk cell_6361 ( .C (clk), .D (signal_8906), .Q (signal_8907) ) ;
    buf_clk cell_6377 ( .C (clk), .D (signal_8922), .Q (signal_8923) ) ;
    buf_clk cell_6393 ( .C (clk), .D (signal_8938), .Q (signal_8939) ) ;
    buf_clk cell_6409 ( .C (clk), .D (signal_8954), .Q (signal_8955) ) ;
    buf_clk cell_6425 ( .C (clk), .D (signal_8970), .Q (signal_8971) ) ;
    buf_clk cell_6441 ( .C (clk), .D (signal_8986), .Q (signal_8987) ) ;
    buf_clk cell_6457 ( .C (clk), .D (signal_9002), .Q (signal_9003) ) ;
    buf_clk cell_6473 ( .C (clk), .D (signal_9018), .Q (signal_9019) ) ;
    buf_clk cell_6489 ( .C (clk), .D (signal_9034), .Q (signal_9035) ) ;
    buf_clk cell_6505 ( .C (clk), .D (signal_9050), .Q (signal_9051) ) ;
    buf_clk cell_6521 ( .C (clk), .D (signal_9066), .Q (signal_9067) ) ;
    buf_clk cell_6537 ( .C (clk), .D (signal_9082), .Q (signal_9083) ) ;
    buf_clk cell_6553 ( .C (clk), .D (signal_9098), .Q (signal_9099) ) ;
    buf_clk cell_6569 ( .C (clk), .D (signal_9114), .Q (signal_9115) ) ;
    buf_clk cell_6585 ( .C (clk), .D (signal_9130), .Q (signal_9131) ) ;
    buf_clk cell_6601 ( .C (clk), .D (signal_9146), .Q (signal_9147) ) ;
    buf_clk cell_6617 ( .C (clk), .D (signal_9162), .Q (signal_9163) ) ;
    buf_clk cell_6633 ( .C (clk), .D (signal_9178), .Q (signal_9179) ) ;
    buf_clk cell_6649 ( .C (clk), .D (signal_9194), .Q (signal_9195) ) ;
    buf_clk cell_6665 ( .C (clk), .D (signal_9210), .Q (signal_9211) ) ;
    buf_clk cell_6681 ( .C (clk), .D (signal_9226), .Q (signal_9227) ) ;
    buf_clk cell_6697 ( .C (clk), .D (signal_9242), .Q (signal_9243) ) ;
    buf_clk cell_6713 ( .C (clk), .D (signal_9258), .Q (signal_9259) ) ;
    buf_clk cell_6729 ( .C (clk), .D (signal_9274), .Q (signal_9275) ) ;
    buf_clk cell_6745 ( .C (clk), .D (signal_9290), .Q (signal_9291) ) ;
    buf_clk cell_6761 ( .C (clk), .D (signal_9306), .Q (signal_9307) ) ;
    buf_clk cell_6777 ( .C (clk), .D (signal_9322), .Q (signal_9323) ) ;
    buf_clk cell_6793 ( .C (clk), .D (signal_9338), .Q (signal_9339) ) ;
    buf_clk cell_6809 ( .C (clk), .D (signal_9354), .Q (signal_9355) ) ;
    buf_clk cell_6825 ( .C (clk), .D (signal_9370), .Q (signal_9371) ) ;
    buf_clk cell_6841 ( .C (clk), .D (signal_9386), .Q (signal_9387) ) ;
    buf_clk cell_6857 ( .C (clk), .D (signal_9402), .Q (signal_9403) ) ;
    buf_clk cell_6873 ( .C (clk), .D (signal_9418), .Q (signal_9419) ) ;
    buf_clk cell_6889 ( .C (clk), .D (signal_9434), .Q (signal_9435) ) ;
    buf_clk cell_6905 ( .C (clk), .D (signal_9450), .Q (signal_9451) ) ;
    buf_clk cell_6921 ( .C (clk), .D (signal_9466), .Q (signal_9467) ) ;
    buf_clk cell_6937 ( .C (clk), .D (signal_9482), .Q (signal_9483) ) ;
    buf_clk cell_6953 ( .C (clk), .D (signal_9498), .Q (signal_9499) ) ;
    buf_clk cell_6969 ( .C (clk), .D (signal_9514), .Q (signal_9515) ) ;
    buf_clk cell_6985 ( .C (clk), .D (signal_9530), .Q (signal_9531) ) ;
    buf_clk cell_7001 ( .C (clk), .D (signal_9546), .Q (signal_9547) ) ;
    buf_clk cell_7017 ( .C (clk), .D (signal_9562), .Q (signal_9563) ) ;
    buf_clk cell_7033 ( .C (clk), .D (signal_9578), .Q (signal_9579) ) ;
    buf_clk cell_7049 ( .C (clk), .D (signal_9594), .Q (signal_9595) ) ;
    buf_clk cell_7065 ( .C (clk), .D (signal_9610), .Q (signal_9611) ) ;
    buf_clk cell_7081 ( .C (clk), .D (signal_9626), .Q (signal_9627) ) ;
    buf_clk cell_7097 ( .C (clk), .D (signal_9642), .Q (signal_9643) ) ;
    buf_clk cell_7113 ( .C (clk), .D (signal_9658), .Q (signal_9659) ) ;
    buf_clk cell_7129 ( .C (clk), .D (signal_9674), .Q (signal_9675) ) ;
    buf_clk cell_7145 ( .C (clk), .D (signal_9690), .Q (signal_9691) ) ;
    buf_clk cell_7161 ( .C (clk), .D (signal_9706), .Q (signal_9707) ) ;
    buf_clk cell_7177 ( .C (clk), .D (signal_9722), .Q (signal_9723) ) ;
    buf_clk cell_7193 ( .C (clk), .D (signal_9738), .Q (signal_9739) ) ;
    buf_clk cell_7209 ( .C (clk), .D (signal_9754), .Q (signal_9755) ) ;
    buf_clk cell_7225 ( .C (clk), .D (signal_9770), .Q (signal_9771) ) ;
    buf_clk cell_7241 ( .C (clk), .D (signal_9786), .Q (signal_9787) ) ;
    buf_clk cell_7257 ( .C (clk), .D (signal_9802), .Q (signal_9803) ) ;
    buf_clk cell_7273 ( .C (clk), .D (signal_9818), .Q (signal_9819) ) ;
    buf_clk cell_7289 ( .C (clk), .D (signal_9834), .Q (signal_9835) ) ;
    buf_clk cell_7305 ( .C (clk), .D (signal_9850), .Q (signal_9851) ) ;
    buf_clk cell_7321 ( .C (clk), .D (signal_9866), .Q (signal_9867) ) ;
    buf_clk cell_7337 ( .C (clk), .D (signal_9882), .Q (signal_9883) ) ;
    buf_clk cell_7353 ( .C (clk), .D (signal_9898), .Q (signal_9899) ) ;
    buf_clk cell_7369 ( .C (clk), .D (signal_9914), .Q (signal_9915) ) ;
    buf_clk cell_7385 ( .C (clk), .D (signal_9930), .Q (signal_9931) ) ;
    buf_clk cell_7401 ( .C (clk), .D (signal_9946), .Q (signal_9947) ) ;
    buf_clk cell_7417 ( .C (clk), .D (signal_9962), .Q (signal_9963) ) ;
    buf_clk cell_7433 ( .C (clk), .D (signal_9978), .Q (signal_9979) ) ;
    buf_clk cell_7449 ( .C (clk), .D (signal_9994), .Q (signal_9995) ) ;
    buf_clk cell_7465 ( .C (clk), .D (signal_10010), .Q (signal_10011) ) ;
    buf_clk cell_7481 ( .C (clk), .D (signal_10026), .Q (signal_10027) ) ;
    buf_clk cell_7497 ( .C (clk), .D (signal_10042), .Q (signal_10043) ) ;
    buf_clk cell_7513 ( .C (clk), .D (signal_10058), .Q (signal_10059) ) ;
    buf_clk cell_7529 ( .C (clk), .D (signal_10074), .Q (signal_10075) ) ;
    buf_clk cell_7545 ( .C (clk), .D (signal_10090), .Q (signal_10091) ) ;
    buf_clk cell_7561 ( .C (clk), .D (signal_10106), .Q (signal_10107) ) ;
    buf_clk cell_7577 ( .C (clk), .D (signal_10122), .Q (signal_10123) ) ;
    buf_clk cell_7593 ( .C (clk), .D (signal_10138), .Q (signal_10139) ) ;
    buf_clk cell_7609 ( .C (clk), .D (signal_10154), .Q (signal_10155) ) ;
    buf_clk cell_7625 ( .C (clk), .D (signal_10170), .Q (signal_10171) ) ;
    buf_clk cell_7641 ( .C (clk), .D (signal_10186), .Q (signal_10187) ) ;
    buf_clk cell_7657 ( .C (clk), .D (signal_10202), .Q (signal_10203) ) ;
    buf_clk cell_7673 ( .C (clk), .D (signal_10218), .Q (signal_10219) ) ;
    buf_clk cell_7689 ( .C (clk), .D (signal_10234), .Q (signal_10235) ) ;
    buf_clk cell_7705 ( .C (clk), .D (signal_10250), .Q (signal_10251) ) ;
    buf_clk cell_7721 ( .C (clk), .D (signal_10266), .Q (signal_10267) ) ;
    buf_clk cell_7737 ( .C (clk), .D (signal_10282), .Q (signal_10283) ) ;
    buf_clk cell_7753 ( .C (clk), .D (signal_10298), .Q (signal_10299) ) ;
    buf_clk cell_7769 ( .C (clk), .D (signal_10314), .Q (signal_10315) ) ;
    buf_clk cell_7785 ( .C (clk), .D (signal_10330), .Q (signal_10331) ) ;
    buf_clk cell_7801 ( .C (clk), .D (signal_10346), .Q (signal_10347) ) ;
    buf_clk cell_7817 ( .C (clk), .D (signal_10362), .Q (signal_10363) ) ;
    buf_clk cell_7833 ( .C (clk), .D (signal_10378), .Q (signal_10379) ) ;
    buf_clk cell_7849 ( .C (clk), .D (signal_10394), .Q (signal_10395) ) ;
    buf_clk cell_7865 ( .C (clk), .D (signal_10410), .Q (signal_10411) ) ;
    buf_clk cell_7881 ( .C (clk), .D (signal_10426), .Q (signal_10427) ) ;
    buf_clk cell_7897 ( .C (clk), .D (signal_10442), .Q (signal_10443) ) ;
    buf_clk cell_7913 ( .C (clk), .D (signal_10458), .Q (signal_10459) ) ;
    buf_clk cell_7929 ( .C (clk), .D (signal_10474), .Q (signal_10475) ) ;
    buf_clk cell_7945 ( .C (clk), .D (signal_10490), .Q (signal_10491) ) ;
    buf_clk cell_7961 ( .C (clk), .D (signal_10506), .Q (signal_10507) ) ;
    buf_clk cell_7977 ( .C (clk), .D (signal_10522), .Q (signal_10523) ) ;
    buf_clk cell_7993 ( .C (clk), .D (signal_10538), .Q (signal_10539) ) ;
    buf_clk cell_8009 ( .C (clk), .D (signal_10554), .Q (signal_10555) ) ;
    buf_clk cell_8025 ( .C (clk), .D (signal_10570), .Q (signal_10571) ) ;
    buf_clk cell_8041 ( .C (clk), .D (signal_10586), .Q (signal_10587) ) ;
    buf_clk cell_8057 ( .C (clk), .D (signal_10602), .Q (signal_10603) ) ;
    buf_clk cell_8073 ( .C (clk), .D (signal_10618), .Q (signal_10619) ) ;
    buf_clk cell_8089 ( .C (clk), .D (signal_10634), .Q (signal_10635) ) ;
    buf_clk cell_8105 ( .C (clk), .D (signal_10650), .Q (signal_10651) ) ;
    buf_clk cell_8121 ( .C (clk), .D (signal_10666), .Q (signal_10667) ) ;
    buf_clk cell_8137 ( .C (clk), .D (signal_10682), .Q (signal_10683) ) ;
    buf_clk cell_8153 ( .C (clk), .D (signal_10698), .Q (signal_10699) ) ;
    buf_clk cell_8169 ( .C (clk), .D (signal_10714), .Q (signal_10715) ) ;
    buf_clk cell_8185 ( .C (clk), .D (signal_10730), .Q (signal_10731) ) ;
    buf_clk cell_8201 ( .C (clk), .D (signal_10746), .Q (signal_10747) ) ;
    buf_clk cell_8217 ( .C (clk), .D (signal_10762), .Q (signal_10763) ) ;
    buf_clk cell_8233 ( .C (clk), .D (signal_10778), .Q (signal_10779) ) ;
    buf_clk cell_8249 ( .C (clk), .D (signal_10794), .Q (signal_10795) ) ;
    buf_clk cell_8265 ( .C (clk), .D (signal_10810), .Q (signal_10811) ) ;
    buf_clk cell_8281 ( .C (clk), .D (signal_10826), .Q (signal_10827) ) ;
    buf_clk cell_8297 ( .C (clk), .D (signal_10842), .Q (signal_10843) ) ;
    buf_clk cell_8313 ( .C (clk), .D (signal_10858), .Q (signal_10859) ) ;
    buf_clk cell_8329 ( .C (clk), .D (signal_10874), .Q (signal_10875) ) ;
    buf_clk cell_8345 ( .C (clk), .D (signal_10890), .Q (signal_10891) ) ;
    buf_clk cell_8361 ( .C (clk), .D (signal_10906), .Q (signal_10907) ) ;
    buf_clk cell_8377 ( .C (clk), .D (signal_10922), .Q (signal_10923) ) ;
    buf_clk cell_8393 ( .C (clk), .D (signal_10938), .Q (signal_10939) ) ;
    buf_clk cell_8409 ( .C (clk), .D (signal_10954), .Q (signal_10955) ) ;
    buf_clk cell_8425 ( .C (clk), .D (signal_10970), .Q (signal_10971) ) ;
    buf_clk cell_8441 ( .C (clk), .D (signal_10986), .Q (signal_10987) ) ;
    buf_clk cell_8457 ( .C (clk), .D (signal_11002), .Q (signal_11003) ) ;
    buf_clk cell_8473 ( .C (clk), .D (signal_11018), .Q (signal_11019) ) ;
    buf_clk cell_8489 ( .C (clk), .D (signal_11034), .Q (signal_11035) ) ;
    buf_clk cell_8505 ( .C (clk), .D (signal_11050), .Q (signal_11051) ) ;
    buf_clk cell_8521 ( .C (clk), .D (signal_11066), .Q (signal_11067) ) ;
    buf_clk cell_8537 ( .C (clk), .D (signal_11082), .Q (signal_11083) ) ;
    buf_clk cell_8553 ( .C (clk), .D (signal_11098), .Q (signal_11099) ) ;
    buf_clk cell_8569 ( .C (clk), .D (signal_11114), .Q (signal_11115) ) ;
    buf_clk cell_8585 ( .C (clk), .D (signal_11130), .Q (signal_11131) ) ;
    buf_clk cell_8601 ( .C (clk), .D (signal_11146), .Q (signal_11147) ) ;
    buf_clk cell_8617 ( .C (clk), .D (signal_11162), .Q (signal_11163) ) ;
    buf_clk cell_8633 ( .C (clk), .D (signal_11178), .Q (signal_11179) ) ;
    buf_clk cell_8649 ( .C (clk), .D (signal_11194), .Q (signal_11195) ) ;
    buf_clk cell_8665 ( .C (clk), .D (signal_11210), .Q (signal_11211) ) ;
    buf_clk cell_8681 ( .C (clk), .D (signal_11226), .Q (signal_11227) ) ;
    buf_clk cell_8697 ( .C (clk), .D (signal_11242), .Q (signal_11243) ) ;
    buf_clk cell_8713 ( .C (clk), .D (signal_11258), .Q (signal_11259) ) ;
    buf_clk cell_8729 ( .C (clk), .D (signal_11274), .Q (signal_11275) ) ;
    buf_clk cell_8745 ( .C (clk), .D (signal_11290), .Q (signal_11291) ) ;
    buf_clk cell_8761 ( .C (clk), .D (signal_11306), .Q (signal_11307) ) ;
    buf_clk cell_8777 ( .C (clk), .D (signal_11322), .Q (signal_11323) ) ;
    buf_clk cell_8793 ( .C (clk), .D (signal_11338), .Q (signal_11339) ) ;
    buf_clk cell_8809 ( .C (clk), .D (signal_11354), .Q (signal_11355) ) ;
    buf_clk cell_8825 ( .C (clk), .D (signal_11370), .Q (signal_11371) ) ;
    buf_clk cell_8841 ( .C (clk), .D (signal_11386), .Q (signal_11387) ) ;
    buf_clk cell_8857 ( .C (clk), .D (signal_11402), .Q (signal_11403) ) ;
    buf_clk cell_8873 ( .C (clk), .D (signal_11418), .Q (signal_11419) ) ;
    buf_clk cell_8889 ( .C (clk), .D (signal_11434), .Q (signal_11435) ) ;
    buf_clk cell_8905 ( .C (clk), .D (signal_11450), .Q (signal_11451) ) ;
    buf_clk cell_8921 ( .C (clk), .D (signal_11466), .Q (signal_11467) ) ;
    buf_clk cell_8937 ( .C (clk), .D (signal_11482), .Q (signal_11483) ) ;
    buf_clk cell_8953 ( .C (clk), .D (signal_11498), .Q (signal_11499) ) ;
    buf_clk cell_8969 ( .C (clk), .D (signal_11514), .Q (signal_11515) ) ;
    buf_clk cell_8985 ( .C (clk), .D (signal_11530), .Q (signal_11531) ) ;
    buf_clk cell_9001 ( .C (clk), .D (signal_11546), .Q (signal_11547) ) ;
    buf_clk cell_9017 ( .C (clk), .D (signal_11562), .Q (signal_11563) ) ;
    buf_clk cell_9033 ( .C (clk), .D (signal_11578), .Q (signal_11579) ) ;
    buf_clk cell_9049 ( .C (clk), .D (signal_11594), .Q (signal_11595) ) ;
    buf_clk cell_9065 ( .C (clk), .D (signal_11610), .Q (signal_11611) ) ;
    buf_clk cell_9081 ( .C (clk), .D (signal_11626), .Q (signal_11627) ) ;
    buf_clk cell_9097 ( .C (clk), .D (signal_11642), .Q (signal_11643) ) ;
    buf_clk cell_9113 ( .C (clk), .D (signal_11658), .Q (signal_11659) ) ;
    buf_clk cell_9129 ( .C (clk), .D (signal_11674), .Q (signal_11675) ) ;
    buf_clk cell_9145 ( .C (clk), .D (signal_11690), .Q (signal_11691) ) ;
    buf_clk cell_9161 ( .C (clk), .D (signal_11706), .Q (signal_11707) ) ;
    buf_clk cell_9177 ( .C (clk), .D (signal_11722), .Q (signal_11723) ) ;
    buf_clk cell_9193 ( .C (clk), .D (signal_11738), .Q (signal_11739) ) ;
    buf_clk cell_9209 ( .C (clk), .D (signal_11754), .Q (signal_11755) ) ;
    buf_clk cell_9225 ( .C (clk), .D (signal_11770), .Q (signal_11771) ) ;
    buf_clk cell_9241 ( .C (clk), .D (signal_11786), .Q (signal_11787) ) ;
    buf_clk cell_9257 ( .C (clk), .D (signal_11802), .Q (signal_11803) ) ;
    buf_clk cell_9273 ( .C (clk), .D (signal_11818), .Q (signal_11819) ) ;
    buf_clk cell_9289 ( .C (clk), .D (signal_11834), .Q (signal_11835) ) ;
    buf_clk cell_9305 ( .C (clk), .D (signal_11850), .Q (signal_11851) ) ;
    buf_clk cell_9321 ( .C (clk), .D (signal_11866), .Q (signal_11867) ) ;
    buf_clk cell_9337 ( .C (clk), .D (signal_11882), .Q (signal_11883) ) ;
    buf_clk cell_9353 ( .C (clk), .D (signal_11898), .Q (signal_11899) ) ;
    buf_clk cell_9369 ( .C (clk), .D (signal_11914), .Q (signal_11915) ) ;
    buf_clk cell_9385 ( .C (clk), .D (signal_11930), .Q (signal_11931) ) ;
    buf_clk cell_9401 ( .C (clk), .D (signal_11946), .Q (signal_11947) ) ;
    buf_clk cell_9417 ( .C (clk), .D (signal_11962), .Q (signal_11963) ) ;
    buf_clk cell_9433 ( .C (clk), .D (signal_11978), .Q (signal_11979) ) ;
    buf_clk cell_9449 ( .C (clk), .D (signal_11994), .Q (signal_11995) ) ;
    buf_clk cell_9465 ( .C (clk), .D (signal_12010), .Q (signal_12011) ) ;
    buf_clk cell_9481 ( .C (clk), .D (signal_12026), .Q (signal_12027) ) ;
    buf_clk cell_9497 ( .C (clk), .D (signal_12042), .Q (signal_12043) ) ;
    buf_clk cell_9513 ( .C (clk), .D (signal_12058), .Q (signal_12059) ) ;
    buf_clk cell_9529 ( .C (clk), .D (signal_12074), .Q (signal_12075) ) ;
    buf_clk cell_9545 ( .C (clk), .D (signal_12090), .Q (signal_12091) ) ;
    buf_clk cell_9561 ( .C (clk), .D (signal_12106), .Q (signal_12107) ) ;
    buf_clk cell_9577 ( .C (clk), .D (signal_12122), .Q (signal_12123) ) ;
    buf_clk cell_9593 ( .C (clk), .D (signal_12138), .Q (signal_12139) ) ;
    buf_clk cell_9609 ( .C (clk), .D (signal_12154), .Q (signal_12155) ) ;
    buf_clk cell_9625 ( .C (clk), .D (signal_12170), .Q (signal_12171) ) ;
    buf_clk cell_9641 ( .C (clk), .D (signal_12186), .Q (signal_12187) ) ;
    buf_clk cell_9657 ( .C (clk), .D (signal_12202), .Q (signal_12203) ) ;
    buf_clk cell_9673 ( .C (clk), .D (signal_12218), .Q (signal_12219) ) ;
    buf_clk cell_9689 ( .C (clk), .D (signal_12234), .Q (signal_12235) ) ;
    buf_clk cell_9705 ( .C (clk), .D (signal_12250), .Q (signal_12251) ) ;
    buf_clk cell_9721 ( .C (clk), .D (signal_12266), .Q (signal_12267) ) ;
    buf_clk cell_9737 ( .C (clk), .D (signal_12282), .Q (signal_12283) ) ;
    buf_clk cell_9753 ( .C (clk), .D (signal_12298), .Q (signal_12299) ) ;
    buf_clk cell_9769 ( .C (clk), .D (signal_12314), .Q (signal_12315) ) ;
    buf_clk cell_9785 ( .C (clk), .D (signal_12330), .Q (signal_12331) ) ;
    buf_clk cell_9801 ( .C (clk), .D (signal_12346), .Q (signal_12347) ) ;
    buf_clk cell_9817 ( .C (clk), .D (signal_12362), .Q (signal_12363) ) ;
    buf_clk cell_9833 ( .C (clk), .D (signal_12378), .Q (signal_12379) ) ;
    buf_clk cell_9849 ( .C (clk), .D (signal_12394), .Q (signal_12395) ) ;
    buf_clk cell_9865 ( .C (clk), .D (signal_12410), .Q (signal_12411) ) ;
    buf_clk cell_9881 ( .C (clk), .D (signal_12426), .Q (signal_12427) ) ;
    buf_clk cell_9897 ( .C (clk), .D (signal_12442), .Q (signal_12443) ) ;
    buf_clk cell_9913 ( .C (clk), .D (signal_12458), .Q (signal_12459) ) ;
    buf_clk cell_9929 ( .C (clk), .D (signal_12474), .Q (signal_12475) ) ;
    buf_clk cell_9945 ( .C (clk), .D (signal_12490), .Q (signal_12491) ) ;
    buf_clk cell_9961 ( .C (clk), .D (signal_12506), .Q (signal_12507) ) ;
    buf_clk cell_9977 ( .C (clk), .D (signal_12522), .Q (signal_12523) ) ;
    buf_clk cell_9993 ( .C (clk), .D (signal_12538), .Q (signal_12539) ) ;
    buf_clk cell_10009 ( .C (clk), .D (signal_12554), .Q (signal_12555) ) ;
    buf_clk cell_10025 ( .C (clk), .D (signal_12570), .Q (signal_12571) ) ;
    buf_clk cell_10041 ( .C (clk), .D (signal_12586), .Q (signal_12587) ) ;
    buf_clk cell_10057 ( .C (clk), .D (signal_12602), .Q (signal_12603) ) ;
    buf_clk cell_10073 ( .C (clk), .D (signal_12618), .Q (signal_12619) ) ;
    buf_clk cell_10089 ( .C (clk), .D (signal_12634), .Q (signal_12635) ) ;
    buf_clk cell_10105 ( .C (clk), .D (signal_12650), .Q (signal_12651) ) ;
    buf_clk cell_10121 ( .C (clk), .D (signal_12666), .Q (signal_12667) ) ;
    buf_clk cell_10137 ( .C (clk), .D (signal_12682), .Q (signal_12683) ) ;
    buf_clk cell_10153 ( .C (clk), .D (signal_12698), .Q (signal_12699) ) ;
    buf_clk cell_10169 ( .C (clk), .D (signal_12714), .Q (signal_12715) ) ;
    buf_clk cell_10185 ( .C (clk), .D (signal_12730), .Q (signal_12731) ) ;
    buf_clk cell_10201 ( .C (clk), .D (signal_12746), .Q (signal_12747) ) ;
    buf_clk cell_10217 ( .C (clk), .D (signal_12762), .Q (signal_12763) ) ;
    buf_clk cell_10233 ( .C (clk), .D (signal_12778), .Q (signal_12779) ) ;
    buf_clk cell_10249 ( .C (clk), .D (signal_12794), .Q (signal_12795) ) ;
    buf_clk cell_10265 ( .C (clk), .D (signal_12810), .Q (signal_12811) ) ;
    buf_clk cell_10281 ( .C (clk), .D (signal_12826), .Q (signal_12827) ) ;
    buf_clk cell_10297 ( .C (clk), .D (signal_12842), .Q (signal_12843) ) ;
    buf_clk cell_10313 ( .C (clk), .D (signal_12858), .Q (signal_12859) ) ;
    buf_clk cell_10329 ( .C (clk), .D (signal_12874), .Q (signal_12875) ) ;
    buf_clk cell_10345 ( .C (clk), .D (signal_12890), .Q (signal_12891) ) ;
    buf_clk cell_10361 ( .C (clk), .D (signal_12906), .Q (signal_12907) ) ;
    buf_clk cell_10377 ( .C (clk), .D (signal_12922), .Q (signal_12923) ) ;
    buf_clk cell_10393 ( .C (clk), .D (signal_12938), .Q (signal_12939) ) ;
    buf_clk cell_10409 ( .C (clk), .D (signal_12954), .Q (signal_12955) ) ;
    buf_clk cell_10425 ( .C (clk), .D (signal_12970), .Q (signal_12971) ) ;
    buf_clk cell_10441 ( .C (clk), .D (signal_12986), .Q (signal_12987) ) ;
    buf_clk cell_10457 ( .C (clk), .D (signal_13002), .Q (signal_13003) ) ;
    buf_clk cell_10473 ( .C (clk), .D (signal_13018), .Q (signal_13019) ) ;
    buf_clk cell_10489 ( .C (clk), .D (signal_13034), .Q (signal_13035) ) ;
    buf_clk cell_10505 ( .C (clk), .D (signal_13050), .Q (signal_13051) ) ;
    buf_clk cell_10521 ( .C (clk), .D (signal_13066), .Q (signal_13067) ) ;
    buf_clk cell_10537 ( .C (clk), .D (signal_13082), .Q (signal_13083) ) ;
    buf_clk cell_10553 ( .C (clk), .D (signal_13098), .Q (signal_13099) ) ;
    buf_clk cell_10569 ( .C (clk), .D (signal_13114), .Q (signal_13115) ) ;
    buf_clk cell_10585 ( .C (clk), .D (signal_13130), .Q (signal_13131) ) ;
    buf_clk cell_10601 ( .C (clk), .D (signal_13146), .Q (signal_13147) ) ;
    buf_clk cell_10617 ( .C (clk), .D (signal_13162), .Q (signal_13163) ) ;
    buf_clk cell_10633 ( .C (clk), .D (signal_13178), .Q (signal_13179) ) ;
    buf_clk cell_10649 ( .C (clk), .D (signal_13194), .Q (signal_13195) ) ;
    buf_clk cell_10665 ( .C (clk), .D (signal_13210), .Q (signal_13211) ) ;
    buf_clk cell_10681 ( .C (clk), .D (signal_13226), .Q (signal_13227) ) ;
    buf_clk cell_10697 ( .C (clk), .D (signal_13242), .Q (signal_13243) ) ;
    buf_clk cell_10713 ( .C (clk), .D (signal_13258), .Q (signal_13259) ) ;
    buf_clk cell_10729 ( .C (clk), .D (signal_13274), .Q (signal_13275) ) ;
    buf_clk cell_10745 ( .C (clk), .D (signal_13290), .Q (signal_13291) ) ;
    buf_clk cell_10761 ( .C (clk), .D (signal_13306), .Q (signal_13307) ) ;
    buf_clk cell_10777 ( .C (clk), .D (signal_13322), .Q (signal_13323) ) ;
    buf_clk cell_10793 ( .C (clk), .D (signal_13338), .Q (signal_13339) ) ;
    buf_clk cell_10809 ( .C (clk), .D (signal_13354), .Q (signal_13355) ) ;
    buf_clk cell_10825 ( .C (clk), .D (signal_13370), .Q (signal_13371) ) ;
    buf_clk cell_10841 ( .C (clk), .D (signal_13386), .Q (signal_13387) ) ;
    buf_clk cell_10857 ( .C (clk), .D (signal_13402), .Q (signal_13403) ) ;
    buf_clk cell_10873 ( .C (clk), .D (signal_13418), .Q (signal_13419) ) ;
    buf_clk cell_10889 ( .C (clk), .D (signal_13434), .Q (signal_13435) ) ;
    buf_clk cell_10905 ( .C (clk), .D (signal_13450), .Q (signal_13451) ) ;
    buf_clk cell_10921 ( .C (clk), .D (signal_13466), .Q (signal_13467) ) ;
    buf_clk cell_10937 ( .C (clk), .D (signal_13482), .Q (signal_13483) ) ;
    buf_clk cell_10953 ( .C (clk), .D (signal_13498), .Q (signal_13499) ) ;
    buf_clk cell_10969 ( .C (clk), .D (signal_13514), .Q (signal_13515) ) ;
    buf_clk cell_10985 ( .C (clk), .D (signal_13530), .Q (signal_13531) ) ;
    buf_clk cell_11001 ( .C (clk), .D (signal_13546), .Q (signal_13547) ) ;
    buf_clk cell_11017 ( .C (clk), .D (signal_13562), .Q (signal_13563) ) ;
    buf_clk cell_11033 ( .C (clk), .D (signal_13578), .Q (signal_13579) ) ;
    buf_clk cell_11049 ( .C (clk), .D (signal_13594), .Q (signal_13595) ) ;
    buf_clk cell_11065 ( .C (clk), .D (signal_13610), .Q (signal_13611) ) ;
    buf_clk cell_11081 ( .C (clk), .D (signal_13626), .Q (signal_13627) ) ;
    buf_clk cell_11097 ( .C (clk), .D (signal_13642), .Q (signal_13643) ) ;
    buf_clk cell_11113 ( .C (clk), .D (signal_13658), .Q (signal_13659) ) ;
    buf_clk cell_11129 ( .C (clk), .D (signal_13674), .Q (signal_13675) ) ;
    buf_clk cell_11145 ( .C (clk), .D (signal_13690), .Q (signal_13691) ) ;
    buf_clk cell_11161 ( .C (clk), .D (signal_13706), .Q (signal_13707) ) ;
    buf_clk cell_11177 ( .C (clk), .D (signal_13722), .Q (signal_13723) ) ;
    buf_clk cell_11193 ( .C (clk), .D (signal_13738), .Q (signal_13739) ) ;
    buf_clk cell_11209 ( .C (clk), .D (signal_13754), .Q (signal_13755) ) ;
    buf_clk cell_11225 ( .C (clk), .D (signal_13770), .Q (signal_13771) ) ;
    buf_clk cell_11241 ( .C (clk), .D (signal_13786), .Q (signal_13787) ) ;
    buf_clk cell_11257 ( .C (clk), .D (signal_13802), .Q (signal_13803) ) ;
    buf_clk cell_11273 ( .C (clk), .D (signal_13818), .Q (signal_13819) ) ;
    buf_clk cell_11289 ( .C (clk), .D (signal_13834), .Q (signal_13835) ) ;
    buf_clk cell_11305 ( .C (clk), .D (signal_13850), .Q (signal_13851) ) ;
    buf_clk cell_11321 ( .C (clk), .D (signal_13866), .Q (signal_13867) ) ;
    buf_clk cell_11337 ( .C (clk), .D (signal_13882), .Q (signal_13883) ) ;
    buf_clk cell_11353 ( .C (clk), .D (signal_13898), .Q (signal_13899) ) ;
    buf_clk cell_11369 ( .C (clk), .D (signal_13914), .Q (signal_13915) ) ;
    buf_clk cell_11385 ( .C (clk), .D (signal_13930), .Q (signal_13931) ) ;
    buf_clk cell_11401 ( .C (clk), .D (signal_13946), .Q (signal_13947) ) ;
    buf_clk cell_11417 ( .C (clk), .D (signal_13962), .Q (signal_13963) ) ;
    buf_clk cell_11433 ( .C (clk), .D (signal_13978), .Q (signal_13979) ) ;
    buf_clk cell_11449 ( .C (clk), .D (signal_13994), .Q (signal_13995) ) ;
    buf_clk cell_11465 ( .C (clk), .D (signal_14010), .Q (signal_14011) ) ;
    buf_clk cell_11481 ( .C (clk), .D (signal_14026), .Q (signal_14027) ) ;
    buf_clk cell_11497 ( .C (clk), .D (signal_14042), .Q (signal_14043) ) ;
    buf_clk cell_11513 ( .C (clk), .D (signal_14058), .Q (signal_14059) ) ;
    buf_clk cell_11529 ( .C (clk), .D (signal_14074), .Q (signal_14075) ) ;
    buf_clk cell_11545 ( .C (clk), .D (signal_14090), .Q (signal_14091) ) ;
    buf_clk cell_11561 ( .C (clk), .D (signal_14106), .Q (signal_14107) ) ;
    buf_clk cell_11577 ( .C (clk), .D (signal_14122), .Q (signal_14123) ) ;
    buf_clk cell_11593 ( .C (clk), .D (signal_14138), .Q (signal_14139) ) ;
    buf_clk cell_11609 ( .C (clk), .D (signal_14154), .Q (signal_14155) ) ;
    buf_clk cell_11625 ( .C (clk), .D (signal_14170), .Q (signal_14171) ) ;
    buf_clk cell_11641 ( .C (clk), .D (signal_14186), .Q (signal_14187) ) ;
    buf_clk cell_11657 ( .C (clk), .D (signal_14202), .Q (signal_14203) ) ;
    buf_clk cell_11673 ( .C (clk), .D (signal_14218), .Q (signal_14219) ) ;
    buf_clk cell_11689 ( .C (clk), .D (signal_14234), .Q (signal_14235) ) ;
    buf_clk cell_11705 ( .C (clk), .D (signal_14250), .Q (signal_14251) ) ;
    buf_clk cell_11721 ( .C (clk), .D (signal_14266), .Q (signal_14267) ) ;
    buf_clk cell_11737 ( .C (clk), .D (signal_14282), .Q (signal_14283) ) ;
    buf_clk cell_11753 ( .C (clk), .D (signal_14298), .Q (signal_14299) ) ;
    buf_clk cell_11769 ( .C (clk), .D (signal_14314), .Q (signal_14315) ) ;
    buf_clk cell_11785 ( .C (clk), .D (signal_14330), .Q (signal_14331) ) ;
    buf_clk cell_11801 ( .C (clk), .D (signal_14346), .Q (signal_14347) ) ;
    buf_clk cell_11817 ( .C (clk), .D (signal_14362), .Q (signal_14363) ) ;
    buf_clk cell_11833 ( .C (clk), .D (signal_14378), .Q (signal_14379) ) ;
    buf_clk cell_11849 ( .C (clk), .D (signal_14394), .Q (signal_14395) ) ;
    buf_clk cell_11865 ( .C (clk), .D (signal_14410), .Q (signal_14411) ) ;
    buf_clk cell_11881 ( .C (clk), .D (signal_14426), .Q (signal_14427) ) ;
    buf_clk cell_11897 ( .C (clk), .D (signal_14442), .Q (signal_14443) ) ;
    buf_clk cell_11913 ( .C (clk), .D (signal_14458), .Q (signal_14459) ) ;
    buf_clk cell_11929 ( .C (clk), .D (signal_14474), .Q (signal_14475) ) ;
    buf_clk cell_11945 ( .C (clk), .D (signal_14490), .Q (signal_14491) ) ;
    buf_clk cell_11961 ( .C (clk), .D (signal_14506), .Q (signal_14507) ) ;
    buf_clk cell_11977 ( .C (clk), .D (signal_14522), .Q (signal_14523) ) ;
    buf_clk cell_11993 ( .C (clk), .D (signal_14538), .Q (signal_14539) ) ;
    buf_clk cell_12009 ( .C (clk), .D (signal_14554), .Q (signal_14555) ) ;
    buf_clk cell_12025 ( .C (clk), .D (signal_14570), .Q (signal_14571) ) ;
    buf_clk cell_12041 ( .C (clk), .D (signal_14586), .Q (signal_14587) ) ;
    buf_clk cell_12057 ( .C (clk), .D (signal_14602), .Q (signal_14603) ) ;
    buf_clk cell_12073 ( .C (clk), .D (signal_14618), .Q (signal_14619) ) ;
    buf_clk cell_12089 ( .C (clk), .D (signal_14634), .Q (signal_14635) ) ;
    buf_clk cell_12105 ( .C (clk), .D (signal_14650), .Q (signal_14651) ) ;
    buf_clk cell_12121 ( .C (clk), .D (signal_14666), .Q (signal_14667) ) ;
    buf_clk cell_12137 ( .C (clk), .D (signal_14682), .Q (signal_14683) ) ;
    buf_clk cell_12153 ( .C (clk), .D (signal_14698), .Q (signal_14699) ) ;
    buf_clk cell_12169 ( .C (clk), .D (signal_14714), .Q (signal_14715) ) ;
    buf_clk cell_12185 ( .C (clk), .D (signal_14730), .Q (signal_14731) ) ;
    buf_clk cell_12201 ( .C (clk), .D (signal_14746), .Q (signal_14747) ) ;
    buf_clk cell_12217 ( .C (clk), .D (signal_14762), .Q (signal_14763) ) ;
    buf_clk cell_12233 ( .C (clk), .D (signal_14778), .Q (signal_14779) ) ;
    buf_clk cell_12249 ( .C (clk), .D (signal_14794), .Q (signal_14795) ) ;
    buf_clk cell_12265 ( .C (clk), .D (signal_14810), .Q (signal_14811) ) ;
    buf_clk cell_12281 ( .C (clk), .D (signal_14826), .Q (signal_14827) ) ;
    buf_clk cell_12297 ( .C (clk), .D (signal_14842), .Q (signal_14843) ) ;
    buf_clk cell_12313 ( .C (clk), .D (signal_14858), .Q (signal_14859) ) ;
    buf_clk cell_12329 ( .C (clk), .D (signal_14874), .Q (signal_14875) ) ;
    buf_clk cell_12345 ( .C (clk), .D (signal_14890), .Q (signal_14891) ) ;
    buf_clk cell_12361 ( .C (clk), .D (signal_14906), .Q (signal_14907) ) ;
    buf_clk cell_12377 ( .C (clk), .D (signal_14922), .Q (signal_14923) ) ;
    buf_clk cell_12393 ( .C (clk), .D (signal_14938), .Q (signal_14939) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2121 ( .s ({signal_4930, signal_4918}), .b ({signal_4125, signal_2358}), .a ({signal_4124, signal_2357}), .clk (clk), .r (Fresh[407]), .c ({signal_4164, signal_2389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2122 ( .s ({signal_4930, signal_4918}), .b ({signal_4127, signal_2360}), .a ({signal_4126, signal_2359}), .clk (clk), .r (Fresh[408]), .c ({signal_4165, signal_2390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2123 ( .s ({signal_4930, signal_4918}), .b ({signal_4129, signal_2362}), .a ({signal_4128, signal_2361}), .clk (clk), .r (Fresh[409]), .c ({signal_4166, signal_2391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2124 ( .s ({signal_4930, signal_4918}), .b ({signal_4131, signal_2364}), .a ({signal_4130, signal_2363}), .clk (clk), .r (Fresh[410]), .c ({signal_4167, signal_2392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2125 ( .s ({signal_4930, signal_4918}), .b ({signal_4133, signal_2366}), .a ({signal_4132, signal_2365}), .clk (clk), .r (Fresh[411]), .c ({signal_4168, signal_2393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2126 ( .s ({signal_4930, signal_4918}), .b ({signal_4135, signal_2368}), .a ({signal_4134, signal_2367}), .clk (clk), .r (Fresh[412]), .c ({signal_4169, signal_2394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2127 ( .s ({signal_4930, signal_4918}), .b ({signal_4137, signal_2370}), .a ({signal_4136, signal_2369}), .clk (clk), .r (Fresh[413]), .c ({signal_4170, signal_2395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2128 ( .s ({signal_4930, signal_4918}), .b ({signal_4139, signal_2372}), .a ({signal_4138, signal_2371}), .clk (clk), .r (Fresh[414]), .c ({signal_4171, signal_2396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2129 ( .s ({signal_4930, signal_4918}), .b ({signal_4141, signal_2374}), .a ({signal_4140, signal_2373}), .clk (clk), .r (Fresh[415]), .c ({signal_4172, signal_2397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2130 ( .s ({signal_4930, signal_4918}), .b ({signal_4143, signal_2376}), .a ({signal_4142, signal_2375}), .clk (clk), .r (Fresh[416]), .c ({signal_4173, signal_2398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2131 ( .s ({signal_4930, signal_4918}), .b ({signal_4145, signal_2378}), .a ({signal_4144, signal_2377}), .clk (clk), .r (Fresh[417]), .c ({signal_4174, signal_2399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2132 ( .s ({signal_4930, signal_4918}), .b ({signal_4147, signal_2380}), .a ({signal_4146, signal_2379}), .clk (clk), .r (Fresh[418]), .c ({signal_4175, signal_2400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2133 ( .s ({signal_4930, signal_4918}), .b ({signal_4149, signal_2382}), .a ({signal_4148, signal_2381}), .clk (clk), .r (Fresh[419]), .c ({signal_4176, signal_2401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2134 ( .s ({signal_4930, signal_4918}), .b ({signal_4151, signal_2384}), .a ({signal_4150, signal_2383}), .clk (clk), .r (Fresh[420]), .c ({signal_4177, signal_2402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2135 ( .s ({signal_4930, signal_4918}), .b ({signal_4153, signal_2386}), .a ({signal_4152, signal_2385}), .clk (clk), .r (Fresh[421]), .c ({signal_4178, signal_2403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2136 ( .s ({signal_4930, signal_4918}), .b ({signal_4155, signal_2388}), .a ({signal_4154, signal_2387}), .clk (clk), .r (Fresh[422]), .c ({signal_4179, signal_2404}) ) ;
    buf_clk cell_2398 ( .C (clk), .D (signal_4943), .Q (signal_4944) ) ;
    buf_clk cell_2414 ( .C (clk), .D (signal_4959), .Q (signal_4960) ) ;
    buf_clk cell_2430 ( .C (clk), .D (signal_4975), .Q (signal_4976) ) ;
    buf_clk cell_2446 ( .C (clk), .D (signal_4991), .Q (signal_4992) ) ;
    buf_clk cell_2462 ( .C (clk), .D (signal_5007), .Q (signal_5008) ) ;
    buf_clk cell_2478 ( .C (clk), .D (signal_5023), .Q (signal_5024) ) ;
    buf_clk cell_2494 ( .C (clk), .D (signal_5039), .Q (signal_5040) ) ;
    buf_clk cell_2510 ( .C (clk), .D (signal_5055), .Q (signal_5056) ) ;
    buf_clk cell_2526 ( .C (clk), .D (signal_5071), .Q (signal_5072) ) ;
    buf_clk cell_2542 ( .C (clk), .D (signal_5087), .Q (signal_5088) ) ;
    buf_clk cell_2558 ( .C (clk), .D (signal_5103), .Q (signal_5104) ) ;
    buf_clk cell_2574 ( .C (clk), .D (signal_5119), .Q (signal_5120) ) ;
    buf_clk cell_2590 ( .C (clk), .D (signal_5135), .Q (signal_5136) ) ;
    buf_clk cell_2606 ( .C (clk), .D (signal_5151), .Q (signal_5152) ) ;
    buf_clk cell_2622 ( .C (clk), .D (signal_5167), .Q (signal_5168) ) ;
    buf_clk cell_2638 ( .C (clk), .D (signal_5183), .Q (signal_5184) ) ;
    buf_clk cell_2654 ( .C (clk), .D (signal_5199), .Q (signal_5200) ) ;
    buf_clk cell_2670 ( .C (clk), .D (signal_5215), .Q (signal_5216) ) ;
    buf_clk cell_2686 ( .C (clk), .D (signal_5231), .Q (signal_5232) ) ;
    buf_clk cell_2702 ( .C (clk), .D (signal_5247), .Q (signal_5248) ) ;
    buf_clk cell_2718 ( .C (clk), .D (signal_5263), .Q (signal_5264) ) ;
    buf_clk cell_2734 ( .C (clk), .D (signal_5279), .Q (signal_5280) ) ;
    buf_clk cell_2750 ( .C (clk), .D (signal_5295), .Q (signal_5296) ) ;
    buf_clk cell_2766 ( .C (clk), .D (signal_5311), .Q (signal_5312) ) ;
    buf_clk cell_2782 ( .C (clk), .D (signal_5327), .Q (signal_5328) ) ;
    buf_clk cell_2798 ( .C (clk), .D (signal_5343), .Q (signal_5344) ) ;
    buf_clk cell_2814 ( .C (clk), .D (signal_5359), .Q (signal_5360) ) ;
    buf_clk cell_2830 ( .C (clk), .D (signal_5375), .Q (signal_5376) ) ;
    buf_clk cell_2846 ( .C (clk), .D (signal_5391), .Q (signal_5392) ) ;
    buf_clk cell_2862 ( .C (clk), .D (signal_5407), .Q (signal_5408) ) ;
    buf_clk cell_2878 ( .C (clk), .D (signal_5423), .Q (signal_5424) ) ;
    buf_clk cell_2894 ( .C (clk), .D (signal_5439), .Q (signal_5440) ) ;
    buf_clk cell_2910 ( .C (clk), .D (signal_5455), .Q (signal_5456) ) ;
    buf_clk cell_2926 ( .C (clk), .D (signal_5471), .Q (signal_5472) ) ;
    buf_clk cell_2942 ( .C (clk), .D (signal_5487), .Q (signal_5488) ) ;
    buf_clk cell_2958 ( .C (clk), .D (signal_5503), .Q (signal_5504) ) ;
    buf_clk cell_2974 ( .C (clk), .D (signal_5519), .Q (signal_5520) ) ;
    buf_clk cell_2990 ( .C (clk), .D (signal_5535), .Q (signal_5536) ) ;
    buf_clk cell_3006 ( .C (clk), .D (signal_5551), .Q (signal_5552) ) ;
    buf_clk cell_3022 ( .C (clk), .D (signal_5567), .Q (signal_5568) ) ;
    buf_clk cell_3038 ( .C (clk), .D (signal_5583), .Q (signal_5584) ) ;
    buf_clk cell_3054 ( .C (clk), .D (signal_5599), .Q (signal_5600) ) ;
    buf_clk cell_3070 ( .C (clk), .D (signal_5615), .Q (signal_5616) ) ;
    buf_clk cell_3086 ( .C (clk), .D (signal_5631), .Q (signal_5632) ) ;
    buf_clk cell_3102 ( .C (clk), .D (signal_5647), .Q (signal_5648) ) ;
    buf_clk cell_3118 ( .C (clk), .D (signal_5663), .Q (signal_5664) ) ;
    buf_clk cell_3134 ( .C (clk), .D (signal_5679), .Q (signal_5680) ) ;
    buf_clk cell_3150 ( .C (clk), .D (signal_5695), .Q (signal_5696) ) ;
    buf_clk cell_3166 ( .C (clk), .D (signal_5711), .Q (signal_5712) ) ;
    buf_clk cell_3182 ( .C (clk), .D (signal_5727), .Q (signal_5728) ) ;
    buf_clk cell_3198 ( .C (clk), .D (signal_5743), .Q (signal_5744) ) ;
    buf_clk cell_3214 ( .C (clk), .D (signal_5759), .Q (signal_5760) ) ;
    buf_clk cell_3230 ( .C (clk), .D (signal_5775), .Q (signal_5776) ) ;
    buf_clk cell_3246 ( .C (clk), .D (signal_5791), .Q (signal_5792) ) ;
    buf_clk cell_3262 ( .C (clk), .D (signal_5807), .Q (signal_5808) ) ;
    buf_clk cell_3278 ( .C (clk), .D (signal_5823), .Q (signal_5824) ) ;
    buf_clk cell_3294 ( .C (clk), .D (signal_5839), .Q (signal_5840) ) ;
    buf_clk cell_3310 ( .C (clk), .D (signal_5855), .Q (signal_5856) ) ;
    buf_clk cell_3326 ( .C (clk), .D (signal_5871), .Q (signal_5872) ) ;
    buf_clk cell_3342 ( .C (clk), .D (signal_5887), .Q (signal_5888) ) ;
    buf_clk cell_3358 ( .C (clk), .D (signal_5903), .Q (signal_5904) ) ;
    buf_clk cell_3374 ( .C (clk), .D (signal_5919), .Q (signal_5920) ) ;
    buf_clk cell_3390 ( .C (clk), .D (signal_5935), .Q (signal_5936) ) ;
    buf_clk cell_3406 ( .C (clk), .D (signal_5951), .Q (signal_5952) ) ;
    buf_clk cell_3422 ( .C (clk), .D (signal_5967), .Q (signal_5968) ) ;
    buf_clk cell_3438 ( .C (clk), .D (signal_5983), .Q (signal_5984) ) ;
    buf_clk cell_3454 ( .C (clk), .D (signal_5999), .Q (signal_6000) ) ;
    buf_clk cell_3470 ( .C (clk), .D (signal_6015), .Q (signal_6016) ) ;
    buf_clk cell_3486 ( .C (clk), .D (signal_6031), .Q (signal_6032) ) ;
    buf_clk cell_3502 ( .C (clk), .D (signal_6047), .Q (signal_6048) ) ;
    buf_clk cell_3518 ( .C (clk), .D (signal_6063), .Q (signal_6064) ) ;
    buf_clk cell_3534 ( .C (clk), .D (signal_6079), .Q (signal_6080) ) ;
    buf_clk cell_3550 ( .C (clk), .D (signal_6095), .Q (signal_6096) ) ;
    buf_clk cell_3566 ( .C (clk), .D (signal_6111), .Q (signal_6112) ) ;
    buf_clk cell_3582 ( .C (clk), .D (signal_6127), .Q (signal_6128) ) ;
    buf_clk cell_3598 ( .C (clk), .D (signal_6143), .Q (signal_6144) ) ;
    buf_clk cell_3614 ( .C (clk), .D (signal_6159), .Q (signal_6160) ) ;
    buf_clk cell_3630 ( .C (clk), .D (signal_6175), .Q (signal_6176) ) ;
    buf_clk cell_3646 ( .C (clk), .D (signal_6191), .Q (signal_6192) ) ;
    buf_clk cell_3662 ( .C (clk), .D (signal_6207), .Q (signal_6208) ) ;
    buf_clk cell_3678 ( .C (clk), .D (signal_6223), .Q (signal_6224) ) ;
    buf_clk cell_3694 ( .C (clk), .D (signal_6239), .Q (signal_6240) ) ;
    buf_clk cell_3710 ( .C (clk), .D (signal_6255), .Q (signal_6256) ) ;
    buf_clk cell_3726 ( .C (clk), .D (signal_6271), .Q (signal_6272) ) ;
    buf_clk cell_3742 ( .C (clk), .D (signal_6287), .Q (signal_6288) ) ;
    buf_clk cell_3758 ( .C (clk), .D (signal_6303), .Q (signal_6304) ) ;
    buf_clk cell_3774 ( .C (clk), .D (signal_6319), .Q (signal_6320) ) ;
    buf_clk cell_3790 ( .C (clk), .D (signal_6335), .Q (signal_6336) ) ;
    buf_clk cell_3806 ( .C (clk), .D (signal_6351), .Q (signal_6352) ) ;
    buf_clk cell_3822 ( .C (clk), .D (signal_6367), .Q (signal_6368) ) ;
    buf_clk cell_3838 ( .C (clk), .D (signal_6383), .Q (signal_6384) ) ;
    buf_clk cell_3854 ( .C (clk), .D (signal_6399), .Q (signal_6400) ) ;
    buf_clk cell_3870 ( .C (clk), .D (signal_6415), .Q (signal_6416) ) ;
    buf_clk cell_3886 ( .C (clk), .D (signal_6431), .Q (signal_6432) ) ;
    buf_clk cell_3902 ( .C (clk), .D (signal_6447), .Q (signal_6448) ) ;
    buf_clk cell_3918 ( .C (clk), .D (signal_6463), .Q (signal_6464) ) ;
    buf_clk cell_3934 ( .C (clk), .D (signal_6479), .Q (signal_6480) ) ;
    buf_clk cell_3950 ( .C (clk), .D (signal_6495), .Q (signal_6496) ) ;
    buf_clk cell_3966 ( .C (clk), .D (signal_6511), .Q (signal_6512) ) ;
    buf_clk cell_3982 ( .C (clk), .D (signal_6527), .Q (signal_6528) ) ;
    buf_clk cell_3998 ( .C (clk), .D (signal_6543), .Q (signal_6544) ) ;
    buf_clk cell_4014 ( .C (clk), .D (signal_6559), .Q (signal_6560) ) ;
    buf_clk cell_4030 ( .C (clk), .D (signal_6575), .Q (signal_6576) ) ;
    buf_clk cell_4046 ( .C (clk), .D (signal_6591), .Q (signal_6592) ) ;
    buf_clk cell_4062 ( .C (clk), .D (signal_6607), .Q (signal_6608) ) ;
    buf_clk cell_4078 ( .C (clk), .D (signal_6623), .Q (signal_6624) ) ;
    buf_clk cell_4094 ( .C (clk), .D (signal_6639), .Q (signal_6640) ) ;
    buf_clk cell_4110 ( .C (clk), .D (signal_6655), .Q (signal_6656) ) ;
    buf_clk cell_4126 ( .C (clk), .D (signal_6671), .Q (signal_6672) ) ;
    buf_clk cell_4142 ( .C (clk), .D (signal_6687), .Q (signal_6688) ) ;
    buf_clk cell_4158 ( .C (clk), .D (signal_6703), .Q (signal_6704) ) ;
    buf_clk cell_4174 ( .C (clk), .D (signal_6719), .Q (signal_6720) ) ;
    buf_clk cell_4190 ( .C (clk), .D (signal_6735), .Q (signal_6736) ) ;
    buf_clk cell_4206 ( .C (clk), .D (signal_6751), .Q (signal_6752) ) ;
    buf_clk cell_4222 ( .C (clk), .D (signal_6767), .Q (signal_6768) ) ;
    buf_clk cell_4238 ( .C (clk), .D (signal_6783), .Q (signal_6784) ) ;
    buf_clk cell_4254 ( .C (clk), .D (signal_6799), .Q (signal_6800) ) ;
    buf_clk cell_4270 ( .C (clk), .D (signal_6815), .Q (signal_6816) ) ;
    buf_clk cell_4286 ( .C (clk), .D (signal_6831), .Q (signal_6832) ) ;
    buf_clk cell_4302 ( .C (clk), .D (signal_6847), .Q (signal_6848) ) ;
    buf_clk cell_4318 ( .C (clk), .D (signal_6863), .Q (signal_6864) ) ;
    buf_clk cell_4334 ( .C (clk), .D (signal_6879), .Q (signal_6880) ) ;
    buf_clk cell_4350 ( .C (clk), .D (signal_6895), .Q (signal_6896) ) ;
    buf_clk cell_4366 ( .C (clk), .D (signal_6911), .Q (signal_6912) ) ;
    buf_clk cell_4382 ( .C (clk), .D (signal_6927), .Q (signal_6928) ) ;
    buf_clk cell_4398 ( .C (clk), .D (signal_6943), .Q (signal_6944) ) ;
    buf_clk cell_4414 ( .C (clk), .D (signal_6959), .Q (signal_6960) ) ;
    buf_clk cell_4428 ( .C (clk), .D (signal_6973), .Q (signal_6974) ) ;
    buf_clk cell_4442 ( .C (clk), .D (signal_6987), .Q (signal_6988) ) ;
    buf_clk cell_4458 ( .C (clk), .D (signal_7003), .Q (signal_7004) ) ;
    buf_clk cell_4474 ( .C (clk), .D (signal_7019), .Q (signal_7020) ) ;
    buf_clk cell_4490 ( .C (clk), .D (signal_7035), .Q (signal_7036) ) ;
    buf_clk cell_4506 ( .C (clk), .D (signal_7051), .Q (signal_7052) ) ;
    buf_clk cell_4522 ( .C (clk), .D (signal_7067), .Q (signal_7068) ) ;
    buf_clk cell_4538 ( .C (clk), .D (signal_7083), .Q (signal_7084) ) ;
    buf_clk cell_4554 ( .C (clk), .D (signal_7099), .Q (signal_7100) ) ;
    buf_clk cell_4570 ( .C (clk), .D (signal_7115), .Q (signal_7116) ) ;
    buf_clk cell_4586 ( .C (clk), .D (signal_7131), .Q (signal_7132) ) ;
    buf_clk cell_4602 ( .C (clk), .D (signal_7147), .Q (signal_7148) ) ;
    buf_clk cell_4618 ( .C (clk), .D (signal_7163), .Q (signal_7164) ) ;
    buf_clk cell_4634 ( .C (clk), .D (signal_7179), .Q (signal_7180) ) ;
    buf_clk cell_4650 ( .C (clk), .D (signal_7195), .Q (signal_7196) ) ;
    buf_clk cell_4666 ( .C (clk), .D (signal_7211), .Q (signal_7212) ) ;
    buf_clk cell_4682 ( .C (clk), .D (signal_7227), .Q (signal_7228) ) ;
    buf_clk cell_4698 ( .C (clk), .D (signal_7243), .Q (signal_7244) ) ;
    buf_clk cell_4714 ( .C (clk), .D (signal_7259), .Q (signal_7260) ) ;
    buf_clk cell_4730 ( .C (clk), .D (signal_7275), .Q (signal_7276) ) ;
    buf_clk cell_4746 ( .C (clk), .D (signal_7291), .Q (signal_7292) ) ;
    buf_clk cell_4762 ( .C (clk), .D (signal_7307), .Q (signal_7308) ) ;
    buf_clk cell_4778 ( .C (clk), .D (signal_7323), .Q (signal_7324) ) ;
    buf_clk cell_4794 ( .C (clk), .D (signal_7339), .Q (signal_7340) ) ;
    buf_clk cell_4810 ( .C (clk), .D (signal_7355), .Q (signal_7356) ) ;
    buf_clk cell_4826 ( .C (clk), .D (signal_7371), .Q (signal_7372) ) ;
    buf_clk cell_4842 ( .C (clk), .D (signal_7387), .Q (signal_7388) ) ;
    buf_clk cell_4858 ( .C (clk), .D (signal_7403), .Q (signal_7404) ) ;
    buf_clk cell_4874 ( .C (clk), .D (signal_7419), .Q (signal_7420) ) ;
    buf_clk cell_4890 ( .C (clk), .D (signal_7435), .Q (signal_7436) ) ;
    buf_clk cell_4906 ( .C (clk), .D (signal_7451), .Q (signal_7452) ) ;
    buf_clk cell_4922 ( .C (clk), .D (signal_7467), .Q (signal_7468) ) ;
    buf_clk cell_4938 ( .C (clk), .D (signal_7483), .Q (signal_7484) ) ;
    buf_clk cell_4954 ( .C (clk), .D (signal_7499), .Q (signal_7500) ) ;
    buf_clk cell_4970 ( .C (clk), .D (signal_7515), .Q (signal_7516) ) ;
    buf_clk cell_4986 ( .C (clk), .D (signal_7531), .Q (signal_7532) ) ;
    buf_clk cell_5002 ( .C (clk), .D (signal_7547), .Q (signal_7548) ) ;
    buf_clk cell_5018 ( .C (clk), .D (signal_7563), .Q (signal_7564) ) ;
    buf_clk cell_5034 ( .C (clk), .D (signal_7579), .Q (signal_7580) ) ;
    buf_clk cell_5050 ( .C (clk), .D (signal_7595), .Q (signal_7596) ) ;
    buf_clk cell_5066 ( .C (clk), .D (signal_7611), .Q (signal_7612) ) ;
    buf_clk cell_5082 ( .C (clk), .D (signal_7627), .Q (signal_7628) ) ;
    buf_clk cell_5098 ( .C (clk), .D (signal_7643), .Q (signal_7644) ) ;
    buf_clk cell_5114 ( .C (clk), .D (signal_7659), .Q (signal_7660) ) ;
    buf_clk cell_5130 ( .C (clk), .D (signal_7675), .Q (signal_7676) ) ;
    buf_clk cell_5146 ( .C (clk), .D (signal_7691), .Q (signal_7692) ) ;
    buf_clk cell_5162 ( .C (clk), .D (signal_7707), .Q (signal_7708) ) ;
    buf_clk cell_5178 ( .C (clk), .D (signal_7723), .Q (signal_7724) ) ;
    buf_clk cell_5194 ( .C (clk), .D (signal_7739), .Q (signal_7740) ) ;
    buf_clk cell_5210 ( .C (clk), .D (signal_7755), .Q (signal_7756) ) ;
    buf_clk cell_5226 ( .C (clk), .D (signal_7771), .Q (signal_7772) ) ;
    buf_clk cell_5242 ( .C (clk), .D (signal_7787), .Q (signal_7788) ) ;
    buf_clk cell_5258 ( .C (clk), .D (signal_7803), .Q (signal_7804) ) ;
    buf_clk cell_5274 ( .C (clk), .D (signal_7819), .Q (signal_7820) ) ;
    buf_clk cell_5290 ( .C (clk), .D (signal_7835), .Q (signal_7836) ) ;
    buf_clk cell_5306 ( .C (clk), .D (signal_7851), .Q (signal_7852) ) ;
    buf_clk cell_5322 ( .C (clk), .D (signal_7867), .Q (signal_7868) ) ;
    buf_clk cell_5338 ( .C (clk), .D (signal_7883), .Q (signal_7884) ) ;
    buf_clk cell_5354 ( .C (clk), .D (signal_7899), .Q (signal_7900) ) ;
    buf_clk cell_5370 ( .C (clk), .D (signal_7915), .Q (signal_7916) ) ;
    buf_clk cell_5386 ( .C (clk), .D (signal_7931), .Q (signal_7932) ) ;
    buf_clk cell_5402 ( .C (clk), .D (signal_7947), .Q (signal_7948) ) ;
    buf_clk cell_5418 ( .C (clk), .D (signal_7963), .Q (signal_7964) ) ;
    buf_clk cell_5434 ( .C (clk), .D (signal_7979), .Q (signal_7980) ) ;
    buf_clk cell_5450 ( .C (clk), .D (signal_7995), .Q (signal_7996) ) ;
    buf_clk cell_5466 ( .C (clk), .D (signal_8011), .Q (signal_8012) ) ;
    buf_clk cell_5482 ( .C (clk), .D (signal_8027), .Q (signal_8028) ) ;
    buf_clk cell_5498 ( .C (clk), .D (signal_8043), .Q (signal_8044) ) ;
    buf_clk cell_5514 ( .C (clk), .D (signal_8059), .Q (signal_8060) ) ;
    buf_clk cell_5530 ( .C (clk), .D (signal_8075), .Q (signal_8076) ) ;
    buf_clk cell_5546 ( .C (clk), .D (signal_8091), .Q (signal_8092) ) ;
    buf_clk cell_5562 ( .C (clk), .D (signal_8107), .Q (signal_8108) ) ;
    buf_clk cell_5578 ( .C (clk), .D (signal_8123), .Q (signal_8124) ) ;
    buf_clk cell_5594 ( .C (clk), .D (signal_8139), .Q (signal_8140) ) ;
    buf_clk cell_5610 ( .C (clk), .D (signal_8155), .Q (signal_8156) ) ;
    buf_clk cell_5626 ( .C (clk), .D (signal_8171), .Q (signal_8172) ) ;
    buf_clk cell_5642 ( .C (clk), .D (signal_8187), .Q (signal_8188) ) ;
    buf_clk cell_5658 ( .C (clk), .D (signal_8203), .Q (signal_8204) ) ;
    buf_clk cell_5674 ( .C (clk), .D (signal_8219), .Q (signal_8220) ) ;
    buf_clk cell_5690 ( .C (clk), .D (signal_8235), .Q (signal_8236) ) ;
    buf_clk cell_5706 ( .C (clk), .D (signal_8251), .Q (signal_8252) ) ;
    buf_clk cell_5722 ( .C (clk), .D (signal_8267), .Q (signal_8268) ) ;
    buf_clk cell_5738 ( .C (clk), .D (signal_8283), .Q (signal_8284) ) ;
    buf_clk cell_5754 ( .C (clk), .D (signal_8299), .Q (signal_8300) ) ;
    buf_clk cell_5770 ( .C (clk), .D (signal_8315), .Q (signal_8316) ) ;
    buf_clk cell_5786 ( .C (clk), .D (signal_8331), .Q (signal_8332) ) ;
    buf_clk cell_5802 ( .C (clk), .D (signal_8347), .Q (signal_8348) ) ;
    buf_clk cell_5818 ( .C (clk), .D (signal_8363), .Q (signal_8364) ) ;
    buf_clk cell_5834 ( .C (clk), .D (signal_8379), .Q (signal_8380) ) ;
    buf_clk cell_5850 ( .C (clk), .D (signal_8395), .Q (signal_8396) ) ;
    buf_clk cell_5866 ( .C (clk), .D (signal_8411), .Q (signal_8412) ) ;
    buf_clk cell_5882 ( .C (clk), .D (signal_8427), .Q (signal_8428) ) ;
    buf_clk cell_5898 ( .C (clk), .D (signal_8443), .Q (signal_8444) ) ;
    buf_clk cell_5914 ( .C (clk), .D (signal_8459), .Q (signal_8460) ) ;
    buf_clk cell_5930 ( .C (clk), .D (signal_8475), .Q (signal_8476) ) ;
    buf_clk cell_5946 ( .C (clk), .D (signal_8491), .Q (signal_8492) ) ;
    buf_clk cell_5962 ( .C (clk), .D (signal_8507), .Q (signal_8508) ) ;
    buf_clk cell_5978 ( .C (clk), .D (signal_8523), .Q (signal_8524) ) ;
    buf_clk cell_5994 ( .C (clk), .D (signal_8539), .Q (signal_8540) ) ;
    buf_clk cell_6010 ( .C (clk), .D (signal_8555), .Q (signal_8556) ) ;
    buf_clk cell_6026 ( .C (clk), .D (signal_8571), .Q (signal_8572) ) ;
    buf_clk cell_6042 ( .C (clk), .D (signal_8587), .Q (signal_8588) ) ;
    buf_clk cell_6058 ( .C (clk), .D (signal_8603), .Q (signal_8604) ) ;
    buf_clk cell_6074 ( .C (clk), .D (signal_8619), .Q (signal_8620) ) ;
    buf_clk cell_6090 ( .C (clk), .D (signal_8635), .Q (signal_8636) ) ;
    buf_clk cell_6106 ( .C (clk), .D (signal_8651), .Q (signal_8652) ) ;
    buf_clk cell_6122 ( .C (clk), .D (signal_8667), .Q (signal_8668) ) ;
    buf_clk cell_6138 ( .C (clk), .D (signal_8683), .Q (signal_8684) ) ;
    buf_clk cell_6154 ( .C (clk), .D (signal_8699), .Q (signal_8700) ) ;
    buf_clk cell_6170 ( .C (clk), .D (signal_8715), .Q (signal_8716) ) ;
    buf_clk cell_6186 ( .C (clk), .D (signal_8731), .Q (signal_8732) ) ;
    buf_clk cell_6202 ( .C (clk), .D (signal_8747), .Q (signal_8748) ) ;
    buf_clk cell_6218 ( .C (clk), .D (signal_8763), .Q (signal_8764) ) ;
    buf_clk cell_6234 ( .C (clk), .D (signal_8779), .Q (signal_8780) ) ;
    buf_clk cell_6250 ( .C (clk), .D (signal_8795), .Q (signal_8796) ) ;
    buf_clk cell_6266 ( .C (clk), .D (signal_8811), .Q (signal_8812) ) ;
    buf_clk cell_6282 ( .C (clk), .D (signal_8827), .Q (signal_8828) ) ;
    buf_clk cell_6298 ( .C (clk), .D (signal_8843), .Q (signal_8844) ) ;
    buf_clk cell_6314 ( .C (clk), .D (signal_8859), .Q (signal_8860) ) ;
    buf_clk cell_6330 ( .C (clk), .D (signal_8875), .Q (signal_8876) ) ;
    buf_clk cell_6346 ( .C (clk), .D (signal_8891), .Q (signal_8892) ) ;
    buf_clk cell_6362 ( .C (clk), .D (signal_8907), .Q (signal_8908) ) ;
    buf_clk cell_6378 ( .C (clk), .D (signal_8923), .Q (signal_8924) ) ;
    buf_clk cell_6394 ( .C (clk), .D (signal_8939), .Q (signal_8940) ) ;
    buf_clk cell_6410 ( .C (clk), .D (signal_8955), .Q (signal_8956) ) ;
    buf_clk cell_6426 ( .C (clk), .D (signal_8971), .Q (signal_8972) ) ;
    buf_clk cell_6442 ( .C (clk), .D (signal_8987), .Q (signal_8988) ) ;
    buf_clk cell_6458 ( .C (clk), .D (signal_9003), .Q (signal_9004) ) ;
    buf_clk cell_6474 ( .C (clk), .D (signal_9019), .Q (signal_9020) ) ;
    buf_clk cell_6490 ( .C (clk), .D (signal_9035), .Q (signal_9036) ) ;
    buf_clk cell_6506 ( .C (clk), .D (signal_9051), .Q (signal_9052) ) ;
    buf_clk cell_6522 ( .C (clk), .D (signal_9067), .Q (signal_9068) ) ;
    buf_clk cell_6538 ( .C (clk), .D (signal_9083), .Q (signal_9084) ) ;
    buf_clk cell_6554 ( .C (clk), .D (signal_9099), .Q (signal_9100) ) ;
    buf_clk cell_6570 ( .C (clk), .D (signal_9115), .Q (signal_9116) ) ;
    buf_clk cell_6586 ( .C (clk), .D (signal_9131), .Q (signal_9132) ) ;
    buf_clk cell_6602 ( .C (clk), .D (signal_9147), .Q (signal_9148) ) ;
    buf_clk cell_6618 ( .C (clk), .D (signal_9163), .Q (signal_9164) ) ;
    buf_clk cell_6634 ( .C (clk), .D (signal_9179), .Q (signal_9180) ) ;
    buf_clk cell_6650 ( .C (clk), .D (signal_9195), .Q (signal_9196) ) ;
    buf_clk cell_6666 ( .C (clk), .D (signal_9211), .Q (signal_9212) ) ;
    buf_clk cell_6682 ( .C (clk), .D (signal_9227), .Q (signal_9228) ) ;
    buf_clk cell_6698 ( .C (clk), .D (signal_9243), .Q (signal_9244) ) ;
    buf_clk cell_6714 ( .C (clk), .D (signal_9259), .Q (signal_9260) ) ;
    buf_clk cell_6730 ( .C (clk), .D (signal_9275), .Q (signal_9276) ) ;
    buf_clk cell_6746 ( .C (clk), .D (signal_9291), .Q (signal_9292) ) ;
    buf_clk cell_6762 ( .C (clk), .D (signal_9307), .Q (signal_9308) ) ;
    buf_clk cell_6778 ( .C (clk), .D (signal_9323), .Q (signal_9324) ) ;
    buf_clk cell_6794 ( .C (clk), .D (signal_9339), .Q (signal_9340) ) ;
    buf_clk cell_6810 ( .C (clk), .D (signal_9355), .Q (signal_9356) ) ;
    buf_clk cell_6826 ( .C (clk), .D (signal_9371), .Q (signal_9372) ) ;
    buf_clk cell_6842 ( .C (clk), .D (signal_9387), .Q (signal_9388) ) ;
    buf_clk cell_6858 ( .C (clk), .D (signal_9403), .Q (signal_9404) ) ;
    buf_clk cell_6874 ( .C (clk), .D (signal_9419), .Q (signal_9420) ) ;
    buf_clk cell_6890 ( .C (clk), .D (signal_9435), .Q (signal_9436) ) ;
    buf_clk cell_6906 ( .C (clk), .D (signal_9451), .Q (signal_9452) ) ;
    buf_clk cell_6922 ( .C (clk), .D (signal_9467), .Q (signal_9468) ) ;
    buf_clk cell_6938 ( .C (clk), .D (signal_9483), .Q (signal_9484) ) ;
    buf_clk cell_6954 ( .C (clk), .D (signal_9499), .Q (signal_9500) ) ;
    buf_clk cell_6970 ( .C (clk), .D (signal_9515), .Q (signal_9516) ) ;
    buf_clk cell_6986 ( .C (clk), .D (signal_9531), .Q (signal_9532) ) ;
    buf_clk cell_7002 ( .C (clk), .D (signal_9547), .Q (signal_9548) ) ;
    buf_clk cell_7018 ( .C (clk), .D (signal_9563), .Q (signal_9564) ) ;
    buf_clk cell_7034 ( .C (clk), .D (signal_9579), .Q (signal_9580) ) ;
    buf_clk cell_7050 ( .C (clk), .D (signal_9595), .Q (signal_9596) ) ;
    buf_clk cell_7066 ( .C (clk), .D (signal_9611), .Q (signal_9612) ) ;
    buf_clk cell_7082 ( .C (clk), .D (signal_9627), .Q (signal_9628) ) ;
    buf_clk cell_7098 ( .C (clk), .D (signal_9643), .Q (signal_9644) ) ;
    buf_clk cell_7114 ( .C (clk), .D (signal_9659), .Q (signal_9660) ) ;
    buf_clk cell_7130 ( .C (clk), .D (signal_9675), .Q (signal_9676) ) ;
    buf_clk cell_7146 ( .C (clk), .D (signal_9691), .Q (signal_9692) ) ;
    buf_clk cell_7162 ( .C (clk), .D (signal_9707), .Q (signal_9708) ) ;
    buf_clk cell_7178 ( .C (clk), .D (signal_9723), .Q (signal_9724) ) ;
    buf_clk cell_7194 ( .C (clk), .D (signal_9739), .Q (signal_9740) ) ;
    buf_clk cell_7210 ( .C (clk), .D (signal_9755), .Q (signal_9756) ) ;
    buf_clk cell_7226 ( .C (clk), .D (signal_9771), .Q (signal_9772) ) ;
    buf_clk cell_7242 ( .C (clk), .D (signal_9787), .Q (signal_9788) ) ;
    buf_clk cell_7258 ( .C (clk), .D (signal_9803), .Q (signal_9804) ) ;
    buf_clk cell_7274 ( .C (clk), .D (signal_9819), .Q (signal_9820) ) ;
    buf_clk cell_7290 ( .C (clk), .D (signal_9835), .Q (signal_9836) ) ;
    buf_clk cell_7306 ( .C (clk), .D (signal_9851), .Q (signal_9852) ) ;
    buf_clk cell_7322 ( .C (clk), .D (signal_9867), .Q (signal_9868) ) ;
    buf_clk cell_7338 ( .C (clk), .D (signal_9883), .Q (signal_9884) ) ;
    buf_clk cell_7354 ( .C (clk), .D (signal_9899), .Q (signal_9900) ) ;
    buf_clk cell_7370 ( .C (clk), .D (signal_9915), .Q (signal_9916) ) ;
    buf_clk cell_7386 ( .C (clk), .D (signal_9931), .Q (signal_9932) ) ;
    buf_clk cell_7402 ( .C (clk), .D (signal_9947), .Q (signal_9948) ) ;
    buf_clk cell_7418 ( .C (clk), .D (signal_9963), .Q (signal_9964) ) ;
    buf_clk cell_7434 ( .C (clk), .D (signal_9979), .Q (signal_9980) ) ;
    buf_clk cell_7450 ( .C (clk), .D (signal_9995), .Q (signal_9996) ) ;
    buf_clk cell_7466 ( .C (clk), .D (signal_10011), .Q (signal_10012) ) ;
    buf_clk cell_7482 ( .C (clk), .D (signal_10027), .Q (signal_10028) ) ;
    buf_clk cell_7498 ( .C (clk), .D (signal_10043), .Q (signal_10044) ) ;
    buf_clk cell_7514 ( .C (clk), .D (signal_10059), .Q (signal_10060) ) ;
    buf_clk cell_7530 ( .C (clk), .D (signal_10075), .Q (signal_10076) ) ;
    buf_clk cell_7546 ( .C (clk), .D (signal_10091), .Q (signal_10092) ) ;
    buf_clk cell_7562 ( .C (clk), .D (signal_10107), .Q (signal_10108) ) ;
    buf_clk cell_7578 ( .C (clk), .D (signal_10123), .Q (signal_10124) ) ;
    buf_clk cell_7594 ( .C (clk), .D (signal_10139), .Q (signal_10140) ) ;
    buf_clk cell_7610 ( .C (clk), .D (signal_10155), .Q (signal_10156) ) ;
    buf_clk cell_7626 ( .C (clk), .D (signal_10171), .Q (signal_10172) ) ;
    buf_clk cell_7642 ( .C (clk), .D (signal_10187), .Q (signal_10188) ) ;
    buf_clk cell_7658 ( .C (clk), .D (signal_10203), .Q (signal_10204) ) ;
    buf_clk cell_7674 ( .C (clk), .D (signal_10219), .Q (signal_10220) ) ;
    buf_clk cell_7690 ( .C (clk), .D (signal_10235), .Q (signal_10236) ) ;
    buf_clk cell_7706 ( .C (clk), .D (signal_10251), .Q (signal_10252) ) ;
    buf_clk cell_7722 ( .C (clk), .D (signal_10267), .Q (signal_10268) ) ;
    buf_clk cell_7738 ( .C (clk), .D (signal_10283), .Q (signal_10284) ) ;
    buf_clk cell_7754 ( .C (clk), .D (signal_10299), .Q (signal_10300) ) ;
    buf_clk cell_7770 ( .C (clk), .D (signal_10315), .Q (signal_10316) ) ;
    buf_clk cell_7786 ( .C (clk), .D (signal_10331), .Q (signal_10332) ) ;
    buf_clk cell_7802 ( .C (clk), .D (signal_10347), .Q (signal_10348) ) ;
    buf_clk cell_7818 ( .C (clk), .D (signal_10363), .Q (signal_10364) ) ;
    buf_clk cell_7834 ( .C (clk), .D (signal_10379), .Q (signal_10380) ) ;
    buf_clk cell_7850 ( .C (clk), .D (signal_10395), .Q (signal_10396) ) ;
    buf_clk cell_7866 ( .C (clk), .D (signal_10411), .Q (signal_10412) ) ;
    buf_clk cell_7882 ( .C (clk), .D (signal_10427), .Q (signal_10428) ) ;
    buf_clk cell_7898 ( .C (clk), .D (signal_10443), .Q (signal_10444) ) ;
    buf_clk cell_7914 ( .C (clk), .D (signal_10459), .Q (signal_10460) ) ;
    buf_clk cell_7930 ( .C (clk), .D (signal_10475), .Q (signal_10476) ) ;
    buf_clk cell_7946 ( .C (clk), .D (signal_10491), .Q (signal_10492) ) ;
    buf_clk cell_7962 ( .C (clk), .D (signal_10507), .Q (signal_10508) ) ;
    buf_clk cell_7978 ( .C (clk), .D (signal_10523), .Q (signal_10524) ) ;
    buf_clk cell_7994 ( .C (clk), .D (signal_10539), .Q (signal_10540) ) ;
    buf_clk cell_8010 ( .C (clk), .D (signal_10555), .Q (signal_10556) ) ;
    buf_clk cell_8026 ( .C (clk), .D (signal_10571), .Q (signal_10572) ) ;
    buf_clk cell_8042 ( .C (clk), .D (signal_10587), .Q (signal_10588) ) ;
    buf_clk cell_8058 ( .C (clk), .D (signal_10603), .Q (signal_10604) ) ;
    buf_clk cell_8074 ( .C (clk), .D (signal_10619), .Q (signal_10620) ) ;
    buf_clk cell_8090 ( .C (clk), .D (signal_10635), .Q (signal_10636) ) ;
    buf_clk cell_8106 ( .C (clk), .D (signal_10651), .Q (signal_10652) ) ;
    buf_clk cell_8122 ( .C (clk), .D (signal_10667), .Q (signal_10668) ) ;
    buf_clk cell_8138 ( .C (clk), .D (signal_10683), .Q (signal_10684) ) ;
    buf_clk cell_8154 ( .C (clk), .D (signal_10699), .Q (signal_10700) ) ;
    buf_clk cell_8170 ( .C (clk), .D (signal_10715), .Q (signal_10716) ) ;
    buf_clk cell_8186 ( .C (clk), .D (signal_10731), .Q (signal_10732) ) ;
    buf_clk cell_8202 ( .C (clk), .D (signal_10747), .Q (signal_10748) ) ;
    buf_clk cell_8218 ( .C (clk), .D (signal_10763), .Q (signal_10764) ) ;
    buf_clk cell_8234 ( .C (clk), .D (signal_10779), .Q (signal_10780) ) ;
    buf_clk cell_8250 ( .C (clk), .D (signal_10795), .Q (signal_10796) ) ;
    buf_clk cell_8266 ( .C (clk), .D (signal_10811), .Q (signal_10812) ) ;
    buf_clk cell_8282 ( .C (clk), .D (signal_10827), .Q (signal_10828) ) ;
    buf_clk cell_8298 ( .C (clk), .D (signal_10843), .Q (signal_10844) ) ;
    buf_clk cell_8314 ( .C (clk), .D (signal_10859), .Q (signal_10860) ) ;
    buf_clk cell_8330 ( .C (clk), .D (signal_10875), .Q (signal_10876) ) ;
    buf_clk cell_8346 ( .C (clk), .D (signal_10891), .Q (signal_10892) ) ;
    buf_clk cell_8362 ( .C (clk), .D (signal_10907), .Q (signal_10908) ) ;
    buf_clk cell_8378 ( .C (clk), .D (signal_10923), .Q (signal_10924) ) ;
    buf_clk cell_8394 ( .C (clk), .D (signal_10939), .Q (signal_10940) ) ;
    buf_clk cell_8410 ( .C (clk), .D (signal_10955), .Q (signal_10956) ) ;
    buf_clk cell_8426 ( .C (clk), .D (signal_10971), .Q (signal_10972) ) ;
    buf_clk cell_8442 ( .C (clk), .D (signal_10987), .Q (signal_10988) ) ;
    buf_clk cell_8458 ( .C (clk), .D (signal_11003), .Q (signal_11004) ) ;
    buf_clk cell_8474 ( .C (clk), .D (signal_11019), .Q (signal_11020) ) ;
    buf_clk cell_8490 ( .C (clk), .D (signal_11035), .Q (signal_11036) ) ;
    buf_clk cell_8506 ( .C (clk), .D (signal_11051), .Q (signal_11052) ) ;
    buf_clk cell_8522 ( .C (clk), .D (signal_11067), .Q (signal_11068) ) ;
    buf_clk cell_8538 ( .C (clk), .D (signal_11083), .Q (signal_11084) ) ;
    buf_clk cell_8554 ( .C (clk), .D (signal_11099), .Q (signal_11100) ) ;
    buf_clk cell_8570 ( .C (clk), .D (signal_11115), .Q (signal_11116) ) ;
    buf_clk cell_8586 ( .C (clk), .D (signal_11131), .Q (signal_11132) ) ;
    buf_clk cell_8602 ( .C (clk), .D (signal_11147), .Q (signal_11148) ) ;
    buf_clk cell_8618 ( .C (clk), .D (signal_11163), .Q (signal_11164) ) ;
    buf_clk cell_8634 ( .C (clk), .D (signal_11179), .Q (signal_11180) ) ;
    buf_clk cell_8650 ( .C (clk), .D (signal_11195), .Q (signal_11196) ) ;
    buf_clk cell_8666 ( .C (clk), .D (signal_11211), .Q (signal_11212) ) ;
    buf_clk cell_8682 ( .C (clk), .D (signal_11227), .Q (signal_11228) ) ;
    buf_clk cell_8698 ( .C (clk), .D (signal_11243), .Q (signal_11244) ) ;
    buf_clk cell_8714 ( .C (clk), .D (signal_11259), .Q (signal_11260) ) ;
    buf_clk cell_8730 ( .C (clk), .D (signal_11275), .Q (signal_11276) ) ;
    buf_clk cell_8746 ( .C (clk), .D (signal_11291), .Q (signal_11292) ) ;
    buf_clk cell_8762 ( .C (clk), .D (signal_11307), .Q (signal_11308) ) ;
    buf_clk cell_8778 ( .C (clk), .D (signal_11323), .Q (signal_11324) ) ;
    buf_clk cell_8794 ( .C (clk), .D (signal_11339), .Q (signal_11340) ) ;
    buf_clk cell_8810 ( .C (clk), .D (signal_11355), .Q (signal_11356) ) ;
    buf_clk cell_8826 ( .C (clk), .D (signal_11371), .Q (signal_11372) ) ;
    buf_clk cell_8842 ( .C (clk), .D (signal_11387), .Q (signal_11388) ) ;
    buf_clk cell_8858 ( .C (clk), .D (signal_11403), .Q (signal_11404) ) ;
    buf_clk cell_8874 ( .C (clk), .D (signal_11419), .Q (signal_11420) ) ;
    buf_clk cell_8890 ( .C (clk), .D (signal_11435), .Q (signal_11436) ) ;
    buf_clk cell_8906 ( .C (clk), .D (signal_11451), .Q (signal_11452) ) ;
    buf_clk cell_8922 ( .C (clk), .D (signal_11467), .Q (signal_11468) ) ;
    buf_clk cell_8938 ( .C (clk), .D (signal_11483), .Q (signal_11484) ) ;
    buf_clk cell_8954 ( .C (clk), .D (signal_11499), .Q (signal_11500) ) ;
    buf_clk cell_8970 ( .C (clk), .D (signal_11515), .Q (signal_11516) ) ;
    buf_clk cell_8986 ( .C (clk), .D (signal_11531), .Q (signal_11532) ) ;
    buf_clk cell_9002 ( .C (clk), .D (signal_11547), .Q (signal_11548) ) ;
    buf_clk cell_9018 ( .C (clk), .D (signal_11563), .Q (signal_11564) ) ;
    buf_clk cell_9034 ( .C (clk), .D (signal_11579), .Q (signal_11580) ) ;
    buf_clk cell_9050 ( .C (clk), .D (signal_11595), .Q (signal_11596) ) ;
    buf_clk cell_9066 ( .C (clk), .D (signal_11611), .Q (signal_11612) ) ;
    buf_clk cell_9082 ( .C (clk), .D (signal_11627), .Q (signal_11628) ) ;
    buf_clk cell_9098 ( .C (clk), .D (signal_11643), .Q (signal_11644) ) ;
    buf_clk cell_9114 ( .C (clk), .D (signal_11659), .Q (signal_11660) ) ;
    buf_clk cell_9130 ( .C (clk), .D (signal_11675), .Q (signal_11676) ) ;
    buf_clk cell_9146 ( .C (clk), .D (signal_11691), .Q (signal_11692) ) ;
    buf_clk cell_9162 ( .C (clk), .D (signal_11707), .Q (signal_11708) ) ;
    buf_clk cell_9178 ( .C (clk), .D (signal_11723), .Q (signal_11724) ) ;
    buf_clk cell_9194 ( .C (clk), .D (signal_11739), .Q (signal_11740) ) ;
    buf_clk cell_9210 ( .C (clk), .D (signal_11755), .Q (signal_11756) ) ;
    buf_clk cell_9226 ( .C (clk), .D (signal_11771), .Q (signal_11772) ) ;
    buf_clk cell_9242 ( .C (clk), .D (signal_11787), .Q (signal_11788) ) ;
    buf_clk cell_9258 ( .C (clk), .D (signal_11803), .Q (signal_11804) ) ;
    buf_clk cell_9274 ( .C (clk), .D (signal_11819), .Q (signal_11820) ) ;
    buf_clk cell_9290 ( .C (clk), .D (signal_11835), .Q (signal_11836) ) ;
    buf_clk cell_9306 ( .C (clk), .D (signal_11851), .Q (signal_11852) ) ;
    buf_clk cell_9322 ( .C (clk), .D (signal_11867), .Q (signal_11868) ) ;
    buf_clk cell_9338 ( .C (clk), .D (signal_11883), .Q (signal_11884) ) ;
    buf_clk cell_9354 ( .C (clk), .D (signal_11899), .Q (signal_11900) ) ;
    buf_clk cell_9370 ( .C (clk), .D (signal_11915), .Q (signal_11916) ) ;
    buf_clk cell_9386 ( .C (clk), .D (signal_11931), .Q (signal_11932) ) ;
    buf_clk cell_9402 ( .C (clk), .D (signal_11947), .Q (signal_11948) ) ;
    buf_clk cell_9418 ( .C (clk), .D (signal_11963), .Q (signal_11964) ) ;
    buf_clk cell_9434 ( .C (clk), .D (signal_11979), .Q (signal_11980) ) ;
    buf_clk cell_9450 ( .C (clk), .D (signal_11995), .Q (signal_11996) ) ;
    buf_clk cell_9466 ( .C (clk), .D (signal_12011), .Q (signal_12012) ) ;
    buf_clk cell_9482 ( .C (clk), .D (signal_12027), .Q (signal_12028) ) ;
    buf_clk cell_9498 ( .C (clk), .D (signal_12043), .Q (signal_12044) ) ;
    buf_clk cell_9514 ( .C (clk), .D (signal_12059), .Q (signal_12060) ) ;
    buf_clk cell_9530 ( .C (clk), .D (signal_12075), .Q (signal_12076) ) ;
    buf_clk cell_9546 ( .C (clk), .D (signal_12091), .Q (signal_12092) ) ;
    buf_clk cell_9562 ( .C (clk), .D (signal_12107), .Q (signal_12108) ) ;
    buf_clk cell_9578 ( .C (clk), .D (signal_12123), .Q (signal_12124) ) ;
    buf_clk cell_9594 ( .C (clk), .D (signal_12139), .Q (signal_12140) ) ;
    buf_clk cell_9610 ( .C (clk), .D (signal_12155), .Q (signal_12156) ) ;
    buf_clk cell_9626 ( .C (clk), .D (signal_12171), .Q (signal_12172) ) ;
    buf_clk cell_9642 ( .C (clk), .D (signal_12187), .Q (signal_12188) ) ;
    buf_clk cell_9658 ( .C (clk), .D (signal_12203), .Q (signal_12204) ) ;
    buf_clk cell_9674 ( .C (clk), .D (signal_12219), .Q (signal_12220) ) ;
    buf_clk cell_9690 ( .C (clk), .D (signal_12235), .Q (signal_12236) ) ;
    buf_clk cell_9706 ( .C (clk), .D (signal_12251), .Q (signal_12252) ) ;
    buf_clk cell_9722 ( .C (clk), .D (signal_12267), .Q (signal_12268) ) ;
    buf_clk cell_9738 ( .C (clk), .D (signal_12283), .Q (signal_12284) ) ;
    buf_clk cell_9754 ( .C (clk), .D (signal_12299), .Q (signal_12300) ) ;
    buf_clk cell_9770 ( .C (clk), .D (signal_12315), .Q (signal_12316) ) ;
    buf_clk cell_9786 ( .C (clk), .D (signal_12331), .Q (signal_12332) ) ;
    buf_clk cell_9802 ( .C (clk), .D (signal_12347), .Q (signal_12348) ) ;
    buf_clk cell_9818 ( .C (clk), .D (signal_12363), .Q (signal_12364) ) ;
    buf_clk cell_9834 ( .C (clk), .D (signal_12379), .Q (signal_12380) ) ;
    buf_clk cell_9850 ( .C (clk), .D (signal_12395), .Q (signal_12396) ) ;
    buf_clk cell_9866 ( .C (clk), .D (signal_12411), .Q (signal_12412) ) ;
    buf_clk cell_9882 ( .C (clk), .D (signal_12427), .Q (signal_12428) ) ;
    buf_clk cell_9898 ( .C (clk), .D (signal_12443), .Q (signal_12444) ) ;
    buf_clk cell_9914 ( .C (clk), .D (signal_12459), .Q (signal_12460) ) ;
    buf_clk cell_9930 ( .C (clk), .D (signal_12475), .Q (signal_12476) ) ;
    buf_clk cell_9946 ( .C (clk), .D (signal_12491), .Q (signal_12492) ) ;
    buf_clk cell_9962 ( .C (clk), .D (signal_12507), .Q (signal_12508) ) ;
    buf_clk cell_9978 ( .C (clk), .D (signal_12523), .Q (signal_12524) ) ;
    buf_clk cell_9994 ( .C (clk), .D (signal_12539), .Q (signal_12540) ) ;
    buf_clk cell_10010 ( .C (clk), .D (signal_12555), .Q (signal_12556) ) ;
    buf_clk cell_10026 ( .C (clk), .D (signal_12571), .Q (signal_12572) ) ;
    buf_clk cell_10042 ( .C (clk), .D (signal_12587), .Q (signal_12588) ) ;
    buf_clk cell_10058 ( .C (clk), .D (signal_12603), .Q (signal_12604) ) ;
    buf_clk cell_10074 ( .C (clk), .D (signal_12619), .Q (signal_12620) ) ;
    buf_clk cell_10090 ( .C (clk), .D (signal_12635), .Q (signal_12636) ) ;
    buf_clk cell_10106 ( .C (clk), .D (signal_12651), .Q (signal_12652) ) ;
    buf_clk cell_10122 ( .C (clk), .D (signal_12667), .Q (signal_12668) ) ;
    buf_clk cell_10138 ( .C (clk), .D (signal_12683), .Q (signal_12684) ) ;
    buf_clk cell_10154 ( .C (clk), .D (signal_12699), .Q (signal_12700) ) ;
    buf_clk cell_10170 ( .C (clk), .D (signal_12715), .Q (signal_12716) ) ;
    buf_clk cell_10186 ( .C (clk), .D (signal_12731), .Q (signal_12732) ) ;
    buf_clk cell_10202 ( .C (clk), .D (signal_12747), .Q (signal_12748) ) ;
    buf_clk cell_10218 ( .C (clk), .D (signal_12763), .Q (signal_12764) ) ;
    buf_clk cell_10234 ( .C (clk), .D (signal_12779), .Q (signal_12780) ) ;
    buf_clk cell_10250 ( .C (clk), .D (signal_12795), .Q (signal_12796) ) ;
    buf_clk cell_10266 ( .C (clk), .D (signal_12811), .Q (signal_12812) ) ;
    buf_clk cell_10282 ( .C (clk), .D (signal_12827), .Q (signal_12828) ) ;
    buf_clk cell_10298 ( .C (clk), .D (signal_12843), .Q (signal_12844) ) ;
    buf_clk cell_10314 ( .C (clk), .D (signal_12859), .Q (signal_12860) ) ;
    buf_clk cell_10330 ( .C (clk), .D (signal_12875), .Q (signal_12876) ) ;
    buf_clk cell_10346 ( .C (clk), .D (signal_12891), .Q (signal_12892) ) ;
    buf_clk cell_10362 ( .C (clk), .D (signal_12907), .Q (signal_12908) ) ;
    buf_clk cell_10378 ( .C (clk), .D (signal_12923), .Q (signal_12924) ) ;
    buf_clk cell_10394 ( .C (clk), .D (signal_12939), .Q (signal_12940) ) ;
    buf_clk cell_10410 ( .C (clk), .D (signal_12955), .Q (signal_12956) ) ;
    buf_clk cell_10426 ( .C (clk), .D (signal_12971), .Q (signal_12972) ) ;
    buf_clk cell_10442 ( .C (clk), .D (signal_12987), .Q (signal_12988) ) ;
    buf_clk cell_10458 ( .C (clk), .D (signal_13003), .Q (signal_13004) ) ;
    buf_clk cell_10474 ( .C (clk), .D (signal_13019), .Q (signal_13020) ) ;
    buf_clk cell_10490 ( .C (clk), .D (signal_13035), .Q (signal_13036) ) ;
    buf_clk cell_10506 ( .C (clk), .D (signal_13051), .Q (signal_13052) ) ;
    buf_clk cell_10522 ( .C (clk), .D (signal_13067), .Q (signal_13068) ) ;
    buf_clk cell_10538 ( .C (clk), .D (signal_13083), .Q (signal_13084) ) ;
    buf_clk cell_10554 ( .C (clk), .D (signal_13099), .Q (signal_13100) ) ;
    buf_clk cell_10570 ( .C (clk), .D (signal_13115), .Q (signal_13116) ) ;
    buf_clk cell_10586 ( .C (clk), .D (signal_13131), .Q (signal_13132) ) ;
    buf_clk cell_10602 ( .C (clk), .D (signal_13147), .Q (signal_13148) ) ;
    buf_clk cell_10618 ( .C (clk), .D (signal_13163), .Q (signal_13164) ) ;
    buf_clk cell_10634 ( .C (clk), .D (signal_13179), .Q (signal_13180) ) ;
    buf_clk cell_10650 ( .C (clk), .D (signal_13195), .Q (signal_13196) ) ;
    buf_clk cell_10666 ( .C (clk), .D (signal_13211), .Q (signal_13212) ) ;
    buf_clk cell_10682 ( .C (clk), .D (signal_13227), .Q (signal_13228) ) ;
    buf_clk cell_10698 ( .C (clk), .D (signal_13243), .Q (signal_13244) ) ;
    buf_clk cell_10714 ( .C (clk), .D (signal_13259), .Q (signal_13260) ) ;
    buf_clk cell_10730 ( .C (clk), .D (signal_13275), .Q (signal_13276) ) ;
    buf_clk cell_10746 ( .C (clk), .D (signal_13291), .Q (signal_13292) ) ;
    buf_clk cell_10762 ( .C (clk), .D (signal_13307), .Q (signal_13308) ) ;
    buf_clk cell_10778 ( .C (clk), .D (signal_13323), .Q (signal_13324) ) ;
    buf_clk cell_10794 ( .C (clk), .D (signal_13339), .Q (signal_13340) ) ;
    buf_clk cell_10810 ( .C (clk), .D (signal_13355), .Q (signal_13356) ) ;
    buf_clk cell_10826 ( .C (clk), .D (signal_13371), .Q (signal_13372) ) ;
    buf_clk cell_10842 ( .C (clk), .D (signal_13387), .Q (signal_13388) ) ;
    buf_clk cell_10858 ( .C (clk), .D (signal_13403), .Q (signal_13404) ) ;
    buf_clk cell_10874 ( .C (clk), .D (signal_13419), .Q (signal_13420) ) ;
    buf_clk cell_10890 ( .C (clk), .D (signal_13435), .Q (signal_13436) ) ;
    buf_clk cell_10906 ( .C (clk), .D (signal_13451), .Q (signal_13452) ) ;
    buf_clk cell_10922 ( .C (clk), .D (signal_13467), .Q (signal_13468) ) ;
    buf_clk cell_10938 ( .C (clk), .D (signal_13483), .Q (signal_13484) ) ;
    buf_clk cell_10954 ( .C (clk), .D (signal_13499), .Q (signal_13500) ) ;
    buf_clk cell_10970 ( .C (clk), .D (signal_13515), .Q (signal_13516) ) ;
    buf_clk cell_10986 ( .C (clk), .D (signal_13531), .Q (signal_13532) ) ;
    buf_clk cell_11002 ( .C (clk), .D (signal_13547), .Q (signal_13548) ) ;
    buf_clk cell_11018 ( .C (clk), .D (signal_13563), .Q (signal_13564) ) ;
    buf_clk cell_11034 ( .C (clk), .D (signal_13579), .Q (signal_13580) ) ;
    buf_clk cell_11050 ( .C (clk), .D (signal_13595), .Q (signal_13596) ) ;
    buf_clk cell_11066 ( .C (clk), .D (signal_13611), .Q (signal_13612) ) ;
    buf_clk cell_11082 ( .C (clk), .D (signal_13627), .Q (signal_13628) ) ;
    buf_clk cell_11098 ( .C (clk), .D (signal_13643), .Q (signal_13644) ) ;
    buf_clk cell_11114 ( .C (clk), .D (signal_13659), .Q (signal_13660) ) ;
    buf_clk cell_11130 ( .C (clk), .D (signal_13675), .Q (signal_13676) ) ;
    buf_clk cell_11146 ( .C (clk), .D (signal_13691), .Q (signal_13692) ) ;
    buf_clk cell_11162 ( .C (clk), .D (signal_13707), .Q (signal_13708) ) ;
    buf_clk cell_11178 ( .C (clk), .D (signal_13723), .Q (signal_13724) ) ;
    buf_clk cell_11194 ( .C (clk), .D (signal_13739), .Q (signal_13740) ) ;
    buf_clk cell_11210 ( .C (clk), .D (signal_13755), .Q (signal_13756) ) ;
    buf_clk cell_11226 ( .C (clk), .D (signal_13771), .Q (signal_13772) ) ;
    buf_clk cell_11242 ( .C (clk), .D (signal_13787), .Q (signal_13788) ) ;
    buf_clk cell_11258 ( .C (clk), .D (signal_13803), .Q (signal_13804) ) ;
    buf_clk cell_11274 ( .C (clk), .D (signal_13819), .Q (signal_13820) ) ;
    buf_clk cell_11290 ( .C (clk), .D (signal_13835), .Q (signal_13836) ) ;
    buf_clk cell_11306 ( .C (clk), .D (signal_13851), .Q (signal_13852) ) ;
    buf_clk cell_11322 ( .C (clk), .D (signal_13867), .Q (signal_13868) ) ;
    buf_clk cell_11338 ( .C (clk), .D (signal_13883), .Q (signal_13884) ) ;
    buf_clk cell_11354 ( .C (clk), .D (signal_13899), .Q (signal_13900) ) ;
    buf_clk cell_11370 ( .C (clk), .D (signal_13915), .Q (signal_13916) ) ;
    buf_clk cell_11386 ( .C (clk), .D (signal_13931), .Q (signal_13932) ) ;
    buf_clk cell_11402 ( .C (clk), .D (signal_13947), .Q (signal_13948) ) ;
    buf_clk cell_11418 ( .C (clk), .D (signal_13963), .Q (signal_13964) ) ;
    buf_clk cell_11434 ( .C (clk), .D (signal_13979), .Q (signal_13980) ) ;
    buf_clk cell_11450 ( .C (clk), .D (signal_13995), .Q (signal_13996) ) ;
    buf_clk cell_11466 ( .C (clk), .D (signal_14011), .Q (signal_14012) ) ;
    buf_clk cell_11482 ( .C (clk), .D (signal_14027), .Q (signal_14028) ) ;
    buf_clk cell_11498 ( .C (clk), .D (signal_14043), .Q (signal_14044) ) ;
    buf_clk cell_11514 ( .C (clk), .D (signal_14059), .Q (signal_14060) ) ;
    buf_clk cell_11530 ( .C (clk), .D (signal_14075), .Q (signal_14076) ) ;
    buf_clk cell_11546 ( .C (clk), .D (signal_14091), .Q (signal_14092) ) ;
    buf_clk cell_11562 ( .C (clk), .D (signal_14107), .Q (signal_14108) ) ;
    buf_clk cell_11578 ( .C (clk), .D (signal_14123), .Q (signal_14124) ) ;
    buf_clk cell_11594 ( .C (clk), .D (signal_14139), .Q (signal_14140) ) ;
    buf_clk cell_11610 ( .C (clk), .D (signal_14155), .Q (signal_14156) ) ;
    buf_clk cell_11626 ( .C (clk), .D (signal_14171), .Q (signal_14172) ) ;
    buf_clk cell_11642 ( .C (clk), .D (signal_14187), .Q (signal_14188) ) ;
    buf_clk cell_11658 ( .C (clk), .D (signal_14203), .Q (signal_14204) ) ;
    buf_clk cell_11674 ( .C (clk), .D (signal_14219), .Q (signal_14220) ) ;
    buf_clk cell_11690 ( .C (clk), .D (signal_14235), .Q (signal_14236) ) ;
    buf_clk cell_11706 ( .C (clk), .D (signal_14251), .Q (signal_14252) ) ;
    buf_clk cell_11722 ( .C (clk), .D (signal_14267), .Q (signal_14268) ) ;
    buf_clk cell_11738 ( .C (clk), .D (signal_14283), .Q (signal_14284) ) ;
    buf_clk cell_11754 ( .C (clk), .D (signal_14299), .Q (signal_14300) ) ;
    buf_clk cell_11770 ( .C (clk), .D (signal_14315), .Q (signal_14316) ) ;
    buf_clk cell_11786 ( .C (clk), .D (signal_14331), .Q (signal_14332) ) ;
    buf_clk cell_11802 ( .C (clk), .D (signal_14347), .Q (signal_14348) ) ;
    buf_clk cell_11818 ( .C (clk), .D (signal_14363), .Q (signal_14364) ) ;
    buf_clk cell_11834 ( .C (clk), .D (signal_14379), .Q (signal_14380) ) ;
    buf_clk cell_11850 ( .C (clk), .D (signal_14395), .Q (signal_14396) ) ;
    buf_clk cell_11866 ( .C (clk), .D (signal_14411), .Q (signal_14412) ) ;
    buf_clk cell_11882 ( .C (clk), .D (signal_14427), .Q (signal_14428) ) ;
    buf_clk cell_11898 ( .C (clk), .D (signal_14443), .Q (signal_14444) ) ;
    buf_clk cell_11914 ( .C (clk), .D (signal_14459), .Q (signal_14460) ) ;
    buf_clk cell_11930 ( .C (clk), .D (signal_14475), .Q (signal_14476) ) ;
    buf_clk cell_11946 ( .C (clk), .D (signal_14491), .Q (signal_14492) ) ;
    buf_clk cell_11962 ( .C (clk), .D (signal_14507), .Q (signal_14508) ) ;
    buf_clk cell_11978 ( .C (clk), .D (signal_14523), .Q (signal_14524) ) ;
    buf_clk cell_11994 ( .C (clk), .D (signal_14539), .Q (signal_14540) ) ;
    buf_clk cell_12010 ( .C (clk), .D (signal_14555), .Q (signal_14556) ) ;
    buf_clk cell_12026 ( .C (clk), .D (signal_14571), .Q (signal_14572) ) ;
    buf_clk cell_12042 ( .C (clk), .D (signal_14587), .Q (signal_14588) ) ;
    buf_clk cell_12058 ( .C (clk), .D (signal_14603), .Q (signal_14604) ) ;
    buf_clk cell_12074 ( .C (clk), .D (signal_14619), .Q (signal_14620) ) ;
    buf_clk cell_12090 ( .C (clk), .D (signal_14635), .Q (signal_14636) ) ;
    buf_clk cell_12106 ( .C (clk), .D (signal_14651), .Q (signal_14652) ) ;
    buf_clk cell_12122 ( .C (clk), .D (signal_14667), .Q (signal_14668) ) ;
    buf_clk cell_12138 ( .C (clk), .D (signal_14683), .Q (signal_14684) ) ;
    buf_clk cell_12154 ( .C (clk), .D (signal_14699), .Q (signal_14700) ) ;
    buf_clk cell_12170 ( .C (clk), .D (signal_14715), .Q (signal_14716) ) ;
    buf_clk cell_12186 ( .C (clk), .D (signal_14731), .Q (signal_14732) ) ;
    buf_clk cell_12202 ( .C (clk), .D (signal_14747), .Q (signal_14748) ) ;
    buf_clk cell_12218 ( .C (clk), .D (signal_14763), .Q (signal_14764) ) ;
    buf_clk cell_12234 ( .C (clk), .D (signal_14779), .Q (signal_14780) ) ;
    buf_clk cell_12250 ( .C (clk), .D (signal_14795), .Q (signal_14796) ) ;
    buf_clk cell_12266 ( .C (clk), .D (signal_14811), .Q (signal_14812) ) ;
    buf_clk cell_12282 ( .C (clk), .D (signal_14827), .Q (signal_14828) ) ;
    buf_clk cell_12298 ( .C (clk), .D (signal_14843), .Q (signal_14844) ) ;
    buf_clk cell_12314 ( .C (clk), .D (signal_14859), .Q (signal_14860) ) ;
    buf_clk cell_12330 ( .C (clk), .D (signal_14875), .Q (signal_14876) ) ;
    buf_clk cell_12346 ( .C (clk), .D (signal_14891), .Q (signal_14892) ) ;
    buf_clk cell_12362 ( .C (clk), .D (signal_14907), .Q (signal_14908) ) ;
    buf_clk cell_12378 ( .C (clk), .D (signal_14923), .Q (signal_14924) ) ;
    buf_clk cell_12394 ( .C (clk), .D (signal_14939), .Q (signal_14940) ) ;

    /* cells in depth 15 */
    buf_clk cell_2399 ( .C (clk), .D (signal_4944), .Q (signal_4945) ) ;
    buf_clk cell_2415 ( .C (clk), .D (signal_4960), .Q (signal_4961) ) ;
    buf_clk cell_2431 ( .C (clk), .D (signal_4976), .Q (signal_4977) ) ;
    buf_clk cell_2447 ( .C (clk), .D (signal_4992), .Q (signal_4993) ) ;
    buf_clk cell_2463 ( .C (clk), .D (signal_5008), .Q (signal_5009) ) ;
    buf_clk cell_2479 ( .C (clk), .D (signal_5024), .Q (signal_5025) ) ;
    buf_clk cell_2495 ( .C (clk), .D (signal_5040), .Q (signal_5041) ) ;
    buf_clk cell_2511 ( .C (clk), .D (signal_5056), .Q (signal_5057) ) ;
    buf_clk cell_2527 ( .C (clk), .D (signal_5072), .Q (signal_5073) ) ;
    buf_clk cell_2543 ( .C (clk), .D (signal_5088), .Q (signal_5089) ) ;
    buf_clk cell_2559 ( .C (clk), .D (signal_5104), .Q (signal_5105) ) ;
    buf_clk cell_2575 ( .C (clk), .D (signal_5120), .Q (signal_5121) ) ;
    buf_clk cell_2591 ( .C (clk), .D (signal_5136), .Q (signal_5137) ) ;
    buf_clk cell_2607 ( .C (clk), .D (signal_5152), .Q (signal_5153) ) ;
    buf_clk cell_2623 ( .C (clk), .D (signal_5168), .Q (signal_5169) ) ;
    buf_clk cell_2639 ( .C (clk), .D (signal_5184), .Q (signal_5185) ) ;
    buf_clk cell_2655 ( .C (clk), .D (signal_5200), .Q (signal_5201) ) ;
    buf_clk cell_2671 ( .C (clk), .D (signal_5216), .Q (signal_5217) ) ;
    buf_clk cell_2687 ( .C (clk), .D (signal_5232), .Q (signal_5233) ) ;
    buf_clk cell_2703 ( .C (clk), .D (signal_5248), .Q (signal_5249) ) ;
    buf_clk cell_2719 ( .C (clk), .D (signal_5264), .Q (signal_5265) ) ;
    buf_clk cell_2735 ( .C (clk), .D (signal_5280), .Q (signal_5281) ) ;
    buf_clk cell_2751 ( .C (clk), .D (signal_5296), .Q (signal_5297) ) ;
    buf_clk cell_2767 ( .C (clk), .D (signal_5312), .Q (signal_5313) ) ;
    buf_clk cell_2783 ( .C (clk), .D (signal_5328), .Q (signal_5329) ) ;
    buf_clk cell_2799 ( .C (clk), .D (signal_5344), .Q (signal_5345) ) ;
    buf_clk cell_2815 ( .C (clk), .D (signal_5360), .Q (signal_5361) ) ;
    buf_clk cell_2831 ( .C (clk), .D (signal_5376), .Q (signal_5377) ) ;
    buf_clk cell_2847 ( .C (clk), .D (signal_5392), .Q (signal_5393) ) ;
    buf_clk cell_2863 ( .C (clk), .D (signal_5408), .Q (signal_5409) ) ;
    buf_clk cell_2879 ( .C (clk), .D (signal_5424), .Q (signal_5425) ) ;
    buf_clk cell_2895 ( .C (clk), .D (signal_5440), .Q (signal_5441) ) ;
    buf_clk cell_2911 ( .C (clk), .D (signal_5456), .Q (signal_5457) ) ;
    buf_clk cell_2927 ( .C (clk), .D (signal_5472), .Q (signal_5473) ) ;
    buf_clk cell_2943 ( .C (clk), .D (signal_5488), .Q (signal_5489) ) ;
    buf_clk cell_2959 ( .C (clk), .D (signal_5504), .Q (signal_5505) ) ;
    buf_clk cell_2975 ( .C (clk), .D (signal_5520), .Q (signal_5521) ) ;
    buf_clk cell_2991 ( .C (clk), .D (signal_5536), .Q (signal_5537) ) ;
    buf_clk cell_3007 ( .C (clk), .D (signal_5552), .Q (signal_5553) ) ;
    buf_clk cell_3023 ( .C (clk), .D (signal_5568), .Q (signal_5569) ) ;
    buf_clk cell_3039 ( .C (clk), .D (signal_5584), .Q (signal_5585) ) ;
    buf_clk cell_3055 ( .C (clk), .D (signal_5600), .Q (signal_5601) ) ;
    buf_clk cell_3071 ( .C (clk), .D (signal_5616), .Q (signal_5617) ) ;
    buf_clk cell_3087 ( .C (clk), .D (signal_5632), .Q (signal_5633) ) ;
    buf_clk cell_3103 ( .C (clk), .D (signal_5648), .Q (signal_5649) ) ;
    buf_clk cell_3119 ( .C (clk), .D (signal_5664), .Q (signal_5665) ) ;
    buf_clk cell_3135 ( .C (clk), .D (signal_5680), .Q (signal_5681) ) ;
    buf_clk cell_3151 ( .C (clk), .D (signal_5696), .Q (signal_5697) ) ;
    buf_clk cell_3167 ( .C (clk), .D (signal_5712), .Q (signal_5713) ) ;
    buf_clk cell_3183 ( .C (clk), .D (signal_5728), .Q (signal_5729) ) ;
    buf_clk cell_3199 ( .C (clk), .D (signal_5744), .Q (signal_5745) ) ;
    buf_clk cell_3215 ( .C (clk), .D (signal_5760), .Q (signal_5761) ) ;
    buf_clk cell_3231 ( .C (clk), .D (signal_5776), .Q (signal_5777) ) ;
    buf_clk cell_3247 ( .C (clk), .D (signal_5792), .Q (signal_5793) ) ;
    buf_clk cell_3263 ( .C (clk), .D (signal_5808), .Q (signal_5809) ) ;
    buf_clk cell_3279 ( .C (clk), .D (signal_5824), .Q (signal_5825) ) ;
    buf_clk cell_3295 ( .C (clk), .D (signal_5840), .Q (signal_5841) ) ;
    buf_clk cell_3311 ( .C (clk), .D (signal_5856), .Q (signal_5857) ) ;
    buf_clk cell_3327 ( .C (clk), .D (signal_5872), .Q (signal_5873) ) ;
    buf_clk cell_3343 ( .C (clk), .D (signal_5888), .Q (signal_5889) ) ;
    buf_clk cell_3359 ( .C (clk), .D (signal_5904), .Q (signal_5905) ) ;
    buf_clk cell_3375 ( .C (clk), .D (signal_5920), .Q (signal_5921) ) ;
    buf_clk cell_3391 ( .C (clk), .D (signal_5936), .Q (signal_5937) ) ;
    buf_clk cell_3407 ( .C (clk), .D (signal_5952), .Q (signal_5953) ) ;
    buf_clk cell_3423 ( .C (clk), .D (signal_5968), .Q (signal_5969) ) ;
    buf_clk cell_3439 ( .C (clk), .D (signal_5984), .Q (signal_5985) ) ;
    buf_clk cell_3455 ( .C (clk), .D (signal_6000), .Q (signal_6001) ) ;
    buf_clk cell_3471 ( .C (clk), .D (signal_6016), .Q (signal_6017) ) ;
    buf_clk cell_3487 ( .C (clk), .D (signal_6032), .Q (signal_6033) ) ;
    buf_clk cell_3503 ( .C (clk), .D (signal_6048), .Q (signal_6049) ) ;
    buf_clk cell_3519 ( .C (clk), .D (signal_6064), .Q (signal_6065) ) ;
    buf_clk cell_3535 ( .C (clk), .D (signal_6080), .Q (signal_6081) ) ;
    buf_clk cell_3551 ( .C (clk), .D (signal_6096), .Q (signal_6097) ) ;
    buf_clk cell_3567 ( .C (clk), .D (signal_6112), .Q (signal_6113) ) ;
    buf_clk cell_3583 ( .C (clk), .D (signal_6128), .Q (signal_6129) ) ;
    buf_clk cell_3599 ( .C (clk), .D (signal_6144), .Q (signal_6145) ) ;
    buf_clk cell_3615 ( .C (clk), .D (signal_6160), .Q (signal_6161) ) ;
    buf_clk cell_3631 ( .C (clk), .D (signal_6176), .Q (signal_6177) ) ;
    buf_clk cell_3647 ( .C (clk), .D (signal_6192), .Q (signal_6193) ) ;
    buf_clk cell_3663 ( .C (clk), .D (signal_6208), .Q (signal_6209) ) ;
    buf_clk cell_3679 ( .C (clk), .D (signal_6224), .Q (signal_6225) ) ;
    buf_clk cell_3695 ( .C (clk), .D (signal_6240), .Q (signal_6241) ) ;
    buf_clk cell_3711 ( .C (clk), .D (signal_6256), .Q (signal_6257) ) ;
    buf_clk cell_3727 ( .C (clk), .D (signal_6272), .Q (signal_6273) ) ;
    buf_clk cell_3743 ( .C (clk), .D (signal_6288), .Q (signal_6289) ) ;
    buf_clk cell_3759 ( .C (clk), .D (signal_6304), .Q (signal_6305) ) ;
    buf_clk cell_3775 ( .C (clk), .D (signal_6320), .Q (signal_6321) ) ;
    buf_clk cell_3791 ( .C (clk), .D (signal_6336), .Q (signal_6337) ) ;
    buf_clk cell_3807 ( .C (clk), .D (signal_6352), .Q (signal_6353) ) ;
    buf_clk cell_3823 ( .C (clk), .D (signal_6368), .Q (signal_6369) ) ;
    buf_clk cell_3839 ( .C (clk), .D (signal_6384), .Q (signal_6385) ) ;
    buf_clk cell_3855 ( .C (clk), .D (signal_6400), .Q (signal_6401) ) ;
    buf_clk cell_3871 ( .C (clk), .D (signal_6416), .Q (signal_6417) ) ;
    buf_clk cell_3887 ( .C (clk), .D (signal_6432), .Q (signal_6433) ) ;
    buf_clk cell_3903 ( .C (clk), .D (signal_6448), .Q (signal_6449) ) ;
    buf_clk cell_3919 ( .C (clk), .D (signal_6464), .Q (signal_6465) ) ;
    buf_clk cell_3935 ( .C (clk), .D (signal_6480), .Q (signal_6481) ) ;
    buf_clk cell_3951 ( .C (clk), .D (signal_6496), .Q (signal_6497) ) ;
    buf_clk cell_3967 ( .C (clk), .D (signal_6512), .Q (signal_6513) ) ;
    buf_clk cell_3983 ( .C (clk), .D (signal_6528), .Q (signal_6529) ) ;
    buf_clk cell_3999 ( .C (clk), .D (signal_6544), .Q (signal_6545) ) ;
    buf_clk cell_4015 ( .C (clk), .D (signal_6560), .Q (signal_6561) ) ;
    buf_clk cell_4031 ( .C (clk), .D (signal_6576), .Q (signal_6577) ) ;
    buf_clk cell_4047 ( .C (clk), .D (signal_6592), .Q (signal_6593) ) ;
    buf_clk cell_4063 ( .C (clk), .D (signal_6608), .Q (signal_6609) ) ;
    buf_clk cell_4079 ( .C (clk), .D (signal_6624), .Q (signal_6625) ) ;
    buf_clk cell_4095 ( .C (clk), .D (signal_6640), .Q (signal_6641) ) ;
    buf_clk cell_4111 ( .C (clk), .D (signal_6656), .Q (signal_6657) ) ;
    buf_clk cell_4127 ( .C (clk), .D (signal_6672), .Q (signal_6673) ) ;
    buf_clk cell_4143 ( .C (clk), .D (signal_6688), .Q (signal_6689) ) ;
    buf_clk cell_4159 ( .C (clk), .D (signal_6704), .Q (signal_6705) ) ;
    buf_clk cell_4175 ( .C (clk), .D (signal_6720), .Q (signal_6721) ) ;
    buf_clk cell_4191 ( .C (clk), .D (signal_6736), .Q (signal_6737) ) ;
    buf_clk cell_4207 ( .C (clk), .D (signal_6752), .Q (signal_6753) ) ;
    buf_clk cell_4223 ( .C (clk), .D (signal_6768), .Q (signal_6769) ) ;
    buf_clk cell_4239 ( .C (clk), .D (signal_6784), .Q (signal_6785) ) ;
    buf_clk cell_4255 ( .C (clk), .D (signal_6800), .Q (signal_6801) ) ;
    buf_clk cell_4271 ( .C (clk), .D (signal_6816), .Q (signal_6817) ) ;
    buf_clk cell_4287 ( .C (clk), .D (signal_6832), .Q (signal_6833) ) ;
    buf_clk cell_4303 ( .C (clk), .D (signal_6848), .Q (signal_6849) ) ;
    buf_clk cell_4319 ( .C (clk), .D (signal_6864), .Q (signal_6865) ) ;
    buf_clk cell_4335 ( .C (clk), .D (signal_6880), .Q (signal_6881) ) ;
    buf_clk cell_4351 ( .C (clk), .D (signal_6896), .Q (signal_6897) ) ;
    buf_clk cell_4367 ( .C (clk), .D (signal_6912), .Q (signal_6913) ) ;
    buf_clk cell_4383 ( .C (clk), .D (signal_6928), .Q (signal_6929) ) ;
    buf_clk cell_4399 ( .C (clk), .D (signal_6944), .Q (signal_6945) ) ;
    buf_clk cell_4443 ( .C (clk), .D (signal_6988), .Q (signal_6989) ) ;
    buf_clk cell_4459 ( .C (clk), .D (signal_7004), .Q (signal_7005) ) ;
    buf_clk cell_4475 ( .C (clk), .D (signal_7020), .Q (signal_7021) ) ;
    buf_clk cell_4491 ( .C (clk), .D (signal_7036), .Q (signal_7037) ) ;
    buf_clk cell_4507 ( .C (clk), .D (signal_7052), .Q (signal_7053) ) ;
    buf_clk cell_4523 ( .C (clk), .D (signal_7068), .Q (signal_7069) ) ;
    buf_clk cell_4539 ( .C (clk), .D (signal_7084), .Q (signal_7085) ) ;
    buf_clk cell_4555 ( .C (clk), .D (signal_7100), .Q (signal_7101) ) ;
    buf_clk cell_4571 ( .C (clk), .D (signal_7116), .Q (signal_7117) ) ;
    buf_clk cell_4587 ( .C (clk), .D (signal_7132), .Q (signal_7133) ) ;
    buf_clk cell_4603 ( .C (clk), .D (signal_7148), .Q (signal_7149) ) ;
    buf_clk cell_4619 ( .C (clk), .D (signal_7164), .Q (signal_7165) ) ;
    buf_clk cell_4635 ( .C (clk), .D (signal_7180), .Q (signal_7181) ) ;
    buf_clk cell_4651 ( .C (clk), .D (signal_7196), .Q (signal_7197) ) ;
    buf_clk cell_4667 ( .C (clk), .D (signal_7212), .Q (signal_7213) ) ;
    buf_clk cell_4683 ( .C (clk), .D (signal_7228), .Q (signal_7229) ) ;
    buf_clk cell_4699 ( .C (clk), .D (signal_7244), .Q (signal_7245) ) ;
    buf_clk cell_4715 ( .C (clk), .D (signal_7260), .Q (signal_7261) ) ;
    buf_clk cell_4731 ( .C (clk), .D (signal_7276), .Q (signal_7277) ) ;
    buf_clk cell_4747 ( .C (clk), .D (signal_7292), .Q (signal_7293) ) ;
    buf_clk cell_4763 ( .C (clk), .D (signal_7308), .Q (signal_7309) ) ;
    buf_clk cell_4779 ( .C (clk), .D (signal_7324), .Q (signal_7325) ) ;
    buf_clk cell_4795 ( .C (clk), .D (signal_7340), .Q (signal_7341) ) ;
    buf_clk cell_4811 ( .C (clk), .D (signal_7356), .Q (signal_7357) ) ;
    buf_clk cell_4827 ( .C (clk), .D (signal_7372), .Q (signal_7373) ) ;
    buf_clk cell_4843 ( .C (clk), .D (signal_7388), .Q (signal_7389) ) ;
    buf_clk cell_4859 ( .C (clk), .D (signal_7404), .Q (signal_7405) ) ;
    buf_clk cell_4875 ( .C (clk), .D (signal_7420), .Q (signal_7421) ) ;
    buf_clk cell_4891 ( .C (clk), .D (signal_7436), .Q (signal_7437) ) ;
    buf_clk cell_4907 ( .C (clk), .D (signal_7452), .Q (signal_7453) ) ;
    buf_clk cell_4923 ( .C (clk), .D (signal_7468), .Q (signal_7469) ) ;
    buf_clk cell_4939 ( .C (clk), .D (signal_7484), .Q (signal_7485) ) ;
    buf_clk cell_4955 ( .C (clk), .D (signal_7500), .Q (signal_7501) ) ;
    buf_clk cell_4971 ( .C (clk), .D (signal_7516), .Q (signal_7517) ) ;
    buf_clk cell_4987 ( .C (clk), .D (signal_7532), .Q (signal_7533) ) ;
    buf_clk cell_5003 ( .C (clk), .D (signal_7548), .Q (signal_7549) ) ;
    buf_clk cell_5019 ( .C (clk), .D (signal_7564), .Q (signal_7565) ) ;
    buf_clk cell_5035 ( .C (clk), .D (signal_7580), .Q (signal_7581) ) ;
    buf_clk cell_5051 ( .C (clk), .D (signal_7596), .Q (signal_7597) ) ;
    buf_clk cell_5067 ( .C (clk), .D (signal_7612), .Q (signal_7613) ) ;
    buf_clk cell_5083 ( .C (clk), .D (signal_7628), .Q (signal_7629) ) ;
    buf_clk cell_5099 ( .C (clk), .D (signal_7644), .Q (signal_7645) ) ;
    buf_clk cell_5115 ( .C (clk), .D (signal_7660), .Q (signal_7661) ) ;
    buf_clk cell_5131 ( .C (clk), .D (signal_7676), .Q (signal_7677) ) ;
    buf_clk cell_5147 ( .C (clk), .D (signal_7692), .Q (signal_7693) ) ;
    buf_clk cell_5163 ( .C (clk), .D (signal_7708), .Q (signal_7709) ) ;
    buf_clk cell_5179 ( .C (clk), .D (signal_7724), .Q (signal_7725) ) ;
    buf_clk cell_5195 ( .C (clk), .D (signal_7740), .Q (signal_7741) ) ;
    buf_clk cell_5211 ( .C (clk), .D (signal_7756), .Q (signal_7757) ) ;
    buf_clk cell_5227 ( .C (clk), .D (signal_7772), .Q (signal_7773) ) ;
    buf_clk cell_5243 ( .C (clk), .D (signal_7788), .Q (signal_7789) ) ;
    buf_clk cell_5259 ( .C (clk), .D (signal_7804), .Q (signal_7805) ) ;
    buf_clk cell_5275 ( .C (clk), .D (signal_7820), .Q (signal_7821) ) ;
    buf_clk cell_5291 ( .C (clk), .D (signal_7836), .Q (signal_7837) ) ;
    buf_clk cell_5307 ( .C (clk), .D (signal_7852), .Q (signal_7853) ) ;
    buf_clk cell_5323 ( .C (clk), .D (signal_7868), .Q (signal_7869) ) ;
    buf_clk cell_5339 ( .C (clk), .D (signal_7884), .Q (signal_7885) ) ;
    buf_clk cell_5355 ( .C (clk), .D (signal_7900), .Q (signal_7901) ) ;
    buf_clk cell_5371 ( .C (clk), .D (signal_7916), .Q (signal_7917) ) ;
    buf_clk cell_5387 ( .C (clk), .D (signal_7932), .Q (signal_7933) ) ;
    buf_clk cell_5403 ( .C (clk), .D (signal_7948), .Q (signal_7949) ) ;
    buf_clk cell_5419 ( .C (clk), .D (signal_7964), .Q (signal_7965) ) ;
    buf_clk cell_5435 ( .C (clk), .D (signal_7980), .Q (signal_7981) ) ;
    buf_clk cell_5451 ( .C (clk), .D (signal_7996), .Q (signal_7997) ) ;
    buf_clk cell_5467 ( .C (clk), .D (signal_8012), .Q (signal_8013) ) ;
    buf_clk cell_5483 ( .C (clk), .D (signal_8028), .Q (signal_8029) ) ;
    buf_clk cell_5499 ( .C (clk), .D (signal_8044), .Q (signal_8045) ) ;
    buf_clk cell_5515 ( .C (clk), .D (signal_8060), .Q (signal_8061) ) ;
    buf_clk cell_5531 ( .C (clk), .D (signal_8076), .Q (signal_8077) ) ;
    buf_clk cell_5547 ( .C (clk), .D (signal_8092), .Q (signal_8093) ) ;
    buf_clk cell_5563 ( .C (clk), .D (signal_8108), .Q (signal_8109) ) ;
    buf_clk cell_5579 ( .C (clk), .D (signal_8124), .Q (signal_8125) ) ;
    buf_clk cell_5595 ( .C (clk), .D (signal_8140), .Q (signal_8141) ) ;
    buf_clk cell_5611 ( .C (clk), .D (signal_8156), .Q (signal_8157) ) ;
    buf_clk cell_5627 ( .C (clk), .D (signal_8172), .Q (signal_8173) ) ;
    buf_clk cell_5643 ( .C (clk), .D (signal_8188), .Q (signal_8189) ) ;
    buf_clk cell_5659 ( .C (clk), .D (signal_8204), .Q (signal_8205) ) ;
    buf_clk cell_5675 ( .C (clk), .D (signal_8220), .Q (signal_8221) ) ;
    buf_clk cell_5691 ( .C (clk), .D (signal_8236), .Q (signal_8237) ) ;
    buf_clk cell_5707 ( .C (clk), .D (signal_8252), .Q (signal_8253) ) ;
    buf_clk cell_5723 ( .C (clk), .D (signal_8268), .Q (signal_8269) ) ;
    buf_clk cell_5739 ( .C (clk), .D (signal_8284), .Q (signal_8285) ) ;
    buf_clk cell_5755 ( .C (clk), .D (signal_8300), .Q (signal_8301) ) ;
    buf_clk cell_5771 ( .C (clk), .D (signal_8316), .Q (signal_8317) ) ;
    buf_clk cell_5787 ( .C (clk), .D (signal_8332), .Q (signal_8333) ) ;
    buf_clk cell_5803 ( .C (clk), .D (signal_8348), .Q (signal_8349) ) ;
    buf_clk cell_5819 ( .C (clk), .D (signal_8364), .Q (signal_8365) ) ;
    buf_clk cell_5835 ( .C (clk), .D (signal_8380), .Q (signal_8381) ) ;
    buf_clk cell_5851 ( .C (clk), .D (signal_8396), .Q (signal_8397) ) ;
    buf_clk cell_5867 ( .C (clk), .D (signal_8412), .Q (signal_8413) ) ;
    buf_clk cell_5883 ( .C (clk), .D (signal_8428), .Q (signal_8429) ) ;
    buf_clk cell_5899 ( .C (clk), .D (signal_8444), .Q (signal_8445) ) ;
    buf_clk cell_5915 ( .C (clk), .D (signal_8460), .Q (signal_8461) ) ;
    buf_clk cell_5931 ( .C (clk), .D (signal_8476), .Q (signal_8477) ) ;
    buf_clk cell_5947 ( .C (clk), .D (signal_8492), .Q (signal_8493) ) ;
    buf_clk cell_5963 ( .C (clk), .D (signal_8508), .Q (signal_8509) ) ;
    buf_clk cell_5979 ( .C (clk), .D (signal_8524), .Q (signal_8525) ) ;
    buf_clk cell_5995 ( .C (clk), .D (signal_8540), .Q (signal_8541) ) ;
    buf_clk cell_6011 ( .C (clk), .D (signal_8556), .Q (signal_8557) ) ;
    buf_clk cell_6027 ( .C (clk), .D (signal_8572), .Q (signal_8573) ) ;
    buf_clk cell_6043 ( .C (clk), .D (signal_8588), .Q (signal_8589) ) ;
    buf_clk cell_6059 ( .C (clk), .D (signal_8604), .Q (signal_8605) ) ;
    buf_clk cell_6075 ( .C (clk), .D (signal_8620), .Q (signal_8621) ) ;
    buf_clk cell_6091 ( .C (clk), .D (signal_8636), .Q (signal_8637) ) ;
    buf_clk cell_6107 ( .C (clk), .D (signal_8652), .Q (signal_8653) ) ;
    buf_clk cell_6123 ( .C (clk), .D (signal_8668), .Q (signal_8669) ) ;
    buf_clk cell_6139 ( .C (clk), .D (signal_8684), .Q (signal_8685) ) ;
    buf_clk cell_6155 ( .C (clk), .D (signal_8700), .Q (signal_8701) ) ;
    buf_clk cell_6171 ( .C (clk), .D (signal_8716), .Q (signal_8717) ) ;
    buf_clk cell_6187 ( .C (clk), .D (signal_8732), .Q (signal_8733) ) ;
    buf_clk cell_6203 ( .C (clk), .D (signal_8748), .Q (signal_8749) ) ;
    buf_clk cell_6219 ( .C (clk), .D (signal_8764), .Q (signal_8765) ) ;
    buf_clk cell_6235 ( .C (clk), .D (signal_8780), .Q (signal_8781) ) ;
    buf_clk cell_6251 ( .C (clk), .D (signal_8796), .Q (signal_8797) ) ;
    buf_clk cell_6267 ( .C (clk), .D (signal_8812), .Q (signal_8813) ) ;
    buf_clk cell_6283 ( .C (clk), .D (signal_8828), .Q (signal_8829) ) ;
    buf_clk cell_6299 ( .C (clk), .D (signal_8844), .Q (signal_8845) ) ;
    buf_clk cell_6315 ( .C (clk), .D (signal_8860), .Q (signal_8861) ) ;
    buf_clk cell_6331 ( .C (clk), .D (signal_8876), .Q (signal_8877) ) ;
    buf_clk cell_6347 ( .C (clk), .D (signal_8892), .Q (signal_8893) ) ;
    buf_clk cell_6363 ( .C (clk), .D (signal_8908), .Q (signal_8909) ) ;
    buf_clk cell_6379 ( .C (clk), .D (signal_8924), .Q (signal_8925) ) ;
    buf_clk cell_6395 ( .C (clk), .D (signal_8940), .Q (signal_8941) ) ;
    buf_clk cell_6411 ( .C (clk), .D (signal_8956), .Q (signal_8957) ) ;
    buf_clk cell_6427 ( .C (clk), .D (signal_8972), .Q (signal_8973) ) ;
    buf_clk cell_6443 ( .C (clk), .D (signal_8988), .Q (signal_8989) ) ;
    buf_clk cell_6459 ( .C (clk), .D (signal_9004), .Q (signal_9005) ) ;
    buf_clk cell_6475 ( .C (clk), .D (signal_9020), .Q (signal_9021) ) ;
    buf_clk cell_6491 ( .C (clk), .D (signal_9036), .Q (signal_9037) ) ;
    buf_clk cell_6507 ( .C (clk), .D (signal_9052), .Q (signal_9053) ) ;
    buf_clk cell_6523 ( .C (clk), .D (signal_9068), .Q (signal_9069) ) ;
    buf_clk cell_6539 ( .C (clk), .D (signal_9084), .Q (signal_9085) ) ;
    buf_clk cell_6555 ( .C (clk), .D (signal_9100), .Q (signal_9101) ) ;
    buf_clk cell_6571 ( .C (clk), .D (signal_9116), .Q (signal_9117) ) ;
    buf_clk cell_6587 ( .C (clk), .D (signal_9132), .Q (signal_9133) ) ;
    buf_clk cell_6603 ( .C (clk), .D (signal_9148), .Q (signal_9149) ) ;
    buf_clk cell_6619 ( .C (clk), .D (signal_9164), .Q (signal_9165) ) ;
    buf_clk cell_6635 ( .C (clk), .D (signal_9180), .Q (signal_9181) ) ;
    buf_clk cell_6651 ( .C (clk), .D (signal_9196), .Q (signal_9197) ) ;
    buf_clk cell_6667 ( .C (clk), .D (signal_9212), .Q (signal_9213) ) ;
    buf_clk cell_6683 ( .C (clk), .D (signal_9228), .Q (signal_9229) ) ;
    buf_clk cell_6699 ( .C (clk), .D (signal_9244), .Q (signal_9245) ) ;
    buf_clk cell_6715 ( .C (clk), .D (signal_9260), .Q (signal_9261) ) ;
    buf_clk cell_6731 ( .C (clk), .D (signal_9276), .Q (signal_9277) ) ;
    buf_clk cell_6747 ( .C (clk), .D (signal_9292), .Q (signal_9293) ) ;
    buf_clk cell_6763 ( .C (clk), .D (signal_9308), .Q (signal_9309) ) ;
    buf_clk cell_6779 ( .C (clk), .D (signal_9324), .Q (signal_9325) ) ;
    buf_clk cell_6795 ( .C (clk), .D (signal_9340), .Q (signal_9341) ) ;
    buf_clk cell_6811 ( .C (clk), .D (signal_9356), .Q (signal_9357) ) ;
    buf_clk cell_6827 ( .C (clk), .D (signal_9372), .Q (signal_9373) ) ;
    buf_clk cell_6843 ( .C (clk), .D (signal_9388), .Q (signal_9389) ) ;
    buf_clk cell_6859 ( .C (clk), .D (signal_9404), .Q (signal_9405) ) ;
    buf_clk cell_6875 ( .C (clk), .D (signal_9420), .Q (signal_9421) ) ;
    buf_clk cell_6891 ( .C (clk), .D (signal_9436), .Q (signal_9437) ) ;
    buf_clk cell_6907 ( .C (clk), .D (signal_9452), .Q (signal_9453) ) ;
    buf_clk cell_6923 ( .C (clk), .D (signal_9468), .Q (signal_9469) ) ;
    buf_clk cell_6939 ( .C (clk), .D (signal_9484), .Q (signal_9485) ) ;
    buf_clk cell_6955 ( .C (clk), .D (signal_9500), .Q (signal_9501) ) ;
    buf_clk cell_6971 ( .C (clk), .D (signal_9516), .Q (signal_9517) ) ;
    buf_clk cell_6987 ( .C (clk), .D (signal_9532), .Q (signal_9533) ) ;
    buf_clk cell_7003 ( .C (clk), .D (signal_9548), .Q (signal_9549) ) ;
    buf_clk cell_7019 ( .C (clk), .D (signal_9564), .Q (signal_9565) ) ;
    buf_clk cell_7035 ( .C (clk), .D (signal_9580), .Q (signal_9581) ) ;
    buf_clk cell_7051 ( .C (clk), .D (signal_9596), .Q (signal_9597) ) ;
    buf_clk cell_7067 ( .C (clk), .D (signal_9612), .Q (signal_9613) ) ;
    buf_clk cell_7083 ( .C (clk), .D (signal_9628), .Q (signal_9629) ) ;
    buf_clk cell_7099 ( .C (clk), .D (signal_9644), .Q (signal_9645) ) ;
    buf_clk cell_7115 ( .C (clk), .D (signal_9660), .Q (signal_9661) ) ;
    buf_clk cell_7131 ( .C (clk), .D (signal_9676), .Q (signal_9677) ) ;
    buf_clk cell_7147 ( .C (clk), .D (signal_9692), .Q (signal_9693) ) ;
    buf_clk cell_7163 ( .C (clk), .D (signal_9708), .Q (signal_9709) ) ;
    buf_clk cell_7179 ( .C (clk), .D (signal_9724), .Q (signal_9725) ) ;
    buf_clk cell_7195 ( .C (clk), .D (signal_9740), .Q (signal_9741) ) ;
    buf_clk cell_7211 ( .C (clk), .D (signal_9756), .Q (signal_9757) ) ;
    buf_clk cell_7227 ( .C (clk), .D (signal_9772), .Q (signal_9773) ) ;
    buf_clk cell_7243 ( .C (clk), .D (signal_9788), .Q (signal_9789) ) ;
    buf_clk cell_7259 ( .C (clk), .D (signal_9804), .Q (signal_9805) ) ;
    buf_clk cell_7275 ( .C (clk), .D (signal_9820), .Q (signal_9821) ) ;
    buf_clk cell_7291 ( .C (clk), .D (signal_9836), .Q (signal_9837) ) ;
    buf_clk cell_7307 ( .C (clk), .D (signal_9852), .Q (signal_9853) ) ;
    buf_clk cell_7323 ( .C (clk), .D (signal_9868), .Q (signal_9869) ) ;
    buf_clk cell_7339 ( .C (clk), .D (signal_9884), .Q (signal_9885) ) ;
    buf_clk cell_7355 ( .C (clk), .D (signal_9900), .Q (signal_9901) ) ;
    buf_clk cell_7371 ( .C (clk), .D (signal_9916), .Q (signal_9917) ) ;
    buf_clk cell_7387 ( .C (clk), .D (signal_9932), .Q (signal_9933) ) ;
    buf_clk cell_7403 ( .C (clk), .D (signal_9948), .Q (signal_9949) ) ;
    buf_clk cell_7419 ( .C (clk), .D (signal_9964), .Q (signal_9965) ) ;
    buf_clk cell_7435 ( .C (clk), .D (signal_9980), .Q (signal_9981) ) ;
    buf_clk cell_7451 ( .C (clk), .D (signal_9996), .Q (signal_9997) ) ;
    buf_clk cell_7467 ( .C (clk), .D (signal_10012), .Q (signal_10013) ) ;
    buf_clk cell_7483 ( .C (clk), .D (signal_10028), .Q (signal_10029) ) ;
    buf_clk cell_7499 ( .C (clk), .D (signal_10044), .Q (signal_10045) ) ;
    buf_clk cell_7515 ( .C (clk), .D (signal_10060), .Q (signal_10061) ) ;
    buf_clk cell_7531 ( .C (clk), .D (signal_10076), .Q (signal_10077) ) ;
    buf_clk cell_7547 ( .C (clk), .D (signal_10092), .Q (signal_10093) ) ;
    buf_clk cell_7563 ( .C (clk), .D (signal_10108), .Q (signal_10109) ) ;
    buf_clk cell_7579 ( .C (clk), .D (signal_10124), .Q (signal_10125) ) ;
    buf_clk cell_7595 ( .C (clk), .D (signal_10140), .Q (signal_10141) ) ;
    buf_clk cell_7611 ( .C (clk), .D (signal_10156), .Q (signal_10157) ) ;
    buf_clk cell_7627 ( .C (clk), .D (signal_10172), .Q (signal_10173) ) ;
    buf_clk cell_7643 ( .C (clk), .D (signal_10188), .Q (signal_10189) ) ;
    buf_clk cell_7659 ( .C (clk), .D (signal_10204), .Q (signal_10205) ) ;
    buf_clk cell_7675 ( .C (clk), .D (signal_10220), .Q (signal_10221) ) ;
    buf_clk cell_7691 ( .C (clk), .D (signal_10236), .Q (signal_10237) ) ;
    buf_clk cell_7707 ( .C (clk), .D (signal_10252), .Q (signal_10253) ) ;
    buf_clk cell_7723 ( .C (clk), .D (signal_10268), .Q (signal_10269) ) ;
    buf_clk cell_7739 ( .C (clk), .D (signal_10284), .Q (signal_10285) ) ;
    buf_clk cell_7755 ( .C (clk), .D (signal_10300), .Q (signal_10301) ) ;
    buf_clk cell_7771 ( .C (clk), .D (signal_10316), .Q (signal_10317) ) ;
    buf_clk cell_7787 ( .C (clk), .D (signal_10332), .Q (signal_10333) ) ;
    buf_clk cell_7803 ( .C (clk), .D (signal_10348), .Q (signal_10349) ) ;
    buf_clk cell_7819 ( .C (clk), .D (signal_10364), .Q (signal_10365) ) ;
    buf_clk cell_7835 ( .C (clk), .D (signal_10380), .Q (signal_10381) ) ;
    buf_clk cell_7851 ( .C (clk), .D (signal_10396), .Q (signal_10397) ) ;
    buf_clk cell_7867 ( .C (clk), .D (signal_10412), .Q (signal_10413) ) ;
    buf_clk cell_7883 ( .C (clk), .D (signal_10428), .Q (signal_10429) ) ;
    buf_clk cell_7899 ( .C (clk), .D (signal_10444), .Q (signal_10445) ) ;
    buf_clk cell_7915 ( .C (clk), .D (signal_10460), .Q (signal_10461) ) ;
    buf_clk cell_7931 ( .C (clk), .D (signal_10476), .Q (signal_10477) ) ;
    buf_clk cell_7947 ( .C (clk), .D (signal_10492), .Q (signal_10493) ) ;
    buf_clk cell_7963 ( .C (clk), .D (signal_10508), .Q (signal_10509) ) ;
    buf_clk cell_7979 ( .C (clk), .D (signal_10524), .Q (signal_10525) ) ;
    buf_clk cell_7995 ( .C (clk), .D (signal_10540), .Q (signal_10541) ) ;
    buf_clk cell_8011 ( .C (clk), .D (signal_10556), .Q (signal_10557) ) ;
    buf_clk cell_8027 ( .C (clk), .D (signal_10572), .Q (signal_10573) ) ;
    buf_clk cell_8043 ( .C (clk), .D (signal_10588), .Q (signal_10589) ) ;
    buf_clk cell_8059 ( .C (clk), .D (signal_10604), .Q (signal_10605) ) ;
    buf_clk cell_8075 ( .C (clk), .D (signal_10620), .Q (signal_10621) ) ;
    buf_clk cell_8091 ( .C (clk), .D (signal_10636), .Q (signal_10637) ) ;
    buf_clk cell_8107 ( .C (clk), .D (signal_10652), .Q (signal_10653) ) ;
    buf_clk cell_8123 ( .C (clk), .D (signal_10668), .Q (signal_10669) ) ;
    buf_clk cell_8139 ( .C (clk), .D (signal_10684), .Q (signal_10685) ) ;
    buf_clk cell_8155 ( .C (clk), .D (signal_10700), .Q (signal_10701) ) ;
    buf_clk cell_8171 ( .C (clk), .D (signal_10716), .Q (signal_10717) ) ;
    buf_clk cell_8187 ( .C (clk), .D (signal_10732), .Q (signal_10733) ) ;
    buf_clk cell_8203 ( .C (clk), .D (signal_10748), .Q (signal_10749) ) ;
    buf_clk cell_8219 ( .C (clk), .D (signal_10764), .Q (signal_10765) ) ;
    buf_clk cell_8235 ( .C (clk), .D (signal_10780), .Q (signal_10781) ) ;
    buf_clk cell_8251 ( .C (clk), .D (signal_10796), .Q (signal_10797) ) ;
    buf_clk cell_8267 ( .C (clk), .D (signal_10812), .Q (signal_10813) ) ;
    buf_clk cell_8283 ( .C (clk), .D (signal_10828), .Q (signal_10829) ) ;
    buf_clk cell_8299 ( .C (clk), .D (signal_10844), .Q (signal_10845) ) ;
    buf_clk cell_8315 ( .C (clk), .D (signal_10860), .Q (signal_10861) ) ;
    buf_clk cell_8331 ( .C (clk), .D (signal_10876), .Q (signal_10877) ) ;
    buf_clk cell_8347 ( .C (clk), .D (signal_10892), .Q (signal_10893) ) ;
    buf_clk cell_8363 ( .C (clk), .D (signal_10908), .Q (signal_10909) ) ;
    buf_clk cell_8379 ( .C (clk), .D (signal_10924), .Q (signal_10925) ) ;
    buf_clk cell_8395 ( .C (clk), .D (signal_10940), .Q (signal_10941) ) ;
    buf_clk cell_8411 ( .C (clk), .D (signal_10956), .Q (signal_10957) ) ;
    buf_clk cell_8427 ( .C (clk), .D (signal_10972), .Q (signal_10973) ) ;
    buf_clk cell_8443 ( .C (clk), .D (signal_10988), .Q (signal_10989) ) ;
    buf_clk cell_8459 ( .C (clk), .D (signal_11004), .Q (signal_11005) ) ;
    buf_clk cell_8475 ( .C (clk), .D (signal_11020), .Q (signal_11021) ) ;
    buf_clk cell_8491 ( .C (clk), .D (signal_11036), .Q (signal_11037) ) ;
    buf_clk cell_8507 ( .C (clk), .D (signal_11052), .Q (signal_11053) ) ;
    buf_clk cell_8523 ( .C (clk), .D (signal_11068), .Q (signal_11069) ) ;
    buf_clk cell_8539 ( .C (clk), .D (signal_11084), .Q (signal_11085) ) ;
    buf_clk cell_8555 ( .C (clk), .D (signal_11100), .Q (signal_11101) ) ;
    buf_clk cell_8571 ( .C (clk), .D (signal_11116), .Q (signal_11117) ) ;
    buf_clk cell_8587 ( .C (clk), .D (signal_11132), .Q (signal_11133) ) ;
    buf_clk cell_8603 ( .C (clk), .D (signal_11148), .Q (signal_11149) ) ;
    buf_clk cell_8619 ( .C (clk), .D (signal_11164), .Q (signal_11165) ) ;
    buf_clk cell_8635 ( .C (clk), .D (signal_11180), .Q (signal_11181) ) ;
    buf_clk cell_8651 ( .C (clk), .D (signal_11196), .Q (signal_11197) ) ;
    buf_clk cell_8667 ( .C (clk), .D (signal_11212), .Q (signal_11213) ) ;
    buf_clk cell_8683 ( .C (clk), .D (signal_11228), .Q (signal_11229) ) ;
    buf_clk cell_8699 ( .C (clk), .D (signal_11244), .Q (signal_11245) ) ;
    buf_clk cell_8715 ( .C (clk), .D (signal_11260), .Q (signal_11261) ) ;
    buf_clk cell_8731 ( .C (clk), .D (signal_11276), .Q (signal_11277) ) ;
    buf_clk cell_8747 ( .C (clk), .D (signal_11292), .Q (signal_11293) ) ;
    buf_clk cell_8763 ( .C (clk), .D (signal_11308), .Q (signal_11309) ) ;
    buf_clk cell_8779 ( .C (clk), .D (signal_11324), .Q (signal_11325) ) ;
    buf_clk cell_8795 ( .C (clk), .D (signal_11340), .Q (signal_11341) ) ;
    buf_clk cell_8811 ( .C (clk), .D (signal_11356), .Q (signal_11357) ) ;
    buf_clk cell_8827 ( .C (clk), .D (signal_11372), .Q (signal_11373) ) ;
    buf_clk cell_8843 ( .C (clk), .D (signal_11388), .Q (signal_11389) ) ;
    buf_clk cell_8859 ( .C (clk), .D (signal_11404), .Q (signal_11405) ) ;
    buf_clk cell_8875 ( .C (clk), .D (signal_11420), .Q (signal_11421) ) ;
    buf_clk cell_8891 ( .C (clk), .D (signal_11436), .Q (signal_11437) ) ;
    buf_clk cell_8907 ( .C (clk), .D (signal_11452), .Q (signal_11453) ) ;
    buf_clk cell_8923 ( .C (clk), .D (signal_11468), .Q (signal_11469) ) ;
    buf_clk cell_8939 ( .C (clk), .D (signal_11484), .Q (signal_11485) ) ;
    buf_clk cell_8955 ( .C (clk), .D (signal_11500), .Q (signal_11501) ) ;
    buf_clk cell_8971 ( .C (clk), .D (signal_11516), .Q (signal_11517) ) ;
    buf_clk cell_8987 ( .C (clk), .D (signal_11532), .Q (signal_11533) ) ;
    buf_clk cell_9003 ( .C (clk), .D (signal_11548), .Q (signal_11549) ) ;
    buf_clk cell_9019 ( .C (clk), .D (signal_11564), .Q (signal_11565) ) ;
    buf_clk cell_9035 ( .C (clk), .D (signal_11580), .Q (signal_11581) ) ;
    buf_clk cell_9051 ( .C (clk), .D (signal_11596), .Q (signal_11597) ) ;
    buf_clk cell_9067 ( .C (clk), .D (signal_11612), .Q (signal_11613) ) ;
    buf_clk cell_9083 ( .C (clk), .D (signal_11628), .Q (signal_11629) ) ;
    buf_clk cell_9099 ( .C (clk), .D (signal_11644), .Q (signal_11645) ) ;
    buf_clk cell_9115 ( .C (clk), .D (signal_11660), .Q (signal_11661) ) ;
    buf_clk cell_9131 ( .C (clk), .D (signal_11676), .Q (signal_11677) ) ;
    buf_clk cell_9147 ( .C (clk), .D (signal_11692), .Q (signal_11693) ) ;
    buf_clk cell_9163 ( .C (clk), .D (signal_11708), .Q (signal_11709) ) ;
    buf_clk cell_9179 ( .C (clk), .D (signal_11724), .Q (signal_11725) ) ;
    buf_clk cell_9195 ( .C (clk), .D (signal_11740), .Q (signal_11741) ) ;
    buf_clk cell_9211 ( .C (clk), .D (signal_11756), .Q (signal_11757) ) ;
    buf_clk cell_9227 ( .C (clk), .D (signal_11772), .Q (signal_11773) ) ;
    buf_clk cell_9243 ( .C (clk), .D (signal_11788), .Q (signal_11789) ) ;
    buf_clk cell_9259 ( .C (clk), .D (signal_11804), .Q (signal_11805) ) ;
    buf_clk cell_9275 ( .C (clk), .D (signal_11820), .Q (signal_11821) ) ;
    buf_clk cell_9291 ( .C (clk), .D (signal_11836), .Q (signal_11837) ) ;
    buf_clk cell_9307 ( .C (clk), .D (signal_11852), .Q (signal_11853) ) ;
    buf_clk cell_9323 ( .C (clk), .D (signal_11868), .Q (signal_11869) ) ;
    buf_clk cell_9339 ( .C (clk), .D (signal_11884), .Q (signal_11885) ) ;
    buf_clk cell_9355 ( .C (clk), .D (signal_11900), .Q (signal_11901) ) ;
    buf_clk cell_9371 ( .C (clk), .D (signal_11916), .Q (signal_11917) ) ;
    buf_clk cell_9387 ( .C (clk), .D (signal_11932), .Q (signal_11933) ) ;
    buf_clk cell_9403 ( .C (clk), .D (signal_11948), .Q (signal_11949) ) ;
    buf_clk cell_9419 ( .C (clk), .D (signal_11964), .Q (signal_11965) ) ;
    buf_clk cell_9435 ( .C (clk), .D (signal_11980), .Q (signal_11981) ) ;
    buf_clk cell_9451 ( .C (clk), .D (signal_11996), .Q (signal_11997) ) ;
    buf_clk cell_9467 ( .C (clk), .D (signal_12012), .Q (signal_12013) ) ;
    buf_clk cell_9483 ( .C (clk), .D (signal_12028), .Q (signal_12029) ) ;
    buf_clk cell_9499 ( .C (clk), .D (signal_12044), .Q (signal_12045) ) ;
    buf_clk cell_9515 ( .C (clk), .D (signal_12060), .Q (signal_12061) ) ;
    buf_clk cell_9531 ( .C (clk), .D (signal_12076), .Q (signal_12077) ) ;
    buf_clk cell_9547 ( .C (clk), .D (signal_12092), .Q (signal_12093) ) ;
    buf_clk cell_9563 ( .C (clk), .D (signal_12108), .Q (signal_12109) ) ;
    buf_clk cell_9579 ( .C (clk), .D (signal_12124), .Q (signal_12125) ) ;
    buf_clk cell_9595 ( .C (clk), .D (signal_12140), .Q (signal_12141) ) ;
    buf_clk cell_9611 ( .C (clk), .D (signal_12156), .Q (signal_12157) ) ;
    buf_clk cell_9627 ( .C (clk), .D (signal_12172), .Q (signal_12173) ) ;
    buf_clk cell_9643 ( .C (clk), .D (signal_12188), .Q (signal_12189) ) ;
    buf_clk cell_9659 ( .C (clk), .D (signal_12204), .Q (signal_12205) ) ;
    buf_clk cell_9675 ( .C (clk), .D (signal_12220), .Q (signal_12221) ) ;
    buf_clk cell_9691 ( .C (clk), .D (signal_12236), .Q (signal_12237) ) ;
    buf_clk cell_9707 ( .C (clk), .D (signal_12252), .Q (signal_12253) ) ;
    buf_clk cell_9723 ( .C (clk), .D (signal_12268), .Q (signal_12269) ) ;
    buf_clk cell_9739 ( .C (clk), .D (signal_12284), .Q (signal_12285) ) ;
    buf_clk cell_9755 ( .C (clk), .D (signal_12300), .Q (signal_12301) ) ;
    buf_clk cell_9771 ( .C (clk), .D (signal_12316), .Q (signal_12317) ) ;
    buf_clk cell_9787 ( .C (clk), .D (signal_12332), .Q (signal_12333) ) ;
    buf_clk cell_9803 ( .C (clk), .D (signal_12348), .Q (signal_12349) ) ;
    buf_clk cell_9819 ( .C (clk), .D (signal_12364), .Q (signal_12365) ) ;
    buf_clk cell_9835 ( .C (clk), .D (signal_12380), .Q (signal_12381) ) ;
    buf_clk cell_9851 ( .C (clk), .D (signal_12396), .Q (signal_12397) ) ;
    buf_clk cell_9867 ( .C (clk), .D (signal_12412), .Q (signal_12413) ) ;
    buf_clk cell_9883 ( .C (clk), .D (signal_12428), .Q (signal_12429) ) ;
    buf_clk cell_9899 ( .C (clk), .D (signal_12444), .Q (signal_12445) ) ;
    buf_clk cell_9915 ( .C (clk), .D (signal_12460), .Q (signal_12461) ) ;
    buf_clk cell_9931 ( .C (clk), .D (signal_12476), .Q (signal_12477) ) ;
    buf_clk cell_9947 ( .C (clk), .D (signal_12492), .Q (signal_12493) ) ;
    buf_clk cell_9963 ( .C (clk), .D (signal_12508), .Q (signal_12509) ) ;
    buf_clk cell_9979 ( .C (clk), .D (signal_12524), .Q (signal_12525) ) ;
    buf_clk cell_9995 ( .C (clk), .D (signal_12540), .Q (signal_12541) ) ;
    buf_clk cell_10011 ( .C (clk), .D (signal_12556), .Q (signal_12557) ) ;
    buf_clk cell_10027 ( .C (clk), .D (signal_12572), .Q (signal_12573) ) ;
    buf_clk cell_10043 ( .C (clk), .D (signal_12588), .Q (signal_12589) ) ;
    buf_clk cell_10059 ( .C (clk), .D (signal_12604), .Q (signal_12605) ) ;
    buf_clk cell_10075 ( .C (clk), .D (signal_12620), .Q (signal_12621) ) ;
    buf_clk cell_10091 ( .C (clk), .D (signal_12636), .Q (signal_12637) ) ;
    buf_clk cell_10107 ( .C (clk), .D (signal_12652), .Q (signal_12653) ) ;
    buf_clk cell_10123 ( .C (clk), .D (signal_12668), .Q (signal_12669) ) ;
    buf_clk cell_10139 ( .C (clk), .D (signal_12684), .Q (signal_12685) ) ;
    buf_clk cell_10155 ( .C (clk), .D (signal_12700), .Q (signal_12701) ) ;
    buf_clk cell_10171 ( .C (clk), .D (signal_12716), .Q (signal_12717) ) ;
    buf_clk cell_10187 ( .C (clk), .D (signal_12732), .Q (signal_12733) ) ;
    buf_clk cell_10203 ( .C (clk), .D (signal_12748), .Q (signal_12749) ) ;
    buf_clk cell_10219 ( .C (clk), .D (signal_12764), .Q (signal_12765) ) ;
    buf_clk cell_10235 ( .C (clk), .D (signal_12780), .Q (signal_12781) ) ;
    buf_clk cell_10251 ( .C (clk), .D (signal_12796), .Q (signal_12797) ) ;
    buf_clk cell_10267 ( .C (clk), .D (signal_12812), .Q (signal_12813) ) ;
    buf_clk cell_10283 ( .C (clk), .D (signal_12828), .Q (signal_12829) ) ;
    buf_clk cell_10299 ( .C (clk), .D (signal_12844), .Q (signal_12845) ) ;
    buf_clk cell_10315 ( .C (clk), .D (signal_12860), .Q (signal_12861) ) ;
    buf_clk cell_10331 ( .C (clk), .D (signal_12876), .Q (signal_12877) ) ;
    buf_clk cell_10347 ( .C (clk), .D (signal_12892), .Q (signal_12893) ) ;
    buf_clk cell_10363 ( .C (clk), .D (signal_12908), .Q (signal_12909) ) ;
    buf_clk cell_10379 ( .C (clk), .D (signal_12924), .Q (signal_12925) ) ;
    buf_clk cell_10395 ( .C (clk), .D (signal_12940), .Q (signal_12941) ) ;
    buf_clk cell_10411 ( .C (clk), .D (signal_12956), .Q (signal_12957) ) ;
    buf_clk cell_10427 ( .C (clk), .D (signal_12972), .Q (signal_12973) ) ;
    buf_clk cell_10443 ( .C (clk), .D (signal_12988), .Q (signal_12989) ) ;
    buf_clk cell_10459 ( .C (clk), .D (signal_13004), .Q (signal_13005) ) ;
    buf_clk cell_10475 ( .C (clk), .D (signal_13020), .Q (signal_13021) ) ;
    buf_clk cell_10491 ( .C (clk), .D (signal_13036), .Q (signal_13037) ) ;
    buf_clk cell_10507 ( .C (clk), .D (signal_13052), .Q (signal_13053) ) ;
    buf_clk cell_10523 ( .C (clk), .D (signal_13068), .Q (signal_13069) ) ;
    buf_clk cell_10539 ( .C (clk), .D (signal_13084), .Q (signal_13085) ) ;
    buf_clk cell_10555 ( .C (clk), .D (signal_13100), .Q (signal_13101) ) ;
    buf_clk cell_10571 ( .C (clk), .D (signal_13116), .Q (signal_13117) ) ;
    buf_clk cell_10587 ( .C (clk), .D (signal_13132), .Q (signal_13133) ) ;
    buf_clk cell_10603 ( .C (clk), .D (signal_13148), .Q (signal_13149) ) ;
    buf_clk cell_10619 ( .C (clk), .D (signal_13164), .Q (signal_13165) ) ;
    buf_clk cell_10635 ( .C (clk), .D (signal_13180), .Q (signal_13181) ) ;
    buf_clk cell_10651 ( .C (clk), .D (signal_13196), .Q (signal_13197) ) ;
    buf_clk cell_10667 ( .C (clk), .D (signal_13212), .Q (signal_13213) ) ;
    buf_clk cell_10683 ( .C (clk), .D (signal_13228), .Q (signal_13229) ) ;
    buf_clk cell_10699 ( .C (clk), .D (signal_13244), .Q (signal_13245) ) ;
    buf_clk cell_10715 ( .C (clk), .D (signal_13260), .Q (signal_13261) ) ;
    buf_clk cell_10731 ( .C (clk), .D (signal_13276), .Q (signal_13277) ) ;
    buf_clk cell_10747 ( .C (clk), .D (signal_13292), .Q (signal_13293) ) ;
    buf_clk cell_10763 ( .C (clk), .D (signal_13308), .Q (signal_13309) ) ;
    buf_clk cell_10779 ( .C (clk), .D (signal_13324), .Q (signal_13325) ) ;
    buf_clk cell_10795 ( .C (clk), .D (signal_13340), .Q (signal_13341) ) ;
    buf_clk cell_10811 ( .C (clk), .D (signal_13356), .Q (signal_13357) ) ;
    buf_clk cell_10827 ( .C (clk), .D (signal_13372), .Q (signal_13373) ) ;
    buf_clk cell_10843 ( .C (clk), .D (signal_13388), .Q (signal_13389) ) ;
    buf_clk cell_10859 ( .C (clk), .D (signal_13404), .Q (signal_13405) ) ;
    buf_clk cell_10875 ( .C (clk), .D (signal_13420), .Q (signal_13421) ) ;
    buf_clk cell_10891 ( .C (clk), .D (signal_13436), .Q (signal_13437) ) ;
    buf_clk cell_10907 ( .C (clk), .D (signal_13452), .Q (signal_13453) ) ;
    buf_clk cell_10923 ( .C (clk), .D (signal_13468), .Q (signal_13469) ) ;
    buf_clk cell_10939 ( .C (clk), .D (signal_13484), .Q (signal_13485) ) ;
    buf_clk cell_10955 ( .C (clk), .D (signal_13500), .Q (signal_13501) ) ;
    buf_clk cell_10971 ( .C (clk), .D (signal_13516), .Q (signal_13517) ) ;
    buf_clk cell_10987 ( .C (clk), .D (signal_13532), .Q (signal_13533) ) ;
    buf_clk cell_11003 ( .C (clk), .D (signal_13548), .Q (signal_13549) ) ;
    buf_clk cell_11019 ( .C (clk), .D (signal_13564), .Q (signal_13565) ) ;
    buf_clk cell_11035 ( .C (clk), .D (signal_13580), .Q (signal_13581) ) ;
    buf_clk cell_11051 ( .C (clk), .D (signal_13596), .Q (signal_13597) ) ;
    buf_clk cell_11067 ( .C (clk), .D (signal_13612), .Q (signal_13613) ) ;
    buf_clk cell_11083 ( .C (clk), .D (signal_13628), .Q (signal_13629) ) ;
    buf_clk cell_11099 ( .C (clk), .D (signal_13644), .Q (signal_13645) ) ;
    buf_clk cell_11115 ( .C (clk), .D (signal_13660), .Q (signal_13661) ) ;
    buf_clk cell_11131 ( .C (clk), .D (signal_13676), .Q (signal_13677) ) ;
    buf_clk cell_11147 ( .C (clk), .D (signal_13692), .Q (signal_13693) ) ;
    buf_clk cell_11163 ( .C (clk), .D (signal_13708), .Q (signal_13709) ) ;
    buf_clk cell_11179 ( .C (clk), .D (signal_13724), .Q (signal_13725) ) ;
    buf_clk cell_11195 ( .C (clk), .D (signal_13740), .Q (signal_13741) ) ;
    buf_clk cell_11211 ( .C (clk), .D (signal_13756), .Q (signal_13757) ) ;
    buf_clk cell_11227 ( .C (clk), .D (signal_13772), .Q (signal_13773) ) ;
    buf_clk cell_11243 ( .C (clk), .D (signal_13788), .Q (signal_13789) ) ;
    buf_clk cell_11259 ( .C (clk), .D (signal_13804), .Q (signal_13805) ) ;
    buf_clk cell_11275 ( .C (clk), .D (signal_13820), .Q (signal_13821) ) ;
    buf_clk cell_11291 ( .C (clk), .D (signal_13836), .Q (signal_13837) ) ;
    buf_clk cell_11307 ( .C (clk), .D (signal_13852), .Q (signal_13853) ) ;
    buf_clk cell_11323 ( .C (clk), .D (signal_13868), .Q (signal_13869) ) ;
    buf_clk cell_11339 ( .C (clk), .D (signal_13884), .Q (signal_13885) ) ;
    buf_clk cell_11355 ( .C (clk), .D (signal_13900), .Q (signal_13901) ) ;
    buf_clk cell_11371 ( .C (clk), .D (signal_13916), .Q (signal_13917) ) ;
    buf_clk cell_11387 ( .C (clk), .D (signal_13932), .Q (signal_13933) ) ;
    buf_clk cell_11403 ( .C (clk), .D (signal_13948), .Q (signal_13949) ) ;
    buf_clk cell_11419 ( .C (clk), .D (signal_13964), .Q (signal_13965) ) ;
    buf_clk cell_11435 ( .C (clk), .D (signal_13980), .Q (signal_13981) ) ;
    buf_clk cell_11451 ( .C (clk), .D (signal_13996), .Q (signal_13997) ) ;
    buf_clk cell_11467 ( .C (clk), .D (signal_14012), .Q (signal_14013) ) ;
    buf_clk cell_11483 ( .C (clk), .D (signal_14028), .Q (signal_14029) ) ;
    buf_clk cell_11499 ( .C (clk), .D (signal_14044), .Q (signal_14045) ) ;
    buf_clk cell_11515 ( .C (clk), .D (signal_14060), .Q (signal_14061) ) ;
    buf_clk cell_11531 ( .C (clk), .D (signal_14076), .Q (signal_14077) ) ;
    buf_clk cell_11547 ( .C (clk), .D (signal_14092), .Q (signal_14093) ) ;
    buf_clk cell_11563 ( .C (clk), .D (signal_14108), .Q (signal_14109) ) ;
    buf_clk cell_11579 ( .C (clk), .D (signal_14124), .Q (signal_14125) ) ;
    buf_clk cell_11595 ( .C (clk), .D (signal_14140), .Q (signal_14141) ) ;
    buf_clk cell_11611 ( .C (clk), .D (signal_14156), .Q (signal_14157) ) ;
    buf_clk cell_11627 ( .C (clk), .D (signal_14172), .Q (signal_14173) ) ;
    buf_clk cell_11643 ( .C (clk), .D (signal_14188), .Q (signal_14189) ) ;
    buf_clk cell_11659 ( .C (clk), .D (signal_14204), .Q (signal_14205) ) ;
    buf_clk cell_11675 ( .C (clk), .D (signal_14220), .Q (signal_14221) ) ;
    buf_clk cell_11691 ( .C (clk), .D (signal_14236), .Q (signal_14237) ) ;
    buf_clk cell_11707 ( .C (clk), .D (signal_14252), .Q (signal_14253) ) ;
    buf_clk cell_11723 ( .C (clk), .D (signal_14268), .Q (signal_14269) ) ;
    buf_clk cell_11739 ( .C (clk), .D (signal_14284), .Q (signal_14285) ) ;
    buf_clk cell_11755 ( .C (clk), .D (signal_14300), .Q (signal_14301) ) ;
    buf_clk cell_11771 ( .C (clk), .D (signal_14316), .Q (signal_14317) ) ;
    buf_clk cell_11787 ( .C (clk), .D (signal_14332), .Q (signal_14333) ) ;
    buf_clk cell_11803 ( .C (clk), .D (signal_14348), .Q (signal_14349) ) ;
    buf_clk cell_11819 ( .C (clk), .D (signal_14364), .Q (signal_14365) ) ;
    buf_clk cell_11835 ( .C (clk), .D (signal_14380), .Q (signal_14381) ) ;
    buf_clk cell_11851 ( .C (clk), .D (signal_14396), .Q (signal_14397) ) ;
    buf_clk cell_11867 ( .C (clk), .D (signal_14412), .Q (signal_14413) ) ;
    buf_clk cell_11883 ( .C (clk), .D (signal_14428), .Q (signal_14429) ) ;
    buf_clk cell_11899 ( .C (clk), .D (signal_14444), .Q (signal_14445) ) ;
    buf_clk cell_11915 ( .C (clk), .D (signal_14460), .Q (signal_14461) ) ;
    buf_clk cell_11931 ( .C (clk), .D (signal_14476), .Q (signal_14477) ) ;
    buf_clk cell_11947 ( .C (clk), .D (signal_14492), .Q (signal_14493) ) ;
    buf_clk cell_11963 ( .C (clk), .D (signal_14508), .Q (signal_14509) ) ;
    buf_clk cell_11979 ( .C (clk), .D (signal_14524), .Q (signal_14525) ) ;
    buf_clk cell_11995 ( .C (clk), .D (signal_14540), .Q (signal_14541) ) ;
    buf_clk cell_12011 ( .C (clk), .D (signal_14556), .Q (signal_14557) ) ;
    buf_clk cell_12027 ( .C (clk), .D (signal_14572), .Q (signal_14573) ) ;
    buf_clk cell_12043 ( .C (clk), .D (signal_14588), .Q (signal_14589) ) ;
    buf_clk cell_12059 ( .C (clk), .D (signal_14604), .Q (signal_14605) ) ;
    buf_clk cell_12075 ( .C (clk), .D (signal_14620), .Q (signal_14621) ) ;
    buf_clk cell_12091 ( .C (clk), .D (signal_14636), .Q (signal_14637) ) ;
    buf_clk cell_12107 ( .C (clk), .D (signal_14652), .Q (signal_14653) ) ;
    buf_clk cell_12123 ( .C (clk), .D (signal_14668), .Q (signal_14669) ) ;
    buf_clk cell_12139 ( .C (clk), .D (signal_14684), .Q (signal_14685) ) ;
    buf_clk cell_12155 ( .C (clk), .D (signal_14700), .Q (signal_14701) ) ;
    buf_clk cell_12171 ( .C (clk), .D (signal_14716), .Q (signal_14717) ) ;
    buf_clk cell_12187 ( .C (clk), .D (signal_14732), .Q (signal_14733) ) ;
    buf_clk cell_12203 ( .C (clk), .D (signal_14748), .Q (signal_14749) ) ;
    buf_clk cell_12219 ( .C (clk), .D (signal_14764), .Q (signal_14765) ) ;
    buf_clk cell_12235 ( .C (clk), .D (signal_14780), .Q (signal_14781) ) ;
    buf_clk cell_12251 ( .C (clk), .D (signal_14796), .Q (signal_14797) ) ;
    buf_clk cell_12267 ( .C (clk), .D (signal_14812), .Q (signal_14813) ) ;
    buf_clk cell_12283 ( .C (clk), .D (signal_14828), .Q (signal_14829) ) ;
    buf_clk cell_12299 ( .C (clk), .D (signal_14844), .Q (signal_14845) ) ;
    buf_clk cell_12315 ( .C (clk), .D (signal_14860), .Q (signal_14861) ) ;
    buf_clk cell_12331 ( .C (clk), .D (signal_14876), .Q (signal_14877) ) ;
    buf_clk cell_12347 ( .C (clk), .D (signal_14892), .Q (signal_14893) ) ;
    buf_clk cell_12363 ( .C (clk), .D (signal_14908), .Q (signal_14909) ) ;
    buf_clk cell_12379 ( .C (clk), .D (signal_14924), .Q (signal_14925) ) ;
    buf_clk cell_12395 ( .C (clk), .D (signal_14940), .Q (signal_14941) ) ;

    /* cells in depth 16 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_56 ( .s (signal_4946), .b ({signal_4180, signal_1405}), .a ({signal_4978, signal_4962}), .c ({signal_4188, signal_1421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_57 ( .s (signal_4946), .b ({signal_4181, signal_1404}), .a ({signal_5010, signal_4994}), .c ({signal_4189, signal_1420}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_58 ( .s (signal_4946), .b ({signal_4182, signal_1403}), .a ({signal_5042, signal_5026}), .c ({signal_4190, signal_1419}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_59 ( .s (signal_4946), .b ({signal_4183, signal_1402}), .a ({signal_5074, signal_5058}), .c ({signal_4191, signal_1418}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_60 ( .s (signal_4946), .b ({signal_4184, signal_1401}), .a ({signal_5106, signal_5090}), .c ({signal_4192, signal_1417}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_61 ( .s (signal_4946), .b ({signal_4185, signal_1400}), .a ({signal_5138, signal_5122}), .c ({signal_4193, signal_1416}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_62 ( .s (signal_4946), .b ({signal_4186, signal_1399}), .a ({signal_5170, signal_5154}), .c ({signal_4194, signal_1415}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_63 ( .s (signal_4946), .b ({signal_4187, signal_1398}), .a ({signal_5202, signal_5186}), .c ({signal_4195, signal_1414}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_445 ( .s (signal_5218), .b ({signal_4221, signal_1557}), .a ({signal_5250, signal_5234}), .c ({signal_4244, signal_705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_448 ( .s (signal_5218), .b ({signal_4223, signal_1556}), .a ({signal_5282, signal_5266}), .c ({signal_4245, signal_707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_451 ( .s (signal_5218), .b ({signal_4225, signal_1555}), .a ({signal_5314, signal_5298}), .c ({signal_4246, signal_709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_454 ( .s (signal_5218), .b ({signal_4227, signal_1554}), .a ({signal_5346, signal_5330}), .c ({signal_4247, signal_711}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_457 ( .s (signal_5218), .b ({signal_4229, signal_1553}), .a ({signal_5378, signal_5362}), .c ({signal_4248, signal_713}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_460 ( .s (signal_5218), .b ({signal_4231, signal_1552}), .a ({signal_5410, signal_5394}), .c ({signal_4249, signal_715}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_463 ( .s (signal_5218), .b ({signal_4233, signal_1551}), .a ({signal_5442, signal_5426}), .c ({signal_4250, signal_717}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_466 ( .s (signal_5218), .b ({signal_4235, signal_1550}), .a ({signal_5474, signal_5458}), .c ({signal_4251, signal_719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_613 ( .s (signal_5490), .b ({signal_4188, signal_1421}), .a ({signal_5522, signal_5506}), .c ({signal_4204, signal_1525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_614 ( .s (signal_5490), .b ({signal_4189, signal_1420}), .a ({signal_5554, signal_5538}), .c ({signal_4205, signal_1524}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_615 ( .s (signal_5490), .b ({signal_4190, signal_1419}), .a ({signal_5586, signal_5570}), .c ({signal_4206, signal_1523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_616 ( .s (signal_5490), .b ({signal_4191, signal_1418}), .a ({signal_5618, signal_5602}), .c ({signal_4207, signal_1522}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_617 ( .s (signal_5490), .b ({signal_4192, signal_1417}), .a ({signal_5650, signal_5634}), .c ({signal_4208, signal_1521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_618 ( .s (signal_5490), .b ({signal_4193, signal_1416}), .a ({signal_5682, signal_5666}), .c ({signal_4209, signal_1520}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_619 ( .s (signal_5490), .b ({signal_4194, signal_1415}), .a ({signal_5714, signal_5698}), .c ({signal_4210, signal_1519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_620 ( .s (signal_5490), .b ({signal_4195, signal_1414}), .a ({signal_5746, signal_5730}), .c ({signal_4211, signal_1518}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_621 ( .s (signal_5762), .b ({signal_5794, signal_5778}), .a ({signal_4204, signal_1525}), .c ({signal_4221, signal_1557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_622 ( .s (signal_5762), .b ({signal_5826, signal_5810}), .a ({signal_4205, signal_1524}), .c ({signal_4223, signal_1556}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_623 ( .s (signal_5762), .b ({signal_5858, signal_5842}), .a ({signal_4206, signal_1523}), .c ({signal_4225, signal_1555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_624 ( .s (signal_5762), .b ({signal_5890, signal_5874}), .a ({signal_4207, signal_1522}), .c ({signal_4227, signal_1554}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_625 ( .s (signal_5762), .b ({signal_5922, signal_5906}), .a ({signal_4208, signal_1521}), .c ({signal_4229, signal_1553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_626 ( .s (signal_5762), .b ({signal_5954, signal_5938}), .a ({signal_4209, signal_1520}), .c ({signal_4231, signal_1552}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_627 ( .s (signal_5762), .b ({signal_5986, signal_5970}), .a ({signal_4210, signal_1519}), .c ({signal_4233, signal_1551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_628 ( .s (signal_5762), .b ({signal_6018, signal_6002}), .a ({signal_4211, signal_1518}), .c ({signal_4235, signal_1550}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_672 ( .a ({signal_4196, signal_724}), .b ({signal_6050, signal_6034}), .c ({signal_4212, signal_1750}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_673 ( .a ({1'b0, signal_6066}), .b ({signal_4187, signal_1398}), .c ({signal_4196, signal_724}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_674 ( .a ({signal_4197, signal_725}), .b ({signal_6098, signal_6082}), .c ({signal_4213, signal_1751}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_675 ( .a ({1'b0, signal_6114}), .b ({signal_4186, signal_1399}), .c ({signal_4197, signal_725}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_676 ( .a ({signal_4198, signal_726}), .b ({signal_6146, signal_6130}), .c ({signal_4214, signal_1752}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_677 ( .a ({1'b0, signal_6162}), .b ({signal_4185, signal_1400}), .c ({signal_4198, signal_726}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_678 ( .a ({signal_4199, signal_727}), .b ({signal_6194, signal_6178}), .c ({signal_4215, signal_1753}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_679 ( .a ({1'b0, signal_6210}), .b ({signal_4184, signal_1401}), .c ({signal_4199, signal_727}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_680 ( .a ({signal_4200, signal_728}), .b ({signal_6242, signal_6226}), .c ({signal_4216, signal_1754}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_681 ( .a ({1'b0, signal_6258}), .b ({signal_4183, signal_1402}), .c ({signal_4200, signal_728}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_682 ( .a ({signal_4201, signal_729}), .b ({signal_6290, signal_6274}), .c ({signal_4217, signal_1755}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_683 ( .a ({1'b0, signal_6306}), .b ({signal_4182, signal_1403}), .c ({signal_4201, signal_729}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_684 ( .a ({signal_4202, signal_730}), .b ({signal_6338, signal_6322}), .c ({signal_4218, signal_1756}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_685 ( .a ({1'b0, signal_6354}), .b ({signal_4181, signal_1404}), .c ({signal_4202, signal_730}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_686 ( .a ({signal_4203, signal_731}), .b ({signal_6386, signal_6370}), .c ({signal_4219, signal_1757}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_687 ( .a ({1'b0, signal_6402}), .b ({signal_4180, signal_1405}), .c ({signal_4203, signal_731}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1098 ( .s (signal_6418), .b ({signal_6450, signal_6434}), .a ({signal_4236, signal_1055}), .c ({signal_4252, signal_1054}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1099 ( .s (signal_6466), .b ({signal_6498, signal_6482}), .a ({signal_4219, signal_1757}), .c ({signal_4236, signal_1055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1102 ( .s (signal_6418), .b ({signal_6530, signal_6514}), .a ({signal_4237, signal_1058}), .c ({signal_4253, signal_1057}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1103 ( .s (signal_6466), .b ({signal_6562, signal_6546}), .a ({signal_4218, signal_1756}), .c ({signal_4237, signal_1058}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1106 ( .s (signal_6418), .b ({signal_6594, signal_6578}), .a ({signal_4238, signal_1061}), .c ({signal_4254, signal_1060}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1107 ( .s (signal_6466), .b ({signal_6626, signal_6610}), .a ({signal_4217, signal_1755}), .c ({signal_4238, signal_1061}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1110 ( .s (signal_6418), .b ({signal_6658, signal_6642}), .a ({signal_4239, signal_1064}), .c ({signal_4255, signal_1063}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1111 ( .s (signal_6466), .b ({signal_6690, signal_6674}), .a ({signal_4216, signal_1754}), .c ({signal_4239, signal_1064}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1114 ( .s (signal_6418), .b ({signal_6722, signal_6706}), .a ({signal_4240, signal_1067}), .c ({signal_4256, signal_1066}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1115 ( .s (signal_6466), .b ({signal_6754, signal_6738}), .a ({signal_4215, signal_1753}), .c ({signal_4240, signal_1067}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1118 ( .s (signal_6418), .b ({signal_6786, signal_6770}), .a ({signal_4241, signal_1070}), .c ({signal_4257, signal_1069}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1119 ( .s (signal_6466), .b ({signal_6818, signal_6802}), .a ({signal_4214, signal_1752}), .c ({signal_4241, signal_1070}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1122 ( .s (signal_6418), .b ({signal_6850, signal_6834}), .a ({signal_4242, signal_1073}), .c ({signal_4258, signal_1072}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1123 ( .s (signal_6466), .b ({signal_6882, signal_6866}), .a ({signal_4213, signal_1751}), .c ({signal_4242, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1126 ( .s (signal_6418), .b ({signal_6914, signal_6898}), .a ({signal_4243, signal_1076}), .c ({signal_4259, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1127 ( .s (signal_6466), .b ({signal_6946, signal_6930}), .a ({signal_4212, signal_1750}), .c ({signal_4243, signal_1076}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2137 ( .s ({signal_6974, signal_6960}), .b ({signal_4165, signal_2390}), .a ({signal_4164, signal_2389}), .clk (clk), .r (Fresh[423]), .c ({signal_4180, signal_1405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2138 ( .s ({signal_6974, signal_6960}), .b ({signal_4167, signal_2392}), .a ({signal_4166, signal_2391}), .clk (clk), .r (Fresh[424]), .c ({signal_4181, signal_1404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2139 ( .s ({signal_6974, signal_6960}), .b ({signal_4169, signal_2394}), .a ({signal_4168, signal_2393}), .clk (clk), .r (Fresh[425]), .c ({signal_4182, signal_1403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2140 ( .s ({signal_6974, signal_6960}), .b ({signal_4171, signal_2396}), .a ({signal_4170, signal_2395}), .clk (clk), .r (Fresh[426]), .c ({signal_4183, signal_1402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2141 ( .s ({signal_6974, signal_6960}), .b ({signal_4173, signal_2398}), .a ({signal_4172, signal_2397}), .clk (clk), .r (Fresh[427]), .c ({signal_4184, signal_1401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2142 ( .s ({signal_6974, signal_6960}), .b ({signal_4175, signal_2400}), .a ({signal_4174, signal_2399}), .clk (clk), .r (Fresh[428]), .c ({signal_4185, signal_1400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2143 ( .s ({signal_6974, signal_6960}), .b ({signal_4177, signal_2402}), .a ({signal_4176, signal_2401}), .clk (clk), .r (Fresh[429]), .c ({signal_4186, signal_1399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_2144 ( .s ({signal_6974, signal_6960}), .b ({signal_4179, signal_2404}), .a ({signal_4178, signal_2403}), .clk (clk), .r (Fresh[430]), .c ({signal_4187, signal_1398}) ) ;
    buf_clk cell_2400 ( .C (clk), .D (signal_4945), .Q (signal_4946) ) ;
    buf_clk cell_2416 ( .C (clk), .D (signal_4961), .Q (signal_4962) ) ;
    buf_clk cell_2432 ( .C (clk), .D (signal_4977), .Q (signal_4978) ) ;
    buf_clk cell_2448 ( .C (clk), .D (signal_4993), .Q (signal_4994) ) ;
    buf_clk cell_2464 ( .C (clk), .D (signal_5009), .Q (signal_5010) ) ;
    buf_clk cell_2480 ( .C (clk), .D (signal_5025), .Q (signal_5026) ) ;
    buf_clk cell_2496 ( .C (clk), .D (signal_5041), .Q (signal_5042) ) ;
    buf_clk cell_2512 ( .C (clk), .D (signal_5057), .Q (signal_5058) ) ;
    buf_clk cell_2528 ( .C (clk), .D (signal_5073), .Q (signal_5074) ) ;
    buf_clk cell_2544 ( .C (clk), .D (signal_5089), .Q (signal_5090) ) ;
    buf_clk cell_2560 ( .C (clk), .D (signal_5105), .Q (signal_5106) ) ;
    buf_clk cell_2576 ( .C (clk), .D (signal_5121), .Q (signal_5122) ) ;
    buf_clk cell_2592 ( .C (clk), .D (signal_5137), .Q (signal_5138) ) ;
    buf_clk cell_2608 ( .C (clk), .D (signal_5153), .Q (signal_5154) ) ;
    buf_clk cell_2624 ( .C (clk), .D (signal_5169), .Q (signal_5170) ) ;
    buf_clk cell_2640 ( .C (clk), .D (signal_5185), .Q (signal_5186) ) ;
    buf_clk cell_2656 ( .C (clk), .D (signal_5201), .Q (signal_5202) ) ;
    buf_clk cell_2672 ( .C (clk), .D (signal_5217), .Q (signal_5218) ) ;
    buf_clk cell_2688 ( .C (clk), .D (signal_5233), .Q (signal_5234) ) ;
    buf_clk cell_2704 ( .C (clk), .D (signal_5249), .Q (signal_5250) ) ;
    buf_clk cell_2720 ( .C (clk), .D (signal_5265), .Q (signal_5266) ) ;
    buf_clk cell_2736 ( .C (clk), .D (signal_5281), .Q (signal_5282) ) ;
    buf_clk cell_2752 ( .C (clk), .D (signal_5297), .Q (signal_5298) ) ;
    buf_clk cell_2768 ( .C (clk), .D (signal_5313), .Q (signal_5314) ) ;
    buf_clk cell_2784 ( .C (clk), .D (signal_5329), .Q (signal_5330) ) ;
    buf_clk cell_2800 ( .C (clk), .D (signal_5345), .Q (signal_5346) ) ;
    buf_clk cell_2816 ( .C (clk), .D (signal_5361), .Q (signal_5362) ) ;
    buf_clk cell_2832 ( .C (clk), .D (signal_5377), .Q (signal_5378) ) ;
    buf_clk cell_2848 ( .C (clk), .D (signal_5393), .Q (signal_5394) ) ;
    buf_clk cell_2864 ( .C (clk), .D (signal_5409), .Q (signal_5410) ) ;
    buf_clk cell_2880 ( .C (clk), .D (signal_5425), .Q (signal_5426) ) ;
    buf_clk cell_2896 ( .C (clk), .D (signal_5441), .Q (signal_5442) ) ;
    buf_clk cell_2912 ( .C (clk), .D (signal_5457), .Q (signal_5458) ) ;
    buf_clk cell_2928 ( .C (clk), .D (signal_5473), .Q (signal_5474) ) ;
    buf_clk cell_2944 ( .C (clk), .D (signal_5489), .Q (signal_5490) ) ;
    buf_clk cell_2960 ( .C (clk), .D (signal_5505), .Q (signal_5506) ) ;
    buf_clk cell_2976 ( .C (clk), .D (signal_5521), .Q (signal_5522) ) ;
    buf_clk cell_2992 ( .C (clk), .D (signal_5537), .Q (signal_5538) ) ;
    buf_clk cell_3008 ( .C (clk), .D (signal_5553), .Q (signal_5554) ) ;
    buf_clk cell_3024 ( .C (clk), .D (signal_5569), .Q (signal_5570) ) ;
    buf_clk cell_3040 ( .C (clk), .D (signal_5585), .Q (signal_5586) ) ;
    buf_clk cell_3056 ( .C (clk), .D (signal_5601), .Q (signal_5602) ) ;
    buf_clk cell_3072 ( .C (clk), .D (signal_5617), .Q (signal_5618) ) ;
    buf_clk cell_3088 ( .C (clk), .D (signal_5633), .Q (signal_5634) ) ;
    buf_clk cell_3104 ( .C (clk), .D (signal_5649), .Q (signal_5650) ) ;
    buf_clk cell_3120 ( .C (clk), .D (signal_5665), .Q (signal_5666) ) ;
    buf_clk cell_3136 ( .C (clk), .D (signal_5681), .Q (signal_5682) ) ;
    buf_clk cell_3152 ( .C (clk), .D (signal_5697), .Q (signal_5698) ) ;
    buf_clk cell_3168 ( .C (clk), .D (signal_5713), .Q (signal_5714) ) ;
    buf_clk cell_3184 ( .C (clk), .D (signal_5729), .Q (signal_5730) ) ;
    buf_clk cell_3200 ( .C (clk), .D (signal_5745), .Q (signal_5746) ) ;
    buf_clk cell_3216 ( .C (clk), .D (signal_5761), .Q (signal_5762) ) ;
    buf_clk cell_3232 ( .C (clk), .D (signal_5777), .Q (signal_5778) ) ;
    buf_clk cell_3248 ( .C (clk), .D (signal_5793), .Q (signal_5794) ) ;
    buf_clk cell_3264 ( .C (clk), .D (signal_5809), .Q (signal_5810) ) ;
    buf_clk cell_3280 ( .C (clk), .D (signal_5825), .Q (signal_5826) ) ;
    buf_clk cell_3296 ( .C (clk), .D (signal_5841), .Q (signal_5842) ) ;
    buf_clk cell_3312 ( .C (clk), .D (signal_5857), .Q (signal_5858) ) ;
    buf_clk cell_3328 ( .C (clk), .D (signal_5873), .Q (signal_5874) ) ;
    buf_clk cell_3344 ( .C (clk), .D (signal_5889), .Q (signal_5890) ) ;
    buf_clk cell_3360 ( .C (clk), .D (signal_5905), .Q (signal_5906) ) ;
    buf_clk cell_3376 ( .C (clk), .D (signal_5921), .Q (signal_5922) ) ;
    buf_clk cell_3392 ( .C (clk), .D (signal_5937), .Q (signal_5938) ) ;
    buf_clk cell_3408 ( .C (clk), .D (signal_5953), .Q (signal_5954) ) ;
    buf_clk cell_3424 ( .C (clk), .D (signal_5969), .Q (signal_5970) ) ;
    buf_clk cell_3440 ( .C (clk), .D (signal_5985), .Q (signal_5986) ) ;
    buf_clk cell_3456 ( .C (clk), .D (signal_6001), .Q (signal_6002) ) ;
    buf_clk cell_3472 ( .C (clk), .D (signal_6017), .Q (signal_6018) ) ;
    buf_clk cell_3488 ( .C (clk), .D (signal_6033), .Q (signal_6034) ) ;
    buf_clk cell_3504 ( .C (clk), .D (signal_6049), .Q (signal_6050) ) ;
    buf_clk cell_3520 ( .C (clk), .D (signal_6065), .Q (signal_6066) ) ;
    buf_clk cell_3536 ( .C (clk), .D (signal_6081), .Q (signal_6082) ) ;
    buf_clk cell_3552 ( .C (clk), .D (signal_6097), .Q (signal_6098) ) ;
    buf_clk cell_3568 ( .C (clk), .D (signal_6113), .Q (signal_6114) ) ;
    buf_clk cell_3584 ( .C (clk), .D (signal_6129), .Q (signal_6130) ) ;
    buf_clk cell_3600 ( .C (clk), .D (signal_6145), .Q (signal_6146) ) ;
    buf_clk cell_3616 ( .C (clk), .D (signal_6161), .Q (signal_6162) ) ;
    buf_clk cell_3632 ( .C (clk), .D (signal_6177), .Q (signal_6178) ) ;
    buf_clk cell_3648 ( .C (clk), .D (signal_6193), .Q (signal_6194) ) ;
    buf_clk cell_3664 ( .C (clk), .D (signal_6209), .Q (signal_6210) ) ;
    buf_clk cell_3680 ( .C (clk), .D (signal_6225), .Q (signal_6226) ) ;
    buf_clk cell_3696 ( .C (clk), .D (signal_6241), .Q (signal_6242) ) ;
    buf_clk cell_3712 ( .C (clk), .D (signal_6257), .Q (signal_6258) ) ;
    buf_clk cell_3728 ( .C (clk), .D (signal_6273), .Q (signal_6274) ) ;
    buf_clk cell_3744 ( .C (clk), .D (signal_6289), .Q (signal_6290) ) ;
    buf_clk cell_3760 ( .C (clk), .D (signal_6305), .Q (signal_6306) ) ;
    buf_clk cell_3776 ( .C (clk), .D (signal_6321), .Q (signal_6322) ) ;
    buf_clk cell_3792 ( .C (clk), .D (signal_6337), .Q (signal_6338) ) ;
    buf_clk cell_3808 ( .C (clk), .D (signal_6353), .Q (signal_6354) ) ;
    buf_clk cell_3824 ( .C (clk), .D (signal_6369), .Q (signal_6370) ) ;
    buf_clk cell_3840 ( .C (clk), .D (signal_6385), .Q (signal_6386) ) ;
    buf_clk cell_3856 ( .C (clk), .D (signal_6401), .Q (signal_6402) ) ;
    buf_clk cell_3872 ( .C (clk), .D (signal_6417), .Q (signal_6418) ) ;
    buf_clk cell_3888 ( .C (clk), .D (signal_6433), .Q (signal_6434) ) ;
    buf_clk cell_3904 ( .C (clk), .D (signal_6449), .Q (signal_6450) ) ;
    buf_clk cell_3920 ( .C (clk), .D (signal_6465), .Q (signal_6466) ) ;
    buf_clk cell_3936 ( .C (clk), .D (signal_6481), .Q (signal_6482) ) ;
    buf_clk cell_3952 ( .C (clk), .D (signal_6497), .Q (signal_6498) ) ;
    buf_clk cell_3968 ( .C (clk), .D (signal_6513), .Q (signal_6514) ) ;
    buf_clk cell_3984 ( .C (clk), .D (signal_6529), .Q (signal_6530) ) ;
    buf_clk cell_4000 ( .C (clk), .D (signal_6545), .Q (signal_6546) ) ;
    buf_clk cell_4016 ( .C (clk), .D (signal_6561), .Q (signal_6562) ) ;
    buf_clk cell_4032 ( .C (clk), .D (signal_6577), .Q (signal_6578) ) ;
    buf_clk cell_4048 ( .C (clk), .D (signal_6593), .Q (signal_6594) ) ;
    buf_clk cell_4064 ( .C (clk), .D (signal_6609), .Q (signal_6610) ) ;
    buf_clk cell_4080 ( .C (clk), .D (signal_6625), .Q (signal_6626) ) ;
    buf_clk cell_4096 ( .C (clk), .D (signal_6641), .Q (signal_6642) ) ;
    buf_clk cell_4112 ( .C (clk), .D (signal_6657), .Q (signal_6658) ) ;
    buf_clk cell_4128 ( .C (clk), .D (signal_6673), .Q (signal_6674) ) ;
    buf_clk cell_4144 ( .C (clk), .D (signal_6689), .Q (signal_6690) ) ;
    buf_clk cell_4160 ( .C (clk), .D (signal_6705), .Q (signal_6706) ) ;
    buf_clk cell_4176 ( .C (clk), .D (signal_6721), .Q (signal_6722) ) ;
    buf_clk cell_4192 ( .C (clk), .D (signal_6737), .Q (signal_6738) ) ;
    buf_clk cell_4208 ( .C (clk), .D (signal_6753), .Q (signal_6754) ) ;
    buf_clk cell_4224 ( .C (clk), .D (signal_6769), .Q (signal_6770) ) ;
    buf_clk cell_4240 ( .C (clk), .D (signal_6785), .Q (signal_6786) ) ;
    buf_clk cell_4256 ( .C (clk), .D (signal_6801), .Q (signal_6802) ) ;
    buf_clk cell_4272 ( .C (clk), .D (signal_6817), .Q (signal_6818) ) ;
    buf_clk cell_4288 ( .C (clk), .D (signal_6833), .Q (signal_6834) ) ;
    buf_clk cell_4304 ( .C (clk), .D (signal_6849), .Q (signal_6850) ) ;
    buf_clk cell_4320 ( .C (clk), .D (signal_6865), .Q (signal_6866) ) ;
    buf_clk cell_4336 ( .C (clk), .D (signal_6881), .Q (signal_6882) ) ;
    buf_clk cell_4352 ( .C (clk), .D (signal_6897), .Q (signal_6898) ) ;
    buf_clk cell_4368 ( .C (clk), .D (signal_6913), .Q (signal_6914) ) ;
    buf_clk cell_4384 ( .C (clk), .D (signal_6929), .Q (signal_6930) ) ;
    buf_clk cell_4400 ( .C (clk), .D (signal_6945), .Q (signal_6946) ) ;
    buf_clk cell_4444 ( .C (clk), .D (signal_6989), .Q (signal_6990) ) ;
    buf_clk cell_4460 ( .C (clk), .D (signal_7005), .Q (signal_7006) ) ;
    buf_clk cell_4476 ( .C (clk), .D (signal_7021), .Q (signal_7022) ) ;
    buf_clk cell_4492 ( .C (clk), .D (signal_7037), .Q (signal_7038) ) ;
    buf_clk cell_4508 ( .C (clk), .D (signal_7053), .Q (signal_7054) ) ;
    buf_clk cell_4524 ( .C (clk), .D (signal_7069), .Q (signal_7070) ) ;
    buf_clk cell_4540 ( .C (clk), .D (signal_7085), .Q (signal_7086) ) ;
    buf_clk cell_4556 ( .C (clk), .D (signal_7101), .Q (signal_7102) ) ;
    buf_clk cell_4572 ( .C (clk), .D (signal_7117), .Q (signal_7118) ) ;
    buf_clk cell_4588 ( .C (clk), .D (signal_7133), .Q (signal_7134) ) ;
    buf_clk cell_4604 ( .C (clk), .D (signal_7149), .Q (signal_7150) ) ;
    buf_clk cell_4620 ( .C (clk), .D (signal_7165), .Q (signal_7166) ) ;
    buf_clk cell_4636 ( .C (clk), .D (signal_7181), .Q (signal_7182) ) ;
    buf_clk cell_4652 ( .C (clk), .D (signal_7197), .Q (signal_7198) ) ;
    buf_clk cell_4668 ( .C (clk), .D (signal_7213), .Q (signal_7214) ) ;
    buf_clk cell_4684 ( .C (clk), .D (signal_7229), .Q (signal_7230) ) ;
    buf_clk cell_4700 ( .C (clk), .D (signal_7245), .Q (signal_7246) ) ;
    buf_clk cell_4716 ( .C (clk), .D (signal_7261), .Q (signal_7262) ) ;
    buf_clk cell_4732 ( .C (clk), .D (signal_7277), .Q (signal_7278) ) ;
    buf_clk cell_4748 ( .C (clk), .D (signal_7293), .Q (signal_7294) ) ;
    buf_clk cell_4764 ( .C (clk), .D (signal_7309), .Q (signal_7310) ) ;
    buf_clk cell_4780 ( .C (clk), .D (signal_7325), .Q (signal_7326) ) ;
    buf_clk cell_4796 ( .C (clk), .D (signal_7341), .Q (signal_7342) ) ;
    buf_clk cell_4812 ( .C (clk), .D (signal_7357), .Q (signal_7358) ) ;
    buf_clk cell_4828 ( .C (clk), .D (signal_7373), .Q (signal_7374) ) ;
    buf_clk cell_4844 ( .C (clk), .D (signal_7389), .Q (signal_7390) ) ;
    buf_clk cell_4860 ( .C (clk), .D (signal_7405), .Q (signal_7406) ) ;
    buf_clk cell_4876 ( .C (clk), .D (signal_7421), .Q (signal_7422) ) ;
    buf_clk cell_4892 ( .C (clk), .D (signal_7437), .Q (signal_7438) ) ;
    buf_clk cell_4908 ( .C (clk), .D (signal_7453), .Q (signal_7454) ) ;
    buf_clk cell_4924 ( .C (clk), .D (signal_7469), .Q (signal_7470) ) ;
    buf_clk cell_4940 ( .C (clk), .D (signal_7485), .Q (signal_7486) ) ;
    buf_clk cell_4956 ( .C (clk), .D (signal_7501), .Q (signal_7502) ) ;
    buf_clk cell_4972 ( .C (clk), .D (signal_7517), .Q (signal_7518) ) ;
    buf_clk cell_4988 ( .C (clk), .D (signal_7533), .Q (signal_7534) ) ;
    buf_clk cell_5004 ( .C (clk), .D (signal_7549), .Q (signal_7550) ) ;
    buf_clk cell_5020 ( .C (clk), .D (signal_7565), .Q (signal_7566) ) ;
    buf_clk cell_5036 ( .C (clk), .D (signal_7581), .Q (signal_7582) ) ;
    buf_clk cell_5052 ( .C (clk), .D (signal_7597), .Q (signal_7598) ) ;
    buf_clk cell_5068 ( .C (clk), .D (signal_7613), .Q (signal_7614) ) ;
    buf_clk cell_5084 ( .C (clk), .D (signal_7629), .Q (signal_7630) ) ;
    buf_clk cell_5100 ( .C (clk), .D (signal_7645), .Q (signal_7646) ) ;
    buf_clk cell_5116 ( .C (clk), .D (signal_7661), .Q (signal_7662) ) ;
    buf_clk cell_5132 ( .C (clk), .D (signal_7677), .Q (signal_7678) ) ;
    buf_clk cell_5148 ( .C (clk), .D (signal_7693), .Q (signal_7694) ) ;
    buf_clk cell_5164 ( .C (clk), .D (signal_7709), .Q (signal_7710) ) ;
    buf_clk cell_5180 ( .C (clk), .D (signal_7725), .Q (signal_7726) ) ;
    buf_clk cell_5196 ( .C (clk), .D (signal_7741), .Q (signal_7742) ) ;
    buf_clk cell_5212 ( .C (clk), .D (signal_7757), .Q (signal_7758) ) ;
    buf_clk cell_5228 ( .C (clk), .D (signal_7773), .Q (signal_7774) ) ;
    buf_clk cell_5244 ( .C (clk), .D (signal_7789), .Q (signal_7790) ) ;
    buf_clk cell_5260 ( .C (clk), .D (signal_7805), .Q (signal_7806) ) ;
    buf_clk cell_5276 ( .C (clk), .D (signal_7821), .Q (signal_7822) ) ;
    buf_clk cell_5292 ( .C (clk), .D (signal_7837), .Q (signal_7838) ) ;
    buf_clk cell_5308 ( .C (clk), .D (signal_7853), .Q (signal_7854) ) ;
    buf_clk cell_5324 ( .C (clk), .D (signal_7869), .Q (signal_7870) ) ;
    buf_clk cell_5340 ( .C (clk), .D (signal_7885), .Q (signal_7886) ) ;
    buf_clk cell_5356 ( .C (clk), .D (signal_7901), .Q (signal_7902) ) ;
    buf_clk cell_5372 ( .C (clk), .D (signal_7917), .Q (signal_7918) ) ;
    buf_clk cell_5388 ( .C (clk), .D (signal_7933), .Q (signal_7934) ) ;
    buf_clk cell_5404 ( .C (clk), .D (signal_7949), .Q (signal_7950) ) ;
    buf_clk cell_5420 ( .C (clk), .D (signal_7965), .Q (signal_7966) ) ;
    buf_clk cell_5436 ( .C (clk), .D (signal_7981), .Q (signal_7982) ) ;
    buf_clk cell_5452 ( .C (clk), .D (signal_7997), .Q (signal_7998) ) ;
    buf_clk cell_5468 ( .C (clk), .D (signal_8013), .Q (signal_8014) ) ;
    buf_clk cell_5484 ( .C (clk), .D (signal_8029), .Q (signal_8030) ) ;
    buf_clk cell_5500 ( .C (clk), .D (signal_8045), .Q (signal_8046) ) ;
    buf_clk cell_5516 ( .C (clk), .D (signal_8061), .Q (signal_8062) ) ;
    buf_clk cell_5532 ( .C (clk), .D (signal_8077), .Q (signal_8078) ) ;
    buf_clk cell_5548 ( .C (clk), .D (signal_8093), .Q (signal_8094) ) ;
    buf_clk cell_5564 ( .C (clk), .D (signal_8109), .Q (signal_8110) ) ;
    buf_clk cell_5580 ( .C (clk), .D (signal_8125), .Q (signal_8126) ) ;
    buf_clk cell_5596 ( .C (clk), .D (signal_8141), .Q (signal_8142) ) ;
    buf_clk cell_5612 ( .C (clk), .D (signal_8157), .Q (signal_8158) ) ;
    buf_clk cell_5628 ( .C (clk), .D (signal_8173), .Q (signal_8174) ) ;
    buf_clk cell_5644 ( .C (clk), .D (signal_8189), .Q (signal_8190) ) ;
    buf_clk cell_5660 ( .C (clk), .D (signal_8205), .Q (signal_8206) ) ;
    buf_clk cell_5676 ( .C (clk), .D (signal_8221), .Q (signal_8222) ) ;
    buf_clk cell_5692 ( .C (clk), .D (signal_8237), .Q (signal_8238) ) ;
    buf_clk cell_5708 ( .C (clk), .D (signal_8253), .Q (signal_8254) ) ;
    buf_clk cell_5724 ( .C (clk), .D (signal_8269), .Q (signal_8270) ) ;
    buf_clk cell_5740 ( .C (clk), .D (signal_8285), .Q (signal_8286) ) ;
    buf_clk cell_5756 ( .C (clk), .D (signal_8301), .Q (signal_8302) ) ;
    buf_clk cell_5772 ( .C (clk), .D (signal_8317), .Q (signal_8318) ) ;
    buf_clk cell_5788 ( .C (clk), .D (signal_8333), .Q (signal_8334) ) ;
    buf_clk cell_5804 ( .C (clk), .D (signal_8349), .Q (signal_8350) ) ;
    buf_clk cell_5820 ( .C (clk), .D (signal_8365), .Q (signal_8366) ) ;
    buf_clk cell_5836 ( .C (clk), .D (signal_8381), .Q (signal_8382) ) ;
    buf_clk cell_5852 ( .C (clk), .D (signal_8397), .Q (signal_8398) ) ;
    buf_clk cell_5868 ( .C (clk), .D (signal_8413), .Q (signal_8414) ) ;
    buf_clk cell_5884 ( .C (clk), .D (signal_8429), .Q (signal_8430) ) ;
    buf_clk cell_5900 ( .C (clk), .D (signal_8445), .Q (signal_8446) ) ;
    buf_clk cell_5916 ( .C (clk), .D (signal_8461), .Q (signal_8462) ) ;
    buf_clk cell_5932 ( .C (clk), .D (signal_8477), .Q (signal_8478) ) ;
    buf_clk cell_5948 ( .C (clk), .D (signal_8493), .Q (signal_8494) ) ;
    buf_clk cell_5964 ( .C (clk), .D (signal_8509), .Q (signal_8510) ) ;
    buf_clk cell_5980 ( .C (clk), .D (signal_8525), .Q (signal_8526) ) ;
    buf_clk cell_5996 ( .C (clk), .D (signal_8541), .Q (signal_8542) ) ;
    buf_clk cell_6012 ( .C (clk), .D (signal_8557), .Q (signal_8558) ) ;
    buf_clk cell_6028 ( .C (clk), .D (signal_8573), .Q (signal_8574) ) ;
    buf_clk cell_6044 ( .C (clk), .D (signal_8589), .Q (signal_8590) ) ;
    buf_clk cell_6060 ( .C (clk), .D (signal_8605), .Q (signal_8606) ) ;
    buf_clk cell_6076 ( .C (clk), .D (signal_8621), .Q (signal_8622) ) ;
    buf_clk cell_6092 ( .C (clk), .D (signal_8637), .Q (signal_8638) ) ;
    buf_clk cell_6108 ( .C (clk), .D (signal_8653), .Q (signal_8654) ) ;
    buf_clk cell_6124 ( .C (clk), .D (signal_8669), .Q (signal_8670) ) ;
    buf_clk cell_6140 ( .C (clk), .D (signal_8685), .Q (signal_8686) ) ;
    buf_clk cell_6156 ( .C (clk), .D (signal_8701), .Q (signal_8702) ) ;
    buf_clk cell_6172 ( .C (clk), .D (signal_8717), .Q (signal_8718) ) ;
    buf_clk cell_6188 ( .C (clk), .D (signal_8733), .Q (signal_8734) ) ;
    buf_clk cell_6204 ( .C (clk), .D (signal_8749), .Q (signal_8750) ) ;
    buf_clk cell_6220 ( .C (clk), .D (signal_8765), .Q (signal_8766) ) ;
    buf_clk cell_6236 ( .C (clk), .D (signal_8781), .Q (signal_8782) ) ;
    buf_clk cell_6252 ( .C (clk), .D (signal_8797), .Q (signal_8798) ) ;
    buf_clk cell_6268 ( .C (clk), .D (signal_8813), .Q (signal_8814) ) ;
    buf_clk cell_6284 ( .C (clk), .D (signal_8829), .Q (signal_8830) ) ;
    buf_clk cell_6300 ( .C (clk), .D (signal_8845), .Q (signal_8846) ) ;
    buf_clk cell_6316 ( .C (clk), .D (signal_8861), .Q (signal_8862) ) ;
    buf_clk cell_6332 ( .C (clk), .D (signal_8877), .Q (signal_8878) ) ;
    buf_clk cell_6348 ( .C (clk), .D (signal_8893), .Q (signal_8894) ) ;
    buf_clk cell_6364 ( .C (clk), .D (signal_8909), .Q (signal_8910) ) ;
    buf_clk cell_6380 ( .C (clk), .D (signal_8925), .Q (signal_8926) ) ;
    buf_clk cell_6396 ( .C (clk), .D (signal_8941), .Q (signal_8942) ) ;
    buf_clk cell_6412 ( .C (clk), .D (signal_8957), .Q (signal_8958) ) ;
    buf_clk cell_6428 ( .C (clk), .D (signal_8973), .Q (signal_8974) ) ;
    buf_clk cell_6444 ( .C (clk), .D (signal_8989), .Q (signal_8990) ) ;
    buf_clk cell_6460 ( .C (clk), .D (signal_9005), .Q (signal_9006) ) ;
    buf_clk cell_6476 ( .C (clk), .D (signal_9021), .Q (signal_9022) ) ;
    buf_clk cell_6492 ( .C (clk), .D (signal_9037), .Q (signal_9038) ) ;
    buf_clk cell_6508 ( .C (clk), .D (signal_9053), .Q (signal_9054) ) ;
    buf_clk cell_6524 ( .C (clk), .D (signal_9069), .Q (signal_9070) ) ;
    buf_clk cell_6540 ( .C (clk), .D (signal_9085), .Q (signal_9086) ) ;
    buf_clk cell_6556 ( .C (clk), .D (signal_9101), .Q (signal_9102) ) ;
    buf_clk cell_6572 ( .C (clk), .D (signal_9117), .Q (signal_9118) ) ;
    buf_clk cell_6588 ( .C (clk), .D (signal_9133), .Q (signal_9134) ) ;
    buf_clk cell_6604 ( .C (clk), .D (signal_9149), .Q (signal_9150) ) ;
    buf_clk cell_6620 ( .C (clk), .D (signal_9165), .Q (signal_9166) ) ;
    buf_clk cell_6636 ( .C (clk), .D (signal_9181), .Q (signal_9182) ) ;
    buf_clk cell_6652 ( .C (clk), .D (signal_9197), .Q (signal_9198) ) ;
    buf_clk cell_6668 ( .C (clk), .D (signal_9213), .Q (signal_9214) ) ;
    buf_clk cell_6684 ( .C (clk), .D (signal_9229), .Q (signal_9230) ) ;
    buf_clk cell_6700 ( .C (clk), .D (signal_9245), .Q (signal_9246) ) ;
    buf_clk cell_6716 ( .C (clk), .D (signal_9261), .Q (signal_9262) ) ;
    buf_clk cell_6732 ( .C (clk), .D (signal_9277), .Q (signal_9278) ) ;
    buf_clk cell_6748 ( .C (clk), .D (signal_9293), .Q (signal_9294) ) ;
    buf_clk cell_6764 ( .C (clk), .D (signal_9309), .Q (signal_9310) ) ;
    buf_clk cell_6780 ( .C (clk), .D (signal_9325), .Q (signal_9326) ) ;
    buf_clk cell_6796 ( .C (clk), .D (signal_9341), .Q (signal_9342) ) ;
    buf_clk cell_6812 ( .C (clk), .D (signal_9357), .Q (signal_9358) ) ;
    buf_clk cell_6828 ( .C (clk), .D (signal_9373), .Q (signal_9374) ) ;
    buf_clk cell_6844 ( .C (clk), .D (signal_9389), .Q (signal_9390) ) ;
    buf_clk cell_6860 ( .C (clk), .D (signal_9405), .Q (signal_9406) ) ;
    buf_clk cell_6876 ( .C (clk), .D (signal_9421), .Q (signal_9422) ) ;
    buf_clk cell_6892 ( .C (clk), .D (signal_9437), .Q (signal_9438) ) ;
    buf_clk cell_6908 ( .C (clk), .D (signal_9453), .Q (signal_9454) ) ;
    buf_clk cell_6924 ( .C (clk), .D (signal_9469), .Q (signal_9470) ) ;
    buf_clk cell_6940 ( .C (clk), .D (signal_9485), .Q (signal_9486) ) ;
    buf_clk cell_6956 ( .C (clk), .D (signal_9501), .Q (signal_9502) ) ;
    buf_clk cell_6972 ( .C (clk), .D (signal_9517), .Q (signal_9518) ) ;
    buf_clk cell_6988 ( .C (clk), .D (signal_9533), .Q (signal_9534) ) ;
    buf_clk cell_7004 ( .C (clk), .D (signal_9549), .Q (signal_9550) ) ;
    buf_clk cell_7020 ( .C (clk), .D (signal_9565), .Q (signal_9566) ) ;
    buf_clk cell_7036 ( .C (clk), .D (signal_9581), .Q (signal_9582) ) ;
    buf_clk cell_7052 ( .C (clk), .D (signal_9597), .Q (signal_9598) ) ;
    buf_clk cell_7068 ( .C (clk), .D (signal_9613), .Q (signal_9614) ) ;
    buf_clk cell_7084 ( .C (clk), .D (signal_9629), .Q (signal_9630) ) ;
    buf_clk cell_7100 ( .C (clk), .D (signal_9645), .Q (signal_9646) ) ;
    buf_clk cell_7116 ( .C (clk), .D (signal_9661), .Q (signal_9662) ) ;
    buf_clk cell_7132 ( .C (clk), .D (signal_9677), .Q (signal_9678) ) ;
    buf_clk cell_7148 ( .C (clk), .D (signal_9693), .Q (signal_9694) ) ;
    buf_clk cell_7164 ( .C (clk), .D (signal_9709), .Q (signal_9710) ) ;
    buf_clk cell_7180 ( .C (clk), .D (signal_9725), .Q (signal_9726) ) ;
    buf_clk cell_7196 ( .C (clk), .D (signal_9741), .Q (signal_9742) ) ;
    buf_clk cell_7212 ( .C (clk), .D (signal_9757), .Q (signal_9758) ) ;
    buf_clk cell_7228 ( .C (clk), .D (signal_9773), .Q (signal_9774) ) ;
    buf_clk cell_7244 ( .C (clk), .D (signal_9789), .Q (signal_9790) ) ;
    buf_clk cell_7260 ( .C (clk), .D (signal_9805), .Q (signal_9806) ) ;
    buf_clk cell_7276 ( .C (clk), .D (signal_9821), .Q (signal_9822) ) ;
    buf_clk cell_7292 ( .C (clk), .D (signal_9837), .Q (signal_9838) ) ;
    buf_clk cell_7308 ( .C (clk), .D (signal_9853), .Q (signal_9854) ) ;
    buf_clk cell_7324 ( .C (clk), .D (signal_9869), .Q (signal_9870) ) ;
    buf_clk cell_7340 ( .C (clk), .D (signal_9885), .Q (signal_9886) ) ;
    buf_clk cell_7356 ( .C (clk), .D (signal_9901), .Q (signal_9902) ) ;
    buf_clk cell_7372 ( .C (clk), .D (signal_9917), .Q (signal_9918) ) ;
    buf_clk cell_7388 ( .C (clk), .D (signal_9933), .Q (signal_9934) ) ;
    buf_clk cell_7404 ( .C (clk), .D (signal_9949), .Q (signal_9950) ) ;
    buf_clk cell_7420 ( .C (clk), .D (signal_9965), .Q (signal_9966) ) ;
    buf_clk cell_7436 ( .C (clk), .D (signal_9981), .Q (signal_9982) ) ;
    buf_clk cell_7452 ( .C (clk), .D (signal_9997), .Q (signal_9998) ) ;
    buf_clk cell_7468 ( .C (clk), .D (signal_10013), .Q (signal_10014) ) ;
    buf_clk cell_7484 ( .C (clk), .D (signal_10029), .Q (signal_10030) ) ;
    buf_clk cell_7500 ( .C (clk), .D (signal_10045), .Q (signal_10046) ) ;
    buf_clk cell_7516 ( .C (clk), .D (signal_10061), .Q (signal_10062) ) ;
    buf_clk cell_7532 ( .C (clk), .D (signal_10077), .Q (signal_10078) ) ;
    buf_clk cell_7548 ( .C (clk), .D (signal_10093), .Q (signal_10094) ) ;
    buf_clk cell_7564 ( .C (clk), .D (signal_10109), .Q (signal_10110) ) ;
    buf_clk cell_7580 ( .C (clk), .D (signal_10125), .Q (signal_10126) ) ;
    buf_clk cell_7596 ( .C (clk), .D (signal_10141), .Q (signal_10142) ) ;
    buf_clk cell_7612 ( .C (clk), .D (signal_10157), .Q (signal_10158) ) ;
    buf_clk cell_7628 ( .C (clk), .D (signal_10173), .Q (signal_10174) ) ;
    buf_clk cell_7644 ( .C (clk), .D (signal_10189), .Q (signal_10190) ) ;
    buf_clk cell_7660 ( .C (clk), .D (signal_10205), .Q (signal_10206) ) ;
    buf_clk cell_7676 ( .C (clk), .D (signal_10221), .Q (signal_10222) ) ;
    buf_clk cell_7692 ( .C (clk), .D (signal_10237), .Q (signal_10238) ) ;
    buf_clk cell_7708 ( .C (clk), .D (signal_10253), .Q (signal_10254) ) ;
    buf_clk cell_7724 ( .C (clk), .D (signal_10269), .Q (signal_10270) ) ;
    buf_clk cell_7740 ( .C (clk), .D (signal_10285), .Q (signal_10286) ) ;
    buf_clk cell_7756 ( .C (clk), .D (signal_10301), .Q (signal_10302) ) ;
    buf_clk cell_7772 ( .C (clk), .D (signal_10317), .Q (signal_10318) ) ;
    buf_clk cell_7788 ( .C (clk), .D (signal_10333), .Q (signal_10334) ) ;
    buf_clk cell_7804 ( .C (clk), .D (signal_10349), .Q (signal_10350) ) ;
    buf_clk cell_7820 ( .C (clk), .D (signal_10365), .Q (signal_10366) ) ;
    buf_clk cell_7836 ( .C (clk), .D (signal_10381), .Q (signal_10382) ) ;
    buf_clk cell_7852 ( .C (clk), .D (signal_10397), .Q (signal_10398) ) ;
    buf_clk cell_7868 ( .C (clk), .D (signal_10413), .Q (signal_10414) ) ;
    buf_clk cell_7884 ( .C (clk), .D (signal_10429), .Q (signal_10430) ) ;
    buf_clk cell_7900 ( .C (clk), .D (signal_10445), .Q (signal_10446) ) ;
    buf_clk cell_7916 ( .C (clk), .D (signal_10461), .Q (signal_10462) ) ;
    buf_clk cell_7932 ( .C (clk), .D (signal_10477), .Q (signal_10478) ) ;
    buf_clk cell_7948 ( .C (clk), .D (signal_10493), .Q (signal_10494) ) ;
    buf_clk cell_7964 ( .C (clk), .D (signal_10509), .Q (signal_10510) ) ;
    buf_clk cell_7980 ( .C (clk), .D (signal_10525), .Q (signal_10526) ) ;
    buf_clk cell_7996 ( .C (clk), .D (signal_10541), .Q (signal_10542) ) ;
    buf_clk cell_8012 ( .C (clk), .D (signal_10557), .Q (signal_10558) ) ;
    buf_clk cell_8028 ( .C (clk), .D (signal_10573), .Q (signal_10574) ) ;
    buf_clk cell_8044 ( .C (clk), .D (signal_10589), .Q (signal_10590) ) ;
    buf_clk cell_8060 ( .C (clk), .D (signal_10605), .Q (signal_10606) ) ;
    buf_clk cell_8076 ( .C (clk), .D (signal_10621), .Q (signal_10622) ) ;
    buf_clk cell_8092 ( .C (clk), .D (signal_10637), .Q (signal_10638) ) ;
    buf_clk cell_8108 ( .C (clk), .D (signal_10653), .Q (signal_10654) ) ;
    buf_clk cell_8124 ( .C (clk), .D (signal_10669), .Q (signal_10670) ) ;
    buf_clk cell_8140 ( .C (clk), .D (signal_10685), .Q (signal_10686) ) ;
    buf_clk cell_8156 ( .C (clk), .D (signal_10701), .Q (signal_10702) ) ;
    buf_clk cell_8172 ( .C (clk), .D (signal_10717), .Q (signal_10718) ) ;
    buf_clk cell_8188 ( .C (clk), .D (signal_10733), .Q (signal_10734) ) ;
    buf_clk cell_8204 ( .C (clk), .D (signal_10749), .Q (signal_10750) ) ;
    buf_clk cell_8220 ( .C (clk), .D (signal_10765), .Q (signal_10766) ) ;
    buf_clk cell_8236 ( .C (clk), .D (signal_10781), .Q (signal_10782) ) ;
    buf_clk cell_8252 ( .C (clk), .D (signal_10797), .Q (signal_10798) ) ;
    buf_clk cell_8268 ( .C (clk), .D (signal_10813), .Q (signal_10814) ) ;
    buf_clk cell_8284 ( .C (clk), .D (signal_10829), .Q (signal_10830) ) ;
    buf_clk cell_8300 ( .C (clk), .D (signal_10845), .Q (signal_10846) ) ;
    buf_clk cell_8316 ( .C (clk), .D (signal_10861), .Q (signal_10862) ) ;
    buf_clk cell_8332 ( .C (clk), .D (signal_10877), .Q (signal_10878) ) ;
    buf_clk cell_8348 ( .C (clk), .D (signal_10893), .Q (signal_10894) ) ;
    buf_clk cell_8364 ( .C (clk), .D (signal_10909), .Q (signal_10910) ) ;
    buf_clk cell_8380 ( .C (clk), .D (signal_10925), .Q (signal_10926) ) ;
    buf_clk cell_8396 ( .C (clk), .D (signal_10941), .Q (signal_10942) ) ;
    buf_clk cell_8412 ( .C (clk), .D (signal_10957), .Q (signal_10958) ) ;
    buf_clk cell_8428 ( .C (clk), .D (signal_10973), .Q (signal_10974) ) ;
    buf_clk cell_8444 ( .C (clk), .D (signal_10989), .Q (signal_10990) ) ;
    buf_clk cell_8460 ( .C (clk), .D (signal_11005), .Q (signal_11006) ) ;
    buf_clk cell_8476 ( .C (clk), .D (signal_11021), .Q (signal_11022) ) ;
    buf_clk cell_8492 ( .C (clk), .D (signal_11037), .Q (signal_11038) ) ;
    buf_clk cell_8508 ( .C (clk), .D (signal_11053), .Q (signal_11054) ) ;
    buf_clk cell_8524 ( .C (clk), .D (signal_11069), .Q (signal_11070) ) ;
    buf_clk cell_8540 ( .C (clk), .D (signal_11085), .Q (signal_11086) ) ;
    buf_clk cell_8556 ( .C (clk), .D (signal_11101), .Q (signal_11102) ) ;
    buf_clk cell_8572 ( .C (clk), .D (signal_11117), .Q (signal_11118) ) ;
    buf_clk cell_8588 ( .C (clk), .D (signal_11133), .Q (signal_11134) ) ;
    buf_clk cell_8604 ( .C (clk), .D (signal_11149), .Q (signal_11150) ) ;
    buf_clk cell_8620 ( .C (clk), .D (signal_11165), .Q (signal_11166) ) ;
    buf_clk cell_8636 ( .C (clk), .D (signal_11181), .Q (signal_11182) ) ;
    buf_clk cell_8652 ( .C (clk), .D (signal_11197), .Q (signal_11198) ) ;
    buf_clk cell_8668 ( .C (clk), .D (signal_11213), .Q (signal_11214) ) ;
    buf_clk cell_8684 ( .C (clk), .D (signal_11229), .Q (signal_11230) ) ;
    buf_clk cell_8700 ( .C (clk), .D (signal_11245), .Q (signal_11246) ) ;
    buf_clk cell_8716 ( .C (clk), .D (signal_11261), .Q (signal_11262) ) ;
    buf_clk cell_8732 ( .C (clk), .D (signal_11277), .Q (signal_11278) ) ;
    buf_clk cell_8748 ( .C (clk), .D (signal_11293), .Q (signal_11294) ) ;
    buf_clk cell_8764 ( .C (clk), .D (signal_11309), .Q (signal_11310) ) ;
    buf_clk cell_8780 ( .C (clk), .D (signal_11325), .Q (signal_11326) ) ;
    buf_clk cell_8796 ( .C (clk), .D (signal_11341), .Q (signal_11342) ) ;
    buf_clk cell_8812 ( .C (clk), .D (signal_11357), .Q (signal_11358) ) ;
    buf_clk cell_8828 ( .C (clk), .D (signal_11373), .Q (signal_11374) ) ;
    buf_clk cell_8844 ( .C (clk), .D (signal_11389), .Q (signal_11390) ) ;
    buf_clk cell_8860 ( .C (clk), .D (signal_11405), .Q (signal_11406) ) ;
    buf_clk cell_8876 ( .C (clk), .D (signal_11421), .Q (signal_11422) ) ;
    buf_clk cell_8892 ( .C (clk), .D (signal_11437), .Q (signal_11438) ) ;
    buf_clk cell_8908 ( .C (clk), .D (signal_11453), .Q (signal_11454) ) ;
    buf_clk cell_8924 ( .C (clk), .D (signal_11469), .Q (signal_11470) ) ;
    buf_clk cell_8940 ( .C (clk), .D (signal_11485), .Q (signal_11486) ) ;
    buf_clk cell_8956 ( .C (clk), .D (signal_11501), .Q (signal_11502) ) ;
    buf_clk cell_8972 ( .C (clk), .D (signal_11517), .Q (signal_11518) ) ;
    buf_clk cell_8988 ( .C (clk), .D (signal_11533), .Q (signal_11534) ) ;
    buf_clk cell_9004 ( .C (clk), .D (signal_11549), .Q (signal_11550) ) ;
    buf_clk cell_9020 ( .C (clk), .D (signal_11565), .Q (signal_11566) ) ;
    buf_clk cell_9036 ( .C (clk), .D (signal_11581), .Q (signal_11582) ) ;
    buf_clk cell_9052 ( .C (clk), .D (signal_11597), .Q (signal_11598) ) ;
    buf_clk cell_9068 ( .C (clk), .D (signal_11613), .Q (signal_11614) ) ;
    buf_clk cell_9084 ( .C (clk), .D (signal_11629), .Q (signal_11630) ) ;
    buf_clk cell_9100 ( .C (clk), .D (signal_11645), .Q (signal_11646) ) ;
    buf_clk cell_9116 ( .C (clk), .D (signal_11661), .Q (signal_11662) ) ;
    buf_clk cell_9132 ( .C (clk), .D (signal_11677), .Q (signal_11678) ) ;
    buf_clk cell_9148 ( .C (clk), .D (signal_11693), .Q (signal_11694) ) ;
    buf_clk cell_9164 ( .C (clk), .D (signal_11709), .Q (signal_11710) ) ;
    buf_clk cell_9180 ( .C (clk), .D (signal_11725), .Q (signal_11726) ) ;
    buf_clk cell_9196 ( .C (clk), .D (signal_11741), .Q (signal_11742) ) ;
    buf_clk cell_9212 ( .C (clk), .D (signal_11757), .Q (signal_11758) ) ;
    buf_clk cell_9228 ( .C (clk), .D (signal_11773), .Q (signal_11774) ) ;
    buf_clk cell_9244 ( .C (clk), .D (signal_11789), .Q (signal_11790) ) ;
    buf_clk cell_9260 ( .C (clk), .D (signal_11805), .Q (signal_11806) ) ;
    buf_clk cell_9276 ( .C (clk), .D (signal_11821), .Q (signal_11822) ) ;
    buf_clk cell_9292 ( .C (clk), .D (signal_11837), .Q (signal_11838) ) ;
    buf_clk cell_9308 ( .C (clk), .D (signal_11853), .Q (signal_11854) ) ;
    buf_clk cell_9324 ( .C (clk), .D (signal_11869), .Q (signal_11870) ) ;
    buf_clk cell_9340 ( .C (clk), .D (signal_11885), .Q (signal_11886) ) ;
    buf_clk cell_9356 ( .C (clk), .D (signal_11901), .Q (signal_11902) ) ;
    buf_clk cell_9372 ( .C (clk), .D (signal_11917), .Q (signal_11918) ) ;
    buf_clk cell_9388 ( .C (clk), .D (signal_11933), .Q (signal_11934) ) ;
    buf_clk cell_9404 ( .C (clk), .D (signal_11949), .Q (signal_11950) ) ;
    buf_clk cell_9420 ( .C (clk), .D (signal_11965), .Q (signal_11966) ) ;
    buf_clk cell_9436 ( .C (clk), .D (signal_11981), .Q (signal_11982) ) ;
    buf_clk cell_9452 ( .C (clk), .D (signal_11997), .Q (signal_11998) ) ;
    buf_clk cell_9468 ( .C (clk), .D (signal_12013), .Q (signal_12014) ) ;
    buf_clk cell_9484 ( .C (clk), .D (signal_12029), .Q (signal_12030) ) ;
    buf_clk cell_9500 ( .C (clk), .D (signal_12045), .Q (signal_12046) ) ;
    buf_clk cell_9516 ( .C (clk), .D (signal_12061), .Q (signal_12062) ) ;
    buf_clk cell_9532 ( .C (clk), .D (signal_12077), .Q (signal_12078) ) ;
    buf_clk cell_9548 ( .C (clk), .D (signal_12093), .Q (signal_12094) ) ;
    buf_clk cell_9564 ( .C (clk), .D (signal_12109), .Q (signal_12110) ) ;
    buf_clk cell_9580 ( .C (clk), .D (signal_12125), .Q (signal_12126) ) ;
    buf_clk cell_9596 ( .C (clk), .D (signal_12141), .Q (signal_12142) ) ;
    buf_clk cell_9612 ( .C (clk), .D (signal_12157), .Q (signal_12158) ) ;
    buf_clk cell_9628 ( .C (clk), .D (signal_12173), .Q (signal_12174) ) ;
    buf_clk cell_9644 ( .C (clk), .D (signal_12189), .Q (signal_12190) ) ;
    buf_clk cell_9660 ( .C (clk), .D (signal_12205), .Q (signal_12206) ) ;
    buf_clk cell_9676 ( .C (clk), .D (signal_12221), .Q (signal_12222) ) ;
    buf_clk cell_9692 ( .C (clk), .D (signal_12237), .Q (signal_12238) ) ;
    buf_clk cell_9708 ( .C (clk), .D (signal_12253), .Q (signal_12254) ) ;
    buf_clk cell_9724 ( .C (clk), .D (signal_12269), .Q (signal_12270) ) ;
    buf_clk cell_9740 ( .C (clk), .D (signal_12285), .Q (signal_12286) ) ;
    buf_clk cell_9756 ( .C (clk), .D (signal_12301), .Q (signal_12302) ) ;
    buf_clk cell_9772 ( .C (clk), .D (signal_12317), .Q (signal_12318) ) ;
    buf_clk cell_9788 ( .C (clk), .D (signal_12333), .Q (signal_12334) ) ;
    buf_clk cell_9804 ( .C (clk), .D (signal_12349), .Q (signal_12350) ) ;
    buf_clk cell_9820 ( .C (clk), .D (signal_12365), .Q (signal_12366) ) ;
    buf_clk cell_9836 ( .C (clk), .D (signal_12381), .Q (signal_12382) ) ;
    buf_clk cell_9852 ( .C (clk), .D (signal_12397), .Q (signal_12398) ) ;
    buf_clk cell_9868 ( .C (clk), .D (signal_12413), .Q (signal_12414) ) ;
    buf_clk cell_9884 ( .C (clk), .D (signal_12429), .Q (signal_12430) ) ;
    buf_clk cell_9900 ( .C (clk), .D (signal_12445), .Q (signal_12446) ) ;
    buf_clk cell_9916 ( .C (clk), .D (signal_12461), .Q (signal_12462) ) ;
    buf_clk cell_9932 ( .C (clk), .D (signal_12477), .Q (signal_12478) ) ;
    buf_clk cell_9948 ( .C (clk), .D (signal_12493), .Q (signal_12494) ) ;
    buf_clk cell_9964 ( .C (clk), .D (signal_12509), .Q (signal_12510) ) ;
    buf_clk cell_9980 ( .C (clk), .D (signal_12525), .Q (signal_12526) ) ;
    buf_clk cell_9996 ( .C (clk), .D (signal_12541), .Q (signal_12542) ) ;
    buf_clk cell_10012 ( .C (clk), .D (signal_12557), .Q (signal_12558) ) ;
    buf_clk cell_10028 ( .C (clk), .D (signal_12573), .Q (signal_12574) ) ;
    buf_clk cell_10044 ( .C (clk), .D (signal_12589), .Q (signal_12590) ) ;
    buf_clk cell_10060 ( .C (clk), .D (signal_12605), .Q (signal_12606) ) ;
    buf_clk cell_10076 ( .C (clk), .D (signal_12621), .Q (signal_12622) ) ;
    buf_clk cell_10092 ( .C (clk), .D (signal_12637), .Q (signal_12638) ) ;
    buf_clk cell_10108 ( .C (clk), .D (signal_12653), .Q (signal_12654) ) ;
    buf_clk cell_10124 ( .C (clk), .D (signal_12669), .Q (signal_12670) ) ;
    buf_clk cell_10140 ( .C (clk), .D (signal_12685), .Q (signal_12686) ) ;
    buf_clk cell_10156 ( .C (clk), .D (signal_12701), .Q (signal_12702) ) ;
    buf_clk cell_10172 ( .C (clk), .D (signal_12717), .Q (signal_12718) ) ;
    buf_clk cell_10188 ( .C (clk), .D (signal_12733), .Q (signal_12734) ) ;
    buf_clk cell_10204 ( .C (clk), .D (signal_12749), .Q (signal_12750) ) ;
    buf_clk cell_10220 ( .C (clk), .D (signal_12765), .Q (signal_12766) ) ;
    buf_clk cell_10236 ( .C (clk), .D (signal_12781), .Q (signal_12782) ) ;
    buf_clk cell_10252 ( .C (clk), .D (signal_12797), .Q (signal_12798) ) ;
    buf_clk cell_10268 ( .C (clk), .D (signal_12813), .Q (signal_12814) ) ;
    buf_clk cell_10284 ( .C (clk), .D (signal_12829), .Q (signal_12830) ) ;
    buf_clk cell_10300 ( .C (clk), .D (signal_12845), .Q (signal_12846) ) ;
    buf_clk cell_10316 ( .C (clk), .D (signal_12861), .Q (signal_12862) ) ;
    buf_clk cell_10332 ( .C (clk), .D (signal_12877), .Q (signal_12878) ) ;
    buf_clk cell_10348 ( .C (clk), .D (signal_12893), .Q (signal_12894) ) ;
    buf_clk cell_10364 ( .C (clk), .D (signal_12909), .Q (signal_12910) ) ;
    buf_clk cell_10380 ( .C (clk), .D (signal_12925), .Q (signal_12926) ) ;
    buf_clk cell_10396 ( .C (clk), .D (signal_12941), .Q (signal_12942) ) ;
    buf_clk cell_10412 ( .C (clk), .D (signal_12957), .Q (signal_12958) ) ;
    buf_clk cell_10428 ( .C (clk), .D (signal_12973), .Q (signal_12974) ) ;
    buf_clk cell_10444 ( .C (clk), .D (signal_12989), .Q (signal_12990) ) ;
    buf_clk cell_10460 ( .C (clk), .D (signal_13005), .Q (signal_13006) ) ;
    buf_clk cell_10476 ( .C (clk), .D (signal_13021), .Q (signal_13022) ) ;
    buf_clk cell_10492 ( .C (clk), .D (signal_13037), .Q (signal_13038) ) ;
    buf_clk cell_10508 ( .C (clk), .D (signal_13053), .Q (signal_13054) ) ;
    buf_clk cell_10524 ( .C (clk), .D (signal_13069), .Q (signal_13070) ) ;
    buf_clk cell_10540 ( .C (clk), .D (signal_13085), .Q (signal_13086) ) ;
    buf_clk cell_10556 ( .C (clk), .D (signal_13101), .Q (signal_13102) ) ;
    buf_clk cell_10572 ( .C (clk), .D (signal_13117), .Q (signal_13118) ) ;
    buf_clk cell_10588 ( .C (clk), .D (signal_13133), .Q (signal_13134) ) ;
    buf_clk cell_10604 ( .C (clk), .D (signal_13149), .Q (signal_13150) ) ;
    buf_clk cell_10620 ( .C (clk), .D (signal_13165), .Q (signal_13166) ) ;
    buf_clk cell_10636 ( .C (clk), .D (signal_13181), .Q (signal_13182) ) ;
    buf_clk cell_10652 ( .C (clk), .D (signal_13197), .Q (signal_13198) ) ;
    buf_clk cell_10668 ( .C (clk), .D (signal_13213), .Q (signal_13214) ) ;
    buf_clk cell_10684 ( .C (clk), .D (signal_13229), .Q (signal_13230) ) ;
    buf_clk cell_10700 ( .C (clk), .D (signal_13245), .Q (signal_13246) ) ;
    buf_clk cell_10716 ( .C (clk), .D (signal_13261), .Q (signal_13262) ) ;
    buf_clk cell_10732 ( .C (clk), .D (signal_13277), .Q (signal_13278) ) ;
    buf_clk cell_10748 ( .C (clk), .D (signal_13293), .Q (signal_13294) ) ;
    buf_clk cell_10764 ( .C (clk), .D (signal_13309), .Q (signal_13310) ) ;
    buf_clk cell_10780 ( .C (clk), .D (signal_13325), .Q (signal_13326) ) ;
    buf_clk cell_10796 ( .C (clk), .D (signal_13341), .Q (signal_13342) ) ;
    buf_clk cell_10812 ( .C (clk), .D (signal_13357), .Q (signal_13358) ) ;
    buf_clk cell_10828 ( .C (clk), .D (signal_13373), .Q (signal_13374) ) ;
    buf_clk cell_10844 ( .C (clk), .D (signal_13389), .Q (signal_13390) ) ;
    buf_clk cell_10860 ( .C (clk), .D (signal_13405), .Q (signal_13406) ) ;
    buf_clk cell_10876 ( .C (clk), .D (signal_13421), .Q (signal_13422) ) ;
    buf_clk cell_10892 ( .C (clk), .D (signal_13437), .Q (signal_13438) ) ;
    buf_clk cell_10908 ( .C (clk), .D (signal_13453), .Q (signal_13454) ) ;
    buf_clk cell_10924 ( .C (clk), .D (signal_13469), .Q (signal_13470) ) ;
    buf_clk cell_10940 ( .C (clk), .D (signal_13485), .Q (signal_13486) ) ;
    buf_clk cell_10956 ( .C (clk), .D (signal_13501), .Q (signal_13502) ) ;
    buf_clk cell_10972 ( .C (clk), .D (signal_13517), .Q (signal_13518) ) ;
    buf_clk cell_10988 ( .C (clk), .D (signal_13533), .Q (signal_13534) ) ;
    buf_clk cell_11004 ( .C (clk), .D (signal_13549), .Q (signal_13550) ) ;
    buf_clk cell_11020 ( .C (clk), .D (signal_13565), .Q (signal_13566) ) ;
    buf_clk cell_11036 ( .C (clk), .D (signal_13581), .Q (signal_13582) ) ;
    buf_clk cell_11052 ( .C (clk), .D (signal_13597), .Q (signal_13598) ) ;
    buf_clk cell_11068 ( .C (clk), .D (signal_13613), .Q (signal_13614) ) ;
    buf_clk cell_11084 ( .C (clk), .D (signal_13629), .Q (signal_13630) ) ;
    buf_clk cell_11100 ( .C (clk), .D (signal_13645), .Q (signal_13646) ) ;
    buf_clk cell_11116 ( .C (clk), .D (signal_13661), .Q (signal_13662) ) ;
    buf_clk cell_11132 ( .C (clk), .D (signal_13677), .Q (signal_13678) ) ;
    buf_clk cell_11148 ( .C (clk), .D (signal_13693), .Q (signal_13694) ) ;
    buf_clk cell_11164 ( .C (clk), .D (signal_13709), .Q (signal_13710) ) ;
    buf_clk cell_11180 ( .C (clk), .D (signal_13725), .Q (signal_13726) ) ;
    buf_clk cell_11196 ( .C (clk), .D (signal_13741), .Q (signal_13742) ) ;
    buf_clk cell_11212 ( .C (clk), .D (signal_13757), .Q (signal_13758) ) ;
    buf_clk cell_11228 ( .C (clk), .D (signal_13773), .Q (signal_13774) ) ;
    buf_clk cell_11244 ( .C (clk), .D (signal_13789), .Q (signal_13790) ) ;
    buf_clk cell_11260 ( .C (clk), .D (signal_13805), .Q (signal_13806) ) ;
    buf_clk cell_11276 ( .C (clk), .D (signal_13821), .Q (signal_13822) ) ;
    buf_clk cell_11292 ( .C (clk), .D (signal_13837), .Q (signal_13838) ) ;
    buf_clk cell_11308 ( .C (clk), .D (signal_13853), .Q (signal_13854) ) ;
    buf_clk cell_11324 ( .C (clk), .D (signal_13869), .Q (signal_13870) ) ;
    buf_clk cell_11340 ( .C (clk), .D (signal_13885), .Q (signal_13886) ) ;
    buf_clk cell_11356 ( .C (clk), .D (signal_13901), .Q (signal_13902) ) ;
    buf_clk cell_11372 ( .C (clk), .D (signal_13917), .Q (signal_13918) ) ;
    buf_clk cell_11388 ( .C (clk), .D (signal_13933), .Q (signal_13934) ) ;
    buf_clk cell_11404 ( .C (clk), .D (signal_13949), .Q (signal_13950) ) ;
    buf_clk cell_11420 ( .C (clk), .D (signal_13965), .Q (signal_13966) ) ;
    buf_clk cell_11436 ( .C (clk), .D (signal_13981), .Q (signal_13982) ) ;
    buf_clk cell_11452 ( .C (clk), .D (signal_13997), .Q (signal_13998) ) ;
    buf_clk cell_11468 ( .C (clk), .D (signal_14013), .Q (signal_14014) ) ;
    buf_clk cell_11484 ( .C (clk), .D (signal_14029), .Q (signal_14030) ) ;
    buf_clk cell_11500 ( .C (clk), .D (signal_14045), .Q (signal_14046) ) ;
    buf_clk cell_11516 ( .C (clk), .D (signal_14061), .Q (signal_14062) ) ;
    buf_clk cell_11532 ( .C (clk), .D (signal_14077), .Q (signal_14078) ) ;
    buf_clk cell_11548 ( .C (clk), .D (signal_14093), .Q (signal_14094) ) ;
    buf_clk cell_11564 ( .C (clk), .D (signal_14109), .Q (signal_14110) ) ;
    buf_clk cell_11580 ( .C (clk), .D (signal_14125), .Q (signal_14126) ) ;
    buf_clk cell_11596 ( .C (clk), .D (signal_14141), .Q (signal_14142) ) ;
    buf_clk cell_11612 ( .C (clk), .D (signal_14157), .Q (signal_14158) ) ;
    buf_clk cell_11628 ( .C (clk), .D (signal_14173), .Q (signal_14174) ) ;
    buf_clk cell_11644 ( .C (clk), .D (signal_14189), .Q (signal_14190) ) ;
    buf_clk cell_11660 ( .C (clk), .D (signal_14205), .Q (signal_14206) ) ;
    buf_clk cell_11676 ( .C (clk), .D (signal_14221), .Q (signal_14222) ) ;
    buf_clk cell_11692 ( .C (clk), .D (signal_14237), .Q (signal_14238) ) ;
    buf_clk cell_11708 ( .C (clk), .D (signal_14253), .Q (signal_14254) ) ;
    buf_clk cell_11724 ( .C (clk), .D (signal_14269), .Q (signal_14270) ) ;
    buf_clk cell_11740 ( .C (clk), .D (signal_14285), .Q (signal_14286) ) ;
    buf_clk cell_11756 ( .C (clk), .D (signal_14301), .Q (signal_14302) ) ;
    buf_clk cell_11772 ( .C (clk), .D (signal_14317), .Q (signal_14318) ) ;
    buf_clk cell_11788 ( .C (clk), .D (signal_14333), .Q (signal_14334) ) ;
    buf_clk cell_11804 ( .C (clk), .D (signal_14349), .Q (signal_14350) ) ;
    buf_clk cell_11820 ( .C (clk), .D (signal_14365), .Q (signal_14366) ) ;
    buf_clk cell_11836 ( .C (clk), .D (signal_14381), .Q (signal_14382) ) ;
    buf_clk cell_11852 ( .C (clk), .D (signal_14397), .Q (signal_14398) ) ;
    buf_clk cell_11868 ( .C (clk), .D (signal_14413), .Q (signal_14414) ) ;
    buf_clk cell_11884 ( .C (clk), .D (signal_14429), .Q (signal_14430) ) ;
    buf_clk cell_11900 ( .C (clk), .D (signal_14445), .Q (signal_14446) ) ;
    buf_clk cell_11916 ( .C (clk), .D (signal_14461), .Q (signal_14462) ) ;
    buf_clk cell_11932 ( .C (clk), .D (signal_14477), .Q (signal_14478) ) ;
    buf_clk cell_11948 ( .C (clk), .D (signal_14493), .Q (signal_14494) ) ;
    buf_clk cell_11964 ( .C (clk), .D (signal_14509), .Q (signal_14510) ) ;
    buf_clk cell_11980 ( .C (clk), .D (signal_14525), .Q (signal_14526) ) ;
    buf_clk cell_11996 ( .C (clk), .D (signal_14541), .Q (signal_14542) ) ;
    buf_clk cell_12012 ( .C (clk), .D (signal_14557), .Q (signal_14558) ) ;
    buf_clk cell_12028 ( .C (clk), .D (signal_14573), .Q (signal_14574) ) ;
    buf_clk cell_12044 ( .C (clk), .D (signal_14589), .Q (signal_14590) ) ;
    buf_clk cell_12060 ( .C (clk), .D (signal_14605), .Q (signal_14606) ) ;
    buf_clk cell_12076 ( .C (clk), .D (signal_14621), .Q (signal_14622) ) ;
    buf_clk cell_12092 ( .C (clk), .D (signal_14637), .Q (signal_14638) ) ;
    buf_clk cell_12108 ( .C (clk), .D (signal_14653), .Q (signal_14654) ) ;
    buf_clk cell_12124 ( .C (clk), .D (signal_14669), .Q (signal_14670) ) ;
    buf_clk cell_12140 ( .C (clk), .D (signal_14685), .Q (signal_14686) ) ;
    buf_clk cell_12156 ( .C (clk), .D (signal_14701), .Q (signal_14702) ) ;
    buf_clk cell_12172 ( .C (clk), .D (signal_14717), .Q (signal_14718) ) ;
    buf_clk cell_12188 ( .C (clk), .D (signal_14733), .Q (signal_14734) ) ;
    buf_clk cell_12204 ( .C (clk), .D (signal_14749), .Q (signal_14750) ) ;
    buf_clk cell_12220 ( .C (clk), .D (signal_14765), .Q (signal_14766) ) ;
    buf_clk cell_12236 ( .C (clk), .D (signal_14781), .Q (signal_14782) ) ;
    buf_clk cell_12252 ( .C (clk), .D (signal_14797), .Q (signal_14798) ) ;
    buf_clk cell_12268 ( .C (clk), .D (signal_14813), .Q (signal_14814) ) ;
    buf_clk cell_12284 ( .C (clk), .D (signal_14829), .Q (signal_14830) ) ;
    buf_clk cell_12300 ( .C (clk), .D (signal_14845), .Q (signal_14846) ) ;
    buf_clk cell_12316 ( .C (clk), .D (signal_14861), .Q (signal_14862) ) ;
    buf_clk cell_12332 ( .C (clk), .D (signal_14877), .Q (signal_14878) ) ;
    buf_clk cell_12348 ( .C (clk), .D (signal_14893), .Q (signal_14894) ) ;
    buf_clk cell_12364 ( .C (clk), .D (signal_14909), .Q (signal_14910) ) ;
    buf_clk cell_12380 ( .C (clk), .D (signal_14925), .Q (signal_14926) ) ;
    buf_clk cell_12396 ( .C (clk), .D (signal_14941), .Q (signal_14942) ) ;

    /* register cells */
    DFF_X1 cell_33 ( .CK (clk), .D (signal_6990), .Q (signal_425), .QN () ) ;
    DFF_X1 cell_36 ( .CK (clk), .D (signal_7006), .Q (signal_426), .QN () ) ;
    DFF_X1 cell_39 ( .CK (clk), .D (signal_7022), .Q (signal_427), .QN () ) ;
    DFF_X1 cell_42 ( .CK (clk), .D (signal_7038), .Q (signal_428), .QN () ) ;
    DFF_X1 cell_45 ( .CK (clk), .D (signal_7054), .Q (signal_424), .QN () ) ;
    DFF_X1 cell_48 ( .CK (clk), .D (signal_7070), .Q (signal_421), .QN () ) ;
    DFF_X1 cell_51 ( .CK (clk), .D (signal_7086), .Q (signal_420), .QN () ) ;
    DFF_X1 cell_53 ( .CK (clk), .D (signal_7102), .Q (signal_418), .QN () ) ;
    DFF_X1 cell_55 ( .CK (clk), .D (signal_7118), .Q (signal_397), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_87 ( .clk (clk), .D ({signal_7150, signal_7134}), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_90 ( .clk (clk), .D ({signal_7182, signal_7166}), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_93 ( .clk (clk), .D ({signal_7214, signal_7198}), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_96 ( .clk (clk), .D ({signal_7246, signal_7230}), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_99 ( .clk (clk), .D ({signal_7278, signal_7262}), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_102 ( .clk (clk), .D ({signal_7310, signal_7294}), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_105 ( .clk (clk), .D ({signal_7342, signal_7326}), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_108 ( .clk (clk), .D ({signal_7374, signal_7358}), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_111 ( .clk (clk), .D ({signal_7406, signal_7390}), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_114 ( .clk (clk), .D ({signal_7438, signal_7422}), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_117 ( .clk (clk), .D ({signal_7470, signal_7454}), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_120 ( .clk (clk), .D ({signal_7502, signal_7486}), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_123 ( .clk (clk), .D ({signal_7534, signal_7518}), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_126 ( .clk (clk), .D ({signal_7566, signal_7550}), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_129 ( .clk (clk), .D ({signal_7598, signal_7582}), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_132 ( .clk (clk), .D ({signal_7630, signal_7614}), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_135 ( .clk (clk), .D ({signal_7662, signal_7646}), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_138 ( .clk (clk), .D ({signal_7694, signal_7678}), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_141 ( .clk (clk), .D ({signal_7726, signal_7710}), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_144 ( .clk (clk), .D ({signal_7758, signal_7742}), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_147 ( .clk (clk), .D ({signal_7790, signal_7774}), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_150 ( .clk (clk), .D ({signal_7822, signal_7806}), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_153 ( .clk (clk), .D ({signal_7854, signal_7838}), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_156 ( .clk (clk), .D ({signal_7886, signal_7870}), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_159 ( .clk (clk), .D ({signal_7918, signal_7902}), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_162 ( .clk (clk), .D ({signal_7950, signal_7934}), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_165 ( .clk (clk), .D ({signal_7982, signal_7966}), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_168 ( .clk (clk), .D ({signal_8014, signal_7998}), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_171 ( .clk (clk), .D ({signal_8046, signal_8030}), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_174 ( .clk (clk), .D ({signal_8078, signal_8062}), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_177 ( .clk (clk), .D ({signal_8110, signal_8094}), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_180 ( .clk (clk), .D ({signal_8142, signal_8126}), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_183 ( .clk (clk), .D ({signal_8174, signal_8158}), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_186 ( .clk (clk), .D ({signal_8206, signal_8190}), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_189 ( .clk (clk), .D ({signal_8238, signal_8222}), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_192 ( .clk (clk), .D ({signal_8270, signal_8254}), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_195 ( .clk (clk), .D ({signal_8302, signal_8286}), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_198 ( .clk (clk), .D ({signal_8334, signal_8318}), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_201 ( .clk (clk), .D ({signal_8366, signal_8350}), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_204 ( .clk (clk), .D ({signal_8398, signal_8382}), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_207 ( .clk (clk), .D ({signal_8430, signal_8414}), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_210 ( .clk (clk), .D ({signal_8462, signal_8446}), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_213 ( .clk (clk), .D ({signal_8494, signal_8478}), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_216 ( .clk (clk), .D ({signal_8526, signal_8510}), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_219 ( .clk (clk), .D ({signal_8558, signal_8542}), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_222 ( .clk (clk), .D ({signal_8590, signal_8574}), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_225 ( .clk (clk), .D ({signal_8622, signal_8606}), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_228 ( .clk (clk), .D ({signal_8654, signal_8638}), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_231 ( .clk (clk), .D ({signal_8686, signal_8670}), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_234 ( .clk (clk), .D ({signal_8718, signal_8702}), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_237 ( .clk (clk), .D ({signal_8750, signal_8734}), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_240 ( .clk (clk), .D ({signal_8782, signal_8766}), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_243 ( .clk (clk), .D ({signal_8814, signal_8798}), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_246 ( .clk (clk), .D ({signal_8846, signal_8830}), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_249 ( .clk (clk), .D ({signal_8878, signal_8862}), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_252 ( .clk (clk), .D ({signal_8910, signal_8894}), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_255 ( .clk (clk), .D ({signal_8942, signal_8926}), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_258 ( .clk (clk), .D ({signal_8974, signal_8958}), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_261 ( .clk (clk), .D ({signal_9006, signal_8990}), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_264 ( .clk (clk), .D ({signal_9038, signal_9022}), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_267 ( .clk (clk), .D ({signal_9070, signal_9054}), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_270 ( .clk (clk), .D ({signal_9102, signal_9086}), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_273 ( .clk (clk), .D ({signal_9134, signal_9118}), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_276 ( .clk (clk), .D ({signal_9166, signal_9150}), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_279 ( .clk (clk), .D ({signal_9198, signal_9182}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_282 ( .clk (clk), .D ({signal_9230, signal_9214}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_285 ( .clk (clk), .D ({signal_9262, signal_9246}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_288 ( .clk (clk), .D ({signal_9294, signal_9278}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_291 ( .clk (clk), .D ({signal_9326, signal_9310}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_294 ( .clk (clk), .D ({signal_9358, signal_9342}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_297 ( .clk (clk), .D ({signal_9390, signal_9374}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_300 ( .clk (clk), .D ({signal_9422, signal_9406}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_303 ( .clk (clk), .D ({signal_9454, signal_9438}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_306 ( .clk (clk), .D ({signal_9486, signal_9470}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_309 ( .clk (clk), .D ({signal_9518, signal_9502}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_312 ( .clk (clk), .D ({signal_9550, signal_9534}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_315 ( .clk (clk), .D ({signal_9582, signal_9566}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_318 ( .clk (clk), .D ({signal_9614, signal_9598}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_321 ( .clk (clk), .D ({signal_9646, signal_9630}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_324 ( .clk (clk), .D ({signal_9678, signal_9662}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_327 ( .clk (clk), .D ({signal_9710, signal_9694}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_330 ( .clk (clk), .D ({signal_9742, signal_9726}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_333 ( .clk (clk), .D ({signal_9774, signal_9758}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_336 ( .clk (clk), .D ({signal_9806, signal_9790}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_339 ( .clk (clk), .D ({signal_9838, signal_9822}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_342 ( .clk (clk), .D ({signal_9870, signal_9854}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_345 ( .clk (clk), .D ({signal_9902, signal_9886}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_348 ( .clk (clk), .D ({signal_9934, signal_9918}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_351 ( .clk (clk), .D ({signal_9966, signal_9950}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_354 ( .clk (clk), .D ({signal_9998, signal_9982}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_357 ( .clk (clk), .D ({signal_10030, signal_10014}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_360 ( .clk (clk), .D ({signal_10062, signal_10046}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_363 ( .clk (clk), .D ({signal_10094, signal_10078}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_366 ( .clk (clk), .D ({signal_10126, signal_10110}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_369 ( .clk (clk), .D ({signal_10158, signal_10142}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_372 ( .clk (clk), .D ({signal_10190, signal_10174}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_375 ( .clk (clk), .D ({signal_10222, signal_10206}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_378 ( .clk (clk), .D ({signal_10254, signal_10238}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_381 ( .clk (clk), .D ({signal_10286, signal_10270}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_384 ( .clk (clk), .D ({signal_10318, signal_10302}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_387 ( .clk (clk), .D ({signal_10350, signal_10334}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_390 ( .clk (clk), .D ({signal_10382, signal_10366}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_393 ( .clk (clk), .D ({signal_10414, signal_10398}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_396 ( .clk (clk), .D ({signal_10446, signal_10430}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_399 ( .clk (clk), .D ({signal_10478, signal_10462}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_402 ( .clk (clk), .D ({signal_10510, signal_10494}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_405 ( .clk (clk), .D ({signal_10542, signal_10526}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_408 ( .clk (clk), .D ({signal_10574, signal_10558}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_411 ( .clk (clk), .D ({signal_10606, signal_10590}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_414 ( .clk (clk), .D ({signal_10638, signal_10622}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_417 ( .clk (clk), .D ({signal_10670, signal_10654}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_420 ( .clk (clk), .D ({signal_10702, signal_10686}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_423 ( .clk (clk), .D ({signal_10734, signal_10718}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_426 ( .clk (clk), .D ({signal_10766, signal_10750}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_429 ( .clk (clk), .D ({signal_10798, signal_10782}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_432 ( .clk (clk), .D ({signal_10830, signal_10814}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_435 ( .clk (clk), .D ({signal_10862, signal_10846}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_438 ( .clk (clk), .D ({signal_10894, signal_10878}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_441 ( .clk (clk), .D ({signal_10926, signal_10910}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_444 ( .clk (clk), .D ({signal_10958, signal_10942}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_447 ( .clk (clk), .D ({signal_4244, signal_705}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_450 ( .clk (clk), .D ({signal_4245, signal_707}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_453 ( .clk (clk), .D ({signal_4246, signal_709}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_456 ( .clk (clk), .D ({signal_4247, signal_711}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_459 ( .clk (clk), .D ({signal_4248, signal_713}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_462 ( .clk (clk), .D ({signal_4249, signal_715}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_465 ( .clk (clk), .D ({signal_4250, signal_717}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_468 ( .clk (clk), .D ({signal_4251, signal_719}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_717 ( .clk (clk), .D ({signal_10990, signal_10974}), .Q ({signal_2406, signal_1493}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_721 ( .clk (clk), .D ({signal_11022, signal_11006}), .Q ({signal_2409, signal_1492}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_725 ( .clk (clk), .D ({signal_11054, signal_11038}), .Q ({signal_2412, signal_1491}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_729 ( .clk (clk), .D ({signal_11086, signal_11070}), .Q ({signal_2415, signal_1490}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_733 ( .clk (clk), .D ({signal_11118, signal_11102}), .Q ({signal_2418, signal_1489}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_737 ( .clk (clk), .D ({signal_11150, signal_11134}), .Q ({signal_2421, signal_1488}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_741 ( .clk (clk), .D ({signal_11182, signal_11166}), .Q ({signal_2424, signal_1487}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_745 ( .clk (clk), .D ({signal_11214, signal_11198}), .Q ({signal_2427, signal_1486}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_749 ( .clk (clk), .D ({signal_11246, signal_11230}), .Q ({signal_2443, signal_758}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_753 ( .clk (clk), .D ({signal_11278, signal_11262}), .Q ({signal_2441, signal_759}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_757 ( .clk (clk), .D ({signal_11310, signal_11294}), .Q ({signal_2439, signal_760}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_761 ( .clk (clk), .D ({signal_11342, signal_11326}), .Q ({signal_2437, signal_761}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_765 ( .clk (clk), .D ({signal_11374, signal_11358}), .Q ({signal_2435, signal_762}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_769 ( .clk (clk), .D ({signal_11406, signal_11390}), .Q ({signal_2433, signal_763}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_773 ( .clk (clk), .D ({signal_11438, signal_11422}), .Q ({signal_2431, signal_764}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_777 ( .clk (clk), .D ({signal_11470, signal_11454}), .Q ({signal_2429, signal_765}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_781 ( .clk (clk), .D ({signal_11502, signal_11486}), .Q ({signal_2866, signal_1909}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_785 ( .clk (clk), .D ({signal_11534, signal_11518}), .Q ({signal_2869, signal_1908}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_789 ( .clk (clk), .D ({signal_11566, signal_11550}), .Q ({signal_2872, signal_1907}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_793 ( .clk (clk), .D ({signal_11598, signal_11582}), .Q ({signal_2875, signal_1906}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_797 ( .clk (clk), .D ({signal_11630, signal_11614}), .Q ({signal_2878, signal_1905}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_801 ( .clk (clk), .D ({signal_11662, signal_11646}), .Q ({signal_2881, signal_1904}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_805 ( .clk (clk), .D ({signal_11694, signal_11678}), .Q ({signal_2884, signal_1903}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_809 ( .clk (clk), .D ({signal_11726, signal_11710}), .Q ({signal_2887, signal_1902}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_813 ( .clk (clk), .D ({signal_11758, signal_11742}), .Q ({signal_2890, signal_1893}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_817 ( .clk (clk), .D ({signal_11790, signal_11774}), .Q ({signal_2893, signal_1892}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_821 ( .clk (clk), .D ({signal_11822, signal_11806}), .Q ({signal_2896, signal_1891}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_825 ( .clk (clk), .D ({signal_11854, signal_11838}), .Q ({signal_2899, signal_1890}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_829 ( .clk (clk), .D ({signal_11886, signal_11870}), .Q ({signal_2902, signal_1889}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_833 ( .clk (clk), .D ({signal_11918, signal_11902}), .Q ({signal_2905, signal_1888}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_837 ( .clk (clk), .D ({signal_11950, signal_11934}), .Q ({signal_2908, signal_1887}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_841 ( .clk (clk), .D ({signal_11982, signal_11966}), .Q ({signal_2911, signal_1886}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_845 ( .clk (clk), .D ({signal_12014, signal_11998}), .Q ({signal_2914, signal_1877}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_849 ( .clk (clk), .D ({signal_12046, signal_12030}), .Q ({signal_2917, signal_1876}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_853 ( .clk (clk), .D ({signal_12078, signal_12062}), .Q ({signal_2920, signal_1875}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_857 ( .clk (clk), .D ({signal_12110, signal_12094}), .Q ({signal_2923, signal_1874}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_861 ( .clk (clk), .D ({signal_12142, signal_12126}), .Q ({signal_2926, signal_1873}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_865 ( .clk (clk), .D ({signal_12174, signal_12158}), .Q ({signal_2929, signal_1872}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_869 ( .clk (clk), .D ({signal_12206, signal_12190}), .Q ({signal_2932, signal_1871}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_873 ( .clk (clk), .D ({signal_12238, signal_12222}), .Q ({signal_2935, signal_1870}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_877 ( .clk (clk), .D ({signal_12270, signal_12254}), .Q ({signal_2938, signal_1861}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_881 ( .clk (clk), .D ({signal_12302, signal_12286}), .Q ({signal_2941, signal_1860}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_885 ( .clk (clk), .D ({signal_12334, signal_12318}), .Q ({signal_2944, signal_1859}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_889 ( .clk (clk), .D ({signal_12366, signal_12350}), .Q ({signal_2947, signal_1858}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_893 ( .clk (clk), .D ({signal_12398, signal_12382}), .Q ({signal_2950, signal_1857}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_897 ( .clk (clk), .D ({signal_12430, signal_12414}), .Q ({signal_2953, signal_1856}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_901 ( .clk (clk), .D ({signal_12462, signal_12446}), .Q ({signal_2956, signal_1855}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_905 ( .clk (clk), .D ({signal_12494, signal_12478}), .Q ({signal_2959, signal_1854}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_909 ( .clk (clk), .D ({signal_12526, signal_12510}), .Q ({signal_2962, signal_1845}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_913 ( .clk (clk), .D ({signal_12558, signal_12542}), .Q ({signal_2965, signal_1844}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_917 ( .clk (clk), .D ({signal_12590, signal_12574}), .Q ({signal_2968, signal_1843}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_921 ( .clk (clk), .D ({signal_12622, signal_12606}), .Q ({signal_2971, signal_1842}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_925 ( .clk (clk), .D ({signal_12654, signal_12638}), .Q ({signal_2974, signal_1841}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_929 ( .clk (clk), .D ({signal_12686, signal_12670}), .Q ({signal_2977, signal_1840}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_933 ( .clk (clk), .D ({signal_12718, signal_12702}), .Q ({signal_2980, signal_1839}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_937 ( .clk (clk), .D ({signal_12750, signal_12734}), .Q ({signal_2983, signal_1838}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_941 ( .clk (clk), .D ({signal_12782, signal_12766}), .Q ({signal_2986, signal_1509}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_945 ( .clk (clk), .D ({signal_12814, signal_12798}), .Q ({signal_2989, signal_1508}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_949 ( .clk (clk), .D ({signal_12846, signal_12830}), .Q ({signal_2992, signal_1507}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_953 ( .clk (clk), .D ({signal_12878, signal_12862}), .Q ({signal_2995, signal_1506}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_957 ( .clk (clk), .D ({signal_12910, signal_12894}), .Q ({signal_2998, signal_1505}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_961 ( .clk (clk), .D ({signal_12942, signal_12926}), .Q ({signal_3001, signal_1504}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_965 ( .clk (clk), .D ({signal_12974, signal_12958}), .Q ({signal_3004, signal_1503}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_969 ( .clk (clk), .D ({signal_13006, signal_12990}), .Q ({signal_3007, signal_1502}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_973 ( .clk (clk), .D ({signal_13038, signal_13022}), .Q ({signal_3010, signal_1821}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_977 ( .clk (clk), .D ({signal_13070, signal_13054}), .Q ({signal_3013, signal_1820}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_981 ( .clk (clk), .D ({signal_13102, signal_13086}), .Q ({signal_3016, signal_1819}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_985 ( .clk (clk), .D ({signal_13134, signal_13118}), .Q ({signal_3019, signal_1818}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_989 ( .clk (clk), .D ({signal_13166, signal_13150}), .Q ({signal_3022, signal_1817}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_993 ( .clk (clk), .D ({signal_13198, signal_13182}), .Q ({signal_3025, signal_1816}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_997 ( .clk (clk), .D ({signal_13230, signal_13214}), .Q ({signal_3028, signal_1815}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1001 ( .clk (clk), .D ({signal_13262, signal_13246}), .Q ({signal_3031, signal_1814}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1005 ( .clk (clk), .D ({signal_13294, signal_13278}), .Q ({signal_3034, signal_1805}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1009 ( .clk (clk), .D ({signal_13326, signal_13310}), .Q ({signal_3037, signal_1804}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1013 ( .clk (clk), .D ({signal_13358, signal_13342}), .Q ({signal_3040, signal_1803}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1017 ( .clk (clk), .D ({signal_13390, signal_13374}), .Q ({signal_3043, signal_1802}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1021 ( .clk (clk), .D ({signal_13422, signal_13406}), .Q ({signal_3046, signal_1801}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1025 ( .clk (clk), .D ({signal_13454, signal_13438}), .Q ({signal_3049, signal_1800}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1029 ( .clk (clk), .D ({signal_13486, signal_13470}), .Q ({signal_3052, signal_1799}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1033 ( .clk (clk), .D ({signal_13518, signal_13502}), .Q ({signal_3055, signal_1798}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1037 ( .clk (clk), .D ({signal_13550, signal_13534}), .Q ({signal_3058, signal_1789}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1041 ( .clk (clk), .D ({signal_13582, signal_13566}), .Q ({signal_3061, signal_1788}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1045 ( .clk (clk), .D ({signal_13614, signal_13598}), .Q ({signal_3064, signal_1787}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1049 ( .clk (clk), .D ({signal_13646, signal_13630}), .Q ({signal_3067, signal_1786}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1053 ( .clk (clk), .D ({signal_13678, signal_13662}), .Q ({signal_3070, signal_1785}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1057 ( .clk (clk), .D ({signal_13710, signal_13694}), .Q ({signal_3073, signal_1784}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1061 ( .clk (clk), .D ({signal_13742, signal_13726}), .Q ({signal_3076, signal_1783}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1065 ( .clk (clk), .D ({signal_13774, signal_13758}), .Q ({signal_3079, signal_1782}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1069 ( .clk (clk), .D ({signal_13806, signal_13790}), .Q ({signal_3082, signal_1773}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1073 ( .clk (clk), .D ({signal_13838, signal_13822}), .Q ({signal_3085, signal_1772}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1077 ( .clk (clk), .D ({signal_13870, signal_13854}), .Q ({signal_3088, signal_1771}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1081 ( .clk (clk), .D ({signal_13902, signal_13886}), .Q ({signal_3091, signal_1770}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1085 ( .clk (clk), .D ({signal_13934, signal_13918}), .Q ({signal_3094, signal_1769}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1089 ( .clk (clk), .D ({signal_13966, signal_13950}), .Q ({signal_3097, signal_1768}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1093 ( .clk (clk), .D ({signal_13998, signal_13982}), .Q ({signal_3100, signal_1767}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1097 ( .clk (clk), .D ({signal_14030, signal_14014}), .Q ({signal_3103, signal_1766}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1101 ( .clk (clk), .D ({signal_4252, signal_1054}), .Q ({signal_3106, signal_1749}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1105 ( .clk (clk), .D ({signal_4253, signal_1057}), .Q ({signal_3109, signal_1748}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1109 ( .clk (clk), .D ({signal_4254, signal_1060}), .Q ({signal_3112, signal_1747}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1113 ( .clk (clk), .D ({signal_4255, signal_1063}), .Q ({signal_3115, signal_1746}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1117 ( .clk (clk), .D ({signal_4256, signal_1066}), .Q ({signal_3118, signal_1745}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1121 ( .clk (clk), .D ({signal_4257, signal_1069}), .Q ({signal_3121, signal_1744}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1125 ( .clk (clk), .D ({signal_4258, signal_1072}), .Q ({signal_3124, signal_1743}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1129 ( .clk (clk), .D ({signal_4259, signal_1075}), .Q ({signal_3127, signal_1742}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1133 ( .clk (clk), .D ({signal_14062, signal_14046}), .Q ({signal_3130, signal_1733}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1137 ( .clk (clk), .D ({signal_14094, signal_14078}), .Q ({signal_3133, signal_1732}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1141 ( .clk (clk), .D ({signal_14126, signal_14110}), .Q ({signal_3136, signal_1731}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1145 ( .clk (clk), .D ({signal_14158, signal_14142}), .Q ({signal_3139, signal_1730}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1149 ( .clk (clk), .D ({signal_14190, signal_14174}), .Q ({signal_3142, signal_1729}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1153 ( .clk (clk), .D ({signal_14222, signal_14206}), .Q ({signal_3145, signal_1728}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1157 ( .clk (clk), .D ({signal_14254, signal_14238}), .Q ({signal_3148, signal_1727}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1161 ( .clk (clk), .D ({signal_14286, signal_14270}), .Q ({signal_3151, signal_1726}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1165 ( .clk (clk), .D ({signal_14318, signal_14302}), .Q ({signal_3154, signal_1717}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1169 ( .clk (clk), .D ({signal_14350, signal_14334}), .Q ({signal_3157, signal_1716}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1173 ( .clk (clk), .D ({signal_14382, signal_14366}), .Q ({signal_3160, signal_1715}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1177 ( .clk (clk), .D ({signal_14414, signal_14398}), .Q ({signal_3163, signal_1714}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1181 ( .clk (clk), .D ({signal_14446, signal_14430}), .Q ({signal_3166, signal_1713}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1185 ( .clk (clk), .D ({signal_14478, signal_14462}), .Q ({signal_3169, signal_1712}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1189 ( .clk (clk), .D ({signal_14510, signal_14494}), .Q ({signal_3172, signal_1711}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1193 ( .clk (clk), .D ({signal_14542, signal_14526}), .Q ({signal_3175, signal_1710}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1197 ( .clk (clk), .D ({signal_14574, signal_14558}), .Q ({signal_3178, signal_1701}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1201 ( .clk (clk), .D ({signal_14606, signal_14590}), .Q ({signal_3181, signal_1700}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1205 ( .clk (clk), .D ({signal_14638, signal_14622}), .Q ({signal_3184, signal_1699}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1209 ( .clk (clk), .D ({signal_14670, signal_14654}), .Q ({signal_3187, signal_1698}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1213 ( .clk (clk), .D ({signal_14702, signal_14686}), .Q ({signal_3190, signal_1697}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1217 ( .clk (clk), .D ({signal_14734, signal_14718}), .Q ({signal_3193, signal_1696}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1221 ( .clk (clk), .D ({signal_14766, signal_14750}), .Q ({signal_3196, signal_1695}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1225 ( .clk (clk), .D ({signal_14798, signal_14782}), .Q ({signal_3199, signal_1694}) ) ;
    DFF_X1 cell_1561 ( .CK (clk), .D (signal_14814), .Q (signal_1268), .QN () ) ;
    DFF_X1 cell_1563 ( .CK (clk), .D (signal_14830), .Q (signal_1269), .QN () ) ;
    DFF_X1 cell_1565 ( .CK (clk), .D (signal_14846), .Q (signal_1270), .QN () ) ;
    DFF_X1 cell_1567 ( .CK (clk), .D (signal_14862), .Q (signal_1271), .QN () ) ;
    DFF_X1 cell_1569 ( .CK (clk), .D (signal_14878), .Q (signal_1272), .QN () ) ;
    DFF_X1 cell_1571 ( .CK (clk), .D (signal_14894), .Q (signal_1273), .QN () ) ;
    DFF_X1 cell_1573 ( .CK (clk), .D (signal_14910), .Q (signal_1274), .QN () ) ;
    DFF_X1 cell_1575 ( .CK (clk), .D (signal_14926), .Q (signal_1254), .QN () ) ;
    DFF_X1 cell_1713 ( .CK (clk), .D (signal_14942), .Q (signal_393), .QN () ) ;
endmodule
