module Reg1(x, y);
 input [74:0] x;
 output [73:0] y;

  register_stage #(.WIDTH(74)) inst_0(.clk(x[71]), .D({x[72],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[73],x[74],x[0],x[11],x[22],x[33],x[44],x[55],x[60],x[61],x[62],x[63],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[56],x[57],x[58],x[59]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73]}));
endmodule

module Reg2(x, y);
 input [130:0] x;
 output [129:0] y;

  register_stage #(.WIDTH(130)) inst_0(.clk(x[115]), .D({x[116],x[117],x[118],x[119],x[120],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[0],x[1],x[2],x[3],x[4],x[55],x[56],x[57],x[58],x[59],x[75],x[76],x[77],x[78],x[79],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [173:0] x;
 output [99:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx29 Fx29_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx30 Fx30_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx34 Fx34_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx35 Fx35_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx39 Fx39_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx40 Fx40_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx44 Fx44_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx45 Fx45_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx49 Fx49_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx50 Fx50_inst(.x({x[34], x[33], x[32], x[31], x[30]}), .y(y[20]));
  Fx51 Fx51_inst(.x({x[35], x[33]}), .y(y[21]));
  Fx52 Fx52_inst(.x({x[36], x[32]}), .y(y[22]));
  Fx53 Fx53_inst(.x({x[37], x[31]}), .y(y[23]));
  Fx54 Fx54_inst(.x({x[38], x[30]}), .y(y[24]));
  Fx55 Fx55_inst(.x({x[43], x[42], x[41], x[40], x[39]}), .y(y[25]));
  Fx56 Fx56_inst(.x({x[44], x[42]}), .y(y[26]));
  Fx57 Fx57_inst(.x({x[45], x[41]}), .y(y[27]));
  Fx58 Fx58_inst(.x({x[46], x[40]}), .y(y[28]));
  Fx59 Fx59_inst(.x({x[47], x[39]}), .y(y[29]));
  Fx60 Fx60_inst(.x({x[52], x[51], x[50], x[49], x[48]}), .y(y[30]));
  Fx61 Fx61_inst(.x({x[53], x[51]}), .y(y[31]));
  Fx62 Fx62_inst(.x({x[54], x[50]}), .y(y[32]));
  Fx63 Fx63_inst(.x({x[55], x[49]}), .y(y[33]));
  Fx64 Fx64_inst(.x({x[56], x[48]}), .y(y[34]));
  Fx65 Fx65_inst(.x({x[61], x[60], x[59], x[58], x[57]}), .y(y[35]));
  Fx66 Fx66_inst(.x({x[62], x[60]}), .y(y[36]));
  Fx67 Fx67_inst(.x({x[63], x[59]}), .y(y[37]));
  Fx68 Fx68_inst(.x({x[64], x[58]}), .y(y[38]));
  Fx69 Fx69_inst(.x({x[65], x[57]}), .y(y[39]));
  Fx70 Fx70_inst(.x({x[70], x[69], x[68], x[67], x[66]}), .y(y[40]));
  Fx71 Fx71_inst(.x({x[71], x[69]}), .y(y[41]));
  Fx72 Fx72_inst(.x({x[72], x[68]}), .y(y[42]));
  Fx73 Fx73_inst(.x({x[73], x[67]}), .y(y[43]));
  Fx74 Fx74_inst(.x({x[74], x[66]}), .y(y[44]));
  Fx75 Fx75_inst(.x({x[79], x[78], x[77], x[76], x[75]}), .y(y[45]));
  Fx76 Fx76_inst(.x({x[80], x[78]}), .y(y[46]));
  Fx77 Fx77_inst(.x({x[81], x[77]}), .y(y[47]));
  Fx78 Fx78_inst(.x({x[82], x[76]}), .y(y[48]));
  Fx79 Fx79_inst(.x({x[83], x[75]}), .y(y[49]));
  Fx80 Fx80_inst(.x({x[88], x[87], x[86], x[85], x[84]}), .y(y[50]));
  Fx81 Fx81_inst(.x({x[89], x[87]}), .y(y[51]));
  Fx82 Fx82_inst(.x({x[90], x[86]}), .y(y[52]));
  Fx83 Fx83_inst(.x({x[91], x[85]}), .y(y[53]));
  Fx84 Fx84_inst(.x({x[92], x[84]}), .y(y[54]));
  Fx85 Fx85_inst(.x({x[97], x[96], x[95], x[94], x[93]}), .y(y[55]));
  Fx86 Fx86_inst(.x({x[98], x[96]}), .y(y[56]));
  Fx87 Fx87_inst(.x({x[99], x[95]}), .y(y[57]));
  Fx88 Fx88_inst(.x({x[100], x[94]}), .y(y[58]));
  Fx89 Fx89_inst(.x({x[101], x[93]}), .y(y[59]));
  Fx90 Fx90_inst(.x({x[106], x[105], x[104], x[103], x[102]}), .y(y[60]));
  Fx91 Fx91_inst(.x({x[107], x[105]}), .y(y[61]));
  Fx92 Fx92_inst(.x({x[108], x[104]}), .y(y[62]));
  Fx93 Fx93_inst(.x({x[109], x[103]}), .y(y[63]));
  Fx94 Fx94_inst(.x({x[110], x[102]}), .y(y[64]));
  Fx95 Fx95_inst(.x({x[115], x[114], x[113], x[112], x[111]}), .y(y[65]));
  Fx96 Fx96_inst(.x({x[116], x[114]}), .y(y[66]));
  Fx97 Fx97_inst(.x({x[117], x[113]}), .y(y[67]));
  Fx98 Fx98_inst(.x({x[118], x[112]}), .y(y[68]));
  Fx99 Fx99_inst(.x({x[119], x[111]}), .y(y[69]));
  Fx100 Fx100_inst(.x({x[124], x[123], x[122], x[121], x[120]}), .y(y[70]));
  Fx101 Fx101_inst(.x({x[125], x[123]}), .y(y[71]));
  Fx102 Fx102_inst(.x({x[126], x[122]}), .y(y[72]));
  Fx103 Fx103_inst(.x({x[127], x[121]}), .y(y[73]));
  Fx104 Fx104_inst(.x({x[128], x[120]}), .y(y[74]));
  Fx105 Fx105_inst(.x({x[133], x[132], x[131], x[130], x[129]}), .y(y[75]));
  Fx106 Fx106_inst(.x({x[134], x[132]}), .y(y[76]));
  Fx107 Fx107_inst(.x({x[135], x[131]}), .y(y[77]));
  Fx108 Fx108_inst(.x({x[136], x[130]}), .y(y[78]));
  Fx109 Fx109_inst(.x({x[137], x[129]}), .y(y[79]));
  Fx110 Fx110_inst(.x({x[142], x[141], x[140], x[139], x[138]}), .y(y[80]));
  Fx111 Fx111_inst(.x({x[143], x[141]}), .y(y[81]));
  Fx112 Fx112_inst(.x({x[144], x[140]}), .y(y[82]));
  Fx113 Fx113_inst(.x({x[145], x[139]}), .y(y[83]));
  Fx114 Fx114_inst(.x({x[146], x[138]}), .y(y[84]));
  Fx115 Fx115_inst(.x({x[151], x[150], x[149], x[148], x[147]}), .y(y[85]));
  Fx116 Fx116_inst(.x({x[152], x[150]}), .y(y[86]));
  Fx117 Fx117_inst(.x({x[153], x[149]}), .y(y[87]));
  Fx118 Fx118_inst(.x({x[154], x[148]}), .y(y[88]));
  Fx119 Fx119_inst(.x({x[155], x[147]}), .y(y[89]));
  Fx120 Fx120_inst(.x({x[160], x[159], x[158], x[157], x[156]}), .y(y[90]));
  Fx121 Fx121_inst(.x({x[161], x[159]}), .y(y[91]));
  Fx122 Fx122_inst(.x({x[162], x[158]}), .y(y[92]));
  Fx123 Fx123_inst(.x({x[163], x[157]}), .y(y[93]));
  Fx124 Fx124_inst(.x({x[164], x[156]}), .y(y[94]));
  Fx125 Fx125_inst(.x({x[169], x[168], x[167], x[166], x[165]}), .y(y[95]));
  Fx126 Fx126_inst(.x({x[170], x[168]}), .y(y[96]));
  Fx127 Fx127_inst(.x({x[171], x[167]}), .y(y[97]));
  Fx128 Fx128_inst(.x({x[172], x[166]}), .y(y[98]));
  Fx129 Fx129_inst(.x({x[173], x[165]}), .y(y[99]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [21:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~x[0] & t[12];
  assign t[10] = ~x[0] & t[17];
  assign t[11] = ~x[0] & t[18];
  assign t[12] = t[19] ^ x[3];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = t[21] ^ x[9];
  assign t[15] = t[22] ^ x[12];
  assign t[16] = t[23] ^ x[15];
  assign t[17] = t[24] ^ x[18];
  assign t[18] = t[25] ^ x[21];
  assign t[19] = (x[1] & x[2]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[20] = (x[4] & x[5]);
  assign t[21] = (x[7] & x[8]);
  assign t[22] = (x[10] & x[11]);
  assign t[23] = (x[13] & x[14]);
  assign t[24] = (x[16] & x[17]);
  assign t[25] = (x[19] & x[20]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[7]);
  assign t[4] = ~(~x[0] & ~t[13]);
  assign t[5] = ~x[0] & t[14];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~x[0] & t[15];
  assign t[9] = ~(~x[0] & ~t[16]);
  assign y = t[0] & t[1];
endmodule

module R1ind66(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(t[0]);
endmodule

module R1ind67(x, y);
 input [6:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[2];
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = t[5] ^ x[3];
  assign t[4] = t[6] ^ x[6];
  assign t[5] = (x[1] & x[2]);
  assign t[6] = (x[4] & x[5]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind68(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~x[0] & t[2];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = t[4] ^ x[3];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[1] & x[2]);
  assign t[5] = (x[4] & x[5]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind73(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind74(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~(~x[0] & ~t[2]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = t[4] ^ x[3];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[1] & x[2]);
  assign t[5] = (x[4] & x[5]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [15:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[13];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[7] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[12]);
  assign t[21] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[13] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] | t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind76(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind77(x, y);
 input [15:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[13];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[7] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[12]);
  assign t[21] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind78(x, y);
 input [15:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[4] & x[10]);
  assign t[21] = (x[4] & x[12]);
  assign t[22] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind79(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind80(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind81(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind82(x, y);
 input [15:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[4] & x[10]);
  assign t[21] = (x[4] & x[12]);
  assign t[22] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind83(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind84(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind85(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind86(x, y);
 input [15:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[4] & x[10]);
  assign t[21] = (x[4] & x[12]);
  assign t[22] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind87(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind88(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind89(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind90(x, y);
 input [15:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[4] & x[10]);
  assign t[21] = (x[4] & x[12]);
  assign t[22] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind91(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind92(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind93(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind94(x, y);
 input [15:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[4] & x[10]);
  assign t[21] = (x[4] & x[12]);
  assign t[22] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind95(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind96(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind97(x, y);
 input [15:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[13];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[7] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[12]);
  assign t[21] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind98(x, y);
 input [15:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15]);
  assign t[11] = t[16] ^ x[6];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[13];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[7] & x[10]);
  assign t[19] = (x[7] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[11];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = t[9] | t[12];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[10] | t[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind99(x, y);
 input [15:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[13];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[7] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[12]);
  assign t[21] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[13] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] | t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind100(x, y);
 input [13:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~t[2];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[9];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = t[17] ^ x[13];
  assign t[14] = (x[4] & x[5]);
  assign t[15] = (x[7] & x[8]);
  assign t[16] = (x[7] & x[10]);
  assign t[17] = (x[7] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[10];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[11] & t[7]);
  assign t[6] = ~(t[12] & t[8]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[13] & t[9]);
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind101(x, y);
 input [15:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[11];
  assign t[15] = t[20] ^ x[13];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[7] & x[10]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[12]);
  assign t[21] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind102(x, y);
 input [15:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15]);
  assign t[11] = t[16] ^ x[6];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[13];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[7] & x[10]);
  assign t[19] = (x[7] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[11];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = t[9] | t[12];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[10] | t[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind103(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind104(x, y);
 input [13:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[4] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[4] & x[12]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind105(x, y);
 input [15:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[13];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[4] & x[10]);
  assign t[22] = (x[4] & x[12]);
  assign t[23] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind106(x, y);
 input [15:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = t[21] ^ x[13];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[4] & x[10]);
  assign t[21] = (x[4] & x[12]);
  assign t[22] = (x[4] & x[14]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind107(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[26] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[27] | t[20]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[15];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[19];
  assign t[31] = t[40] ^ x[21];
  assign t[32] = t[41] ^ x[23];
  assign t[33] = t[42] ^ x[25];
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[8] & x[9]);
  assign t[36] = (x[11] & x[12]);
  assign t[37] = (x[8] & x[14]);
  assign t[38] = (x[8] & x[16]);
  assign t[39] = (x[11] & x[18]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[11] & x[20]);
  assign t[41] = (x[8] & x[22]);
  assign t[42] = (x[11] & x[24]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind108(x, y);
 input [21:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[21] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[24] & t[17]);
  assign t[15] = ~(t[25]);
  assign t[16] = ~(t[25] & t[18]);
  assign t[17] = ~(t[20]);
  assign t[18] = ~(t[22]);
  assign t[19] = t[26] ^ x[5];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = t[27] ^ x[10];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[15];
  assign t[23] = t[30] ^ x[17];
  assign t[24] = t[31] ^ x[19];
  assign t[25] = t[32] ^ x[21];
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[8] & x[9]);
  assign t[28] = (x[8] & x[11]);
  assign t[29] = (x[13] & x[14]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[13] & x[16]);
  assign t[31] = (x[8] & x[18]);
  assign t[32] = (x[13] & x[20]);
  assign t[3] = ~x[2] & t[19];
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[6] : t[7];
  assign t[6] = x[2] ? x[7] : t[8];
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[20] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind109(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[26]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[29] & t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[31] & t[30]);
  assign t[24] = ~(t[33]);
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[15];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[19];
  assign t[31] = t[40] ^ x[21];
  assign t[32] = t[41] ^ x[23];
  assign t[33] = t[42] ^ x[25];
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[8] & x[9]);
  assign t[36] = (x[11] & x[12]);
  assign t[37] = (x[8] & x[14]);
  assign t[38] = (x[8] & x[16]);
  assign t[39] = (x[11] & x[18]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[11] & x[20]);
  assign t[41] = (x[8] & x[22]);
  assign t[42] = (x[11] & x[24]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind110(x, y);
 input [25:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = t[17] | t[24];
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = t[20] | t[25];
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[21] | t[15]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[29]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[22] | t[18]);
  assign t[21] = ~(t[30]);
  assign t[22] = ~(t[31]);
  assign t[23] = t[32] ^ x[7];
  assign t[24] = t[33] ^ x[10];
  assign t[25] = t[34] ^ x[13];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[17];
  assign t[28] = t[37] ^ x[19];
  assign t[29] = t[38] ^ x[21];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[23];
  assign t[31] = t[40] ^ x[25];
  assign t[32] = (x[5] & x[6]);
  assign t[33] = (x[8] & x[9]);
  assign t[34] = (x[11] & x[12]);
  assign t[35] = (x[8] & x[14]);
  assign t[36] = (x[8] & x[16]);
  assign t[37] = (x[11] & x[18]);
  assign t[38] = (x[11] & x[20]);
  assign t[39] = (x[8] & x[22]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[11] & x[24]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind111(x, y);
 input [25:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[24] | t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[25] | t[18]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[27]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[30]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = t[32] ^ x[5];
  assign t[24] = t[33] ^ x[10];
  assign t[25] = t[34] ^ x[13];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[17];
  assign t[28] = t[37] ^ x[19];
  assign t[29] = t[38] ^ x[21];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[23];
  assign t[31] = t[40] ^ x[25];
  assign t[32] = (x[3] & x[4]);
  assign t[33] = (x[8] & x[9]);
  assign t[34] = (x[11] & x[12]);
  assign t[35] = (x[8] & x[14]);
  assign t[36] = (x[8] & x[16]);
  assign t[37] = (x[11] & x[18]);
  assign t[38] = (x[11] & x[20]);
  assign t[39] = (x[8] & x[22]);
  assign t[3] = ~x[2] & t[23];
  assign t[40] = (x[11] & x[24]);
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[6] : t[7];
  assign t[6] = x[2] ? x[7] : t[8];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13] | t[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind112(x, y);
 input [21:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25] & t[18]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[26] & t[19]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[27] & t[20]);
  assign t[19] = ~(t[22]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[24]);
  assign t[21] = t[28] ^ x[7];
  assign t[22] = t[29] ^ x[10];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[17];
  assign t[26] = t[33] ^ x[19];
  assign t[27] = t[34] ^ x[21];
  assign t[28] = (x[5] & x[6]);
  assign t[29] = (x[8] & x[9]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[8] & x[11]);
  assign t[31] = (x[13] & x[14]);
  assign t[32] = (x[13] & x[16]);
  assign t[33] = (x[8] & x[18]);
  assign t[34] = (x[13] & x[20]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[21];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind113(x, y);
 input [25:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[26]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[29] & t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[31] & t[30]);
  assign t[24] = ~(t[33]);
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[15];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[19];
  assign t[31] = t[40] ^ x[21];
  assign t[32] = t[41] ^ x[23];
  assign t[33] = t[42] ^ x[25];
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[8] & x[9]);
  assign t[36] = (x[11] & x[12]);
  assign t[37] = (x[8] & x[14]);
  assign t[38] = (x[8] & x[16]);
  assign t[39] = (x[11] & x[18]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[11] & x[20]);
  assign t[41] = (x[8] & x[22]);
  assign t[42] = (x[11] & x[24]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind114(x, y);
 input [25:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~t[2];
  assign t[10] = t[15] | t[22];
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = t[18] | t[23];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[19] | t[13]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[20] | t[16]);
  assign t[19] = ~(t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[29]);
  assign t[21] = t[30] ^ x[5];
  assign t[22] = t[31] ^ x[10];
  assign t[23] = t[32] ^ x[13];
  assign t[24] = t[33] ^ x[15];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[19];
  assign t[27] = t[36] ^ x[21];
  assign t[28] = t[37] ^ x[23];
  assign t[29] = t[38] ^ x[25];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[3] & x[4]);
  assign t[31] = (x[8] & x[9]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[8] & x[14]);
  assign t[34] = (x[8] & x[16]);
  assign t[35] = (x[11] & x[18]);
  assign t[36] = (x[11] & x[20]);
  assign t[37] = (x[8] & x[22]);
  assign t[38] = (x[11] & x[24]);
  assign t[3] = ~x[2] & t[21];
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[6] : t[7];
  assign t[6] = x[2] ? x[7] : t[8];
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind115(x, y);
 input [28:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[28] | t[19]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[30] | t[22]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[20];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[24];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[28];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[8] & x[17]);
  assign t[42] = (x[8] & x[19]);
  assign t[43] = (x[14] & x[21]);
  assign t[44] = (x[14] & x[23]);
  assign t[45] = (x[8] & x[25]);
  assign t[46] = (x[14] & x[27]);
  assign t[4] = ~(~x[2] & ~t[27]);
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind116(x, y);
 input [24:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[24] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[27] & t[19]);
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[29] & t[21]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[30] & t[22]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[27]);
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[10];
  assign t[25] = t[33] ^ x[12];
  assign t[26] = t[34] ^ x[15];
  assign t[27] = t[35] ^ x[18];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[22];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[38] ^ x[24];
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[8] & x[9]);
  assign t[33] = (x[8] & x[11]);
  assign t[34] = (x[13] & x[14]);
  assign t[35] = (x[16] & x[17]);
  assign t[36] = (x[16] & x[19]);
  assign t[37] = (x[8] & x[21]);
  assign t[38] = (x[16] & x[23]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[4] = ~x[2] & t[23];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind117(x, y);
 input [28:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[28]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[30]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[32] & t[31]);
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[34] & t[33]);
  assign t[26] = ~(t[36]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[20];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[24];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[28];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[8] & x[17]);
  assign t[42] = (x[8] & x[19]);
  assign t[43] = (x[14] & x[21]);
  assign t[44] = (x[14] & x[23]);
  assign t[45] = (x[8] & x[25]);
  assign t[46] = (x[14] & x[27]);
  assign t[4] = ~x[2] & t[27];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind118(x, y);
 input [25:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = t[18] | t[24];
  assign t[13] = ~x[2] & t[25];
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = t[21] | t[26];
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[22] | t[16]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[23] | t[19]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[32]);
  assign t[24] = t[33] ^ x[7];
  assign t[25] = t[34] ^ x[10];
  assign t[26] = t[35] ^ x[13];
  assign t[27] = t[36] ^ x[15];
  assign t[28] = t[37] ^ x[17];
  assign t[29] = t[38] ^ x[19];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[21];
  assign t[31] = t[40] ^ x[23];
  assign t[32] = t[41] ^ x[25];
  assign t[33] = (x[5] & x[6]);
  assign t[34] = (x[8] & x[9]);
  assign t[35] = (x[11] & x[12]);
  assign t[36] = (x[5] & x[14]);
  assign t[37] = (x[5] & x[16]);
  assign t[38] = (x[11] & x[18]);
  assign t[39] = (x[11] & x[20]);
  assign t[3] = t[6] ? x[1] : x[0];
  assign t[40] = (x[5] & x[22]);
  assign t[41] = (x[11] & x[24]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind119(x, y);
 input [28:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[28] | t[19]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[30] | t[22]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[20];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[24];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[28];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[8] & x[17]);
  assign t[42] = (x[8] & x[19]);
  assign t[43] = (x[14] & x[21]);
  assign t[44] = (x[14] & x[23]);
  assign t[45] = (x[8] & x[25]);
  assign t[46] = (x[14] & x[27]);
  assign t[4] = ~(~x[2] & ~t[27]);
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind120(x, y);
 input [24:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[24] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[27] & t[19]);
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[29] & t[21]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[30] & t[22]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[27]);
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[10];
  assign t[25] = t[33] ^ x[12];
  assign t[26] = t[34] ^ x[15];
  assign t[27] = t[35] ^ x[18];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[22];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[38] ^ x[24];
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[8] & x[9]);
  assign t[33] = (x[8] & x[11]);
  assign t[34] = (x[13] & x[14]);
  assign t[35] = (x[16] & x[17]);
  assign t[36] = (x[16] & x[19]);
  assign t[37] = (x[8] & x[21]);
  assign t[38] = (x[16] & x[23]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[4] = ~x[2] & t[23];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind121(x, y);
 input [28:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[28]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[30]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[32] & t[31]);
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[34] & t[33]);
  assign t[26] = ~(t[36]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[20];
  assign t[33] = t[43] ^ x[22];
  assign t[34] = t[44] ^ x[24];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[28];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[8] & x[17]);
  assign t[42] = (x[8] & x[19]);
  assign t[43] = (x[14] & x[21]);
  assign t[44] = (x[14] & x[23]);
  assign t[45] = (x[8] & x[25]);
  assign t[46] = (x[14] & x[27]);
  assign t[4] = ~x[2] & t[27];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind122(x, y);
 input [28:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[26];
  assign t[14] = ~x[2] & t[27];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = t[22] | t[28];
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[23] | t[17]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[24] | t[20]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34]);
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[16];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[20];
  assign t[31] = t[41] ^ x[22];
  assign t[32] = t[42] ^ x[24];
  assign t[33] = t[43] ^ x[26];
  assign t[34] = t[44] ^ x[28];
  assign t[35] = (x[3] & x[4]);
  assign t[36] = (x[8] & x[9]);
  assign t[37] = (x[11] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[8] & x[17]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[8] & x[19]);
  assign t[41] = (x[14] & x[21]);
  assign t[42] = (x[14] & x[23]);
  assign t[43] = (x[8] & x[25]);
  assign t[44] = (x[14] & x[27]);
  assign t[4] = ~x[2] & t[25];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind123(x, y);
 input [35:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[19];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[21];
  assign t[41] = t[54] ^ x[23];
  assign t[42] = t[55] ^ x[25];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[29];
  assign t[45] = t[58] ^ x[31];
  assign t[46] = t[59] ^ x[33];
  assign t[47] = t[60] ^ x[35];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[9] & x[18]);
  assign t[53] = (x[9] & x[20]);
  assign t[54] = (x[12] & x[22]);
  assign t[55] = (x[12] & x[24]);
  assign t[56] = (x[15] & x[26]);
  assign t[57] = (x[15] & x[28]);
  assign t[58] = (x[9] & x[30]);
  assign t[59] = (x[12] & x[32]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[15] & x[34]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind124(x, y);
 input [29:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[13];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[18];
  assign t[34] = t[44] ^ x[21];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = t[46] ^ x[25];
  assign t[37] = t[47] ^ x[27];
  assign t[38] = t[48] ^ x[29];
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[9] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[14] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[19] & x[22]);
  assign t[46] = (x[9] & x[24]);
  assign t[47] = (x[14] & x[26]);
  assign t[48] = (x[19] & x[28]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind125(x, y);
 input [35:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = ~(t[22] & t[36]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[37]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] & t[34]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[44] & t[43]);
  assign t[34] = ~(t[47]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[19];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[21];
  assign t[41] = t[54] ^ x[23];
  assign t[42] = t[55] ^ x[25];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[29];
  assign t[45] = t[58] ^ x[31];
  assign t[46] = t[59] ^ x[33];
  assign t[47] = t[60] ^ x[35];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[9] & x[18]);
  assign t[53] = (x[9] & x[20]);
  assign t[54] = (x[12] & x[22]);
  assign t[55] = (x[12] & x[24]);
  assign t[56] = (x[15] & x[26]);
  assign t[57] = (x[15] & x[28]);
  assign t[58] = (x[9] & x[30]);
  assign t[59] = (x[12] & x[32]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[15] & x[34]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind126(x, y);
 input [35:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[8];
  assign t[33] = t[46] ^ x[11];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[19];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[23];
  assign t[39] = t[52] ^ x[25];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[27];
  assign t[41] = t[54] ^ x[29];
  assign t[42] = t[55] ^ x[31];
  assign t[43] = t[56] ^ x[33];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = (x[6] & x[7]);
  assign t[46] = (x[9] & x[10]);
  assign t[47] = (x[12] & x[13]);
  assign t[48] = (x[15] & x[16]);
  assign t[49] = (x[9] & x[18]);
  assign t[4] = t[7];
  assign t[50] = (x[9] & x[20]);
  assign t[51] = (x[12] & x[22]);
  assign t[52] = (x[12] & x[24]);
  assign t[53] = (x[15] & x[26]);
  assign t[54] = (x[15] & x[28]);
  assign t[55] = (x[9] & x[30]);
  assign t[56] = (x[12] & x[32]);
  assign t[57] = (x[15] & x[34]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind127(x, y);
 input [35:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[19];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[21];
  assign t[41] = t[54] ^ x[23];
  assign t[42] = t[55] ^ x[25];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[29];
  assign t[45] = t[58] ^ x[31];
  assign t[46] = t[59] ^ x[33];
  assign t[47] = t[60] ^ x[35];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[9] & x[18]);
  assign t[53] = (x[9] & x[20]);
  assign t[54] = (x[12] & x[22]);
  assign t[55] = (x[12] & x[24]);
  assign t[56] = (x[15] & x[26]);
  assign t[57] = (x[15] & x[28]);
  assign t[58] = (x[9] & x[30]);
  assign t[59] = (x[12] & x[32]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[15] & x[34]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind128(x, y);
 input [29:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[28] & t[18]);
  assign t[13] = ~(t[29] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[34] & t[24]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[35] & t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = ~(t[36] & t[26]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[30]);
  assign t[26] = ~(t[32]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[11];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[21];
  assign t[33] = t[43] ^ x[23];
  assign t[34] = t[44] ^ x[25];
  assign t[35] = t[45] ^ x[27];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[9] & x[10]);
  assign t[39] = (x[9] & x[12]);
  assign t[3] = ~x[2] & t[27];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[14] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[19] & x[22]);
  assign t[44] = (x[9] & x[24]);
  assign t[45] = (x[14] & x[26]);
  assign t[46] = (x[19] & x[28]);
  assign t[4] = t[6];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind129(x, y);
 input [35:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = ~(t[20] & t[34]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = ~(t[23] & t[35]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26] & t[36]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] & t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] & t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[38] & t[37]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[45]);
  assign t[33] = t[46] ^ x[5];
  assign t[34] = t[47] ^ x[11];
  assign t[35] = t[48] ^ x[14];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[19];
  assign t[38] = t[51] ^ x[21];
  assign t[39] = t[52] ^ x[23];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[25];
  assign t[41] = t[54] ^ x[27];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[31];
  assign t[44] = t[57] ^ x[33];
  assign t[45] = t[58] ^ x[35];
  assign t[46] = (x[3] & x[4]);
  assign t[47] = (x[9] & x[10]);
  assign t[48] = (x[12] & x[13]);
  assign t[49] = (x[15] & x[16]);
  assign t[4] = t[6];
  assign t[50] = (x[9] & x[18]);
  assign t[51] = (x[9] & x[20]);
  assign t[52] = (x[12] & x[22]);
  assign t[53] = (x[12] & x[24]);
  assign t[54] = (x[15] & x[26]);
  assign t[55] = (x[15] & x[28]);
  assign t[56] = (x[9] & x[30]);
  assign t[57] = (x[12] & x[32]);
  assign t[58] = (x[15] & x[34]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind130(x, y);
 input [35:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[8];
  assign t[33] = t[46] ^ x[11];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[19];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[23];
  assign t[39] = t[52] ^ x[25];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[27];
  assign t[41] = t[54] ^ x[29];
  assign t[42] = t[55] ^ x[31];
  assign t[43] = t[56] ^ x[33];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = (x[6] & x[7]);
  assign t[46] = (x[9] & x[10]);
  assign t[47] = (x[12] & x[13]);
  assign t[48] = (x[15] & x[16]);
  assign t[49] = (x[9] & x[18]);
  assign t[4] = t[7];
  assign t[50] = (x[9] & x[20]);
  assign t[51] = (x[12] & x[22]);
  assign t[52] = (x[12] & x[24]);
  assign t[53] = (x[15] & x[26]);
  assign t[54] = (x[15] & x[28]);
  assign t[55] = (x[9] & x[30]);
  assign t[56] = (x[12] & x[32]);
  assign t[57] = (x[15] & x[34]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind131(x, y);
 input [35:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[18] | t[19]);
  assign t[13] = ~(t[34] | t[20]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[15] = ~(t[35] | t[23]);
  assign t[16] = ~(t[24] | t[25]);
  assign t[17] = ~(t[36] | t[26]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] | t[32]);
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[37] | t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = t[46] ^ x[5];
  assign t[34] = t[47] ^ x[11];
  assign t[35] = t[48] ^ x[14];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[19];
  assign t[38] = t[51] ^ x[21];
  assign t[39] = t[52] ^ x[23];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[25];
  assign t[41] = t[54] ^ x[27];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[31];
  assign t[44] = t[57] ^ x[33];
  assign t[45] = t[58] ^ x[35];
  assign t[46] = (x[3] & x[4]);
  assign t[47] = (x[9] & x[10]);
  assign t[48] = (x[12] & x[13]);
  assign t[49] = (x[15] & x[16]);
  assign t[4] = t[6];
  assign t[50] = (x[9] & x[18]);
  assign t[51] = (x[9] & x[20]);
  assign t[52] = (x[12] & x[22]);
  assign t[53] = (x[12] & x[24]);
  assign t[54] = (x[15] & x[26]);
  assign t[55] = (x[15] & x[28]);
  assign t[56] = (x[9] & x[30]);
  assign t[57] = (x[12] & x[32]);
  assign t[58] = (x[15] & x[34]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind132(x, y);
 input [29:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[13];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[18];
  assign t[34] = t[44] ^ x[21];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = t[46] ^ x[25];
  assign t[37] = t[47] ^ x[27];
  assign t[38] = t[48] ^ x[29];
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[9] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[14] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[19] & x[22]);
  assign t[46] = (x[9] & x[24]);
  assign t[47] = (x[14] & x[26]);
  assign t[48] = (x[19] & x[28]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind133(x, y);
 input [35:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = ~(t[22] & t[36]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[37]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] & t[34]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[44] & t[43]);
  assign t[34] = ~(t[47]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[19];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[21];
  assign t[41] = t[54] ^ x[23];
  assign t[42] = t[55] ^ x[25];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[29];
  assign t[45] = t[58] ^ x[31];
  assign t[46] = t[59] ^ x[33];
  assign t[47] = t[60] ^ x[35];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[9] & x[18]);
  assign t[53] = (x[9] & x[20]);
  assign t[54] = (x[12] & x[22]);
  assign t[55] = (x[12] & x[24]);
  assign t[56] = (x[15] & x[26]);
  assign t[57] = (x[15] & x[28]);
  assign t[58] = (x[9] & x[30]);
  assign t[59] = (x[12] & x[32]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[15] & x[34]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind134(x, y);
 input [35:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = t[20] | t[31];
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = t[23] | t[32];
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = t[26] | t[33];
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[35]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] | t[18]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[28] | t[21]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[29] | t[24]);
  assign t[27] = ~(t[40]);
  assign t[28] = ~(t[41]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ x[5];
  assign t[31] = t[44] ^ x[11];
  assign t[32] = t[45] ^ x[14];
  assign t[33] = t[46] ^ x[17];
  assign t[34] = t[47] ^ x[19];
  assign t[35] = t[48] ^ x[21];
  assign t[36] = t[49] ^ x[23];
  assign t[37] = t[50] ^ x[25];
  assign t[38] = t[51] ^ x[27];
  assign t[39] = t[52] ^ x[29];
  assign t[3] = ~x[2] & t[30];
  assign t[40] = t[53] ^ x[31];
  assign t[41] = t[54] ^ x[33];
  assign t[42] = t[55] ^ x[35];
  assign t[43] = (x[3] & x[4]);
  assign t[44] = (x[9] & x[10]);
  assign t[45] = (x[12] & x[13]);
  assign t[46] = (x[15] & x[16]);
  assign t[47] = (x[9] & x[18]);
  assign t[48] = (x[9] & x[20]);
  assign t[49] = (x[12] & x[22]);
  assign t[4] = t[6];
  assign t[50] = (x[12] & x[24]);
  assign t[51] = (x[15] & x[26]);
  assign t[52] = (x[15] & x[28]);
  assign t[53] = (x[9] & x[30]);
  assign t[54] = (x[12] & x[32]);
  assign t[55] = (x[15] & x[34]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind135(x, y);
 input [35:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[19];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[21];
  assign t[41] = t[54] ^ x[23];
  assign t[42] = t[55] ^ x[25];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[29];
  assign t[45] = t[58] ^ x[31];
  assign t[46] = t[59] ^ x[33];
  assign t[47] = t[60] ^ x[35];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[9] & x[18]);
  assign t[53] = (x[9] & x[20]);
  assign t[54] = (x[12] & x[22]);
  assign t[55] = (x[12] & x[24]);
  assign t[56] = (x[15] & x[26]);
  assign t[57] = (x[15] & x[28]);
  assign t[58] = (x[9] & x[30]);
  assign t[59] = (x[12] & x[32]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[15] & x[34]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind136(x, y);
 input [29:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[13];
  assign t[32] = t[42] ^ x[16];
  assign t[33] = t[43] ^ x[18];
  assign t[34] = t[44] ^ x[21];
  assign t[35] = t[45] ^ x[23];
  assign t[36] = t[46] ^ x[25];
  assign t[37] = t[47] ^ x[27];
  assign t[38] = t[48] ^ x[29];
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[9] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[14] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[19] & x[22]);
  assign t[46] = (x[9] & x[24]);
  assign t[47] = (x[14] & x[26]);
  assign t[48] = (x[19] & x[28]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind137(x, y);
 input [35:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = ~(t[20] & t[34]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = ~(t[23] & t[35]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26] & t[36]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] & t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] & t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[38] & t[37]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[45]);
  assign t[33] = t[46] ^ x[5];
  assign t[34] = t[47] ^ x[11];
  assign t[35] = t[48] ^ x[14];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[19];
  assign t[38] = t[51] ^ x[21];
  assign t[39] = t[52] ^ x[23];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[25];
  assign t[41] = t[54] ^ x[27];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[31];
  assign t[44] = t[57] ^ x[33];
  assign t[45] = t[58] ^ x[35];
  assign t[46] = (x[3] & x[4]);
  assign t[47] = (x[9] & x[10]);
  assign t[48] = (x[12] & x[13]);
  assign t[49] = (x[15] & x[16]);
  assign t[4] = t[6];
  assign t[50] = (x[9] & x[18]);
  assign t[51] = (x[9] & x[20]);
  assign t[52] = (x[12] & x[22]);
  assign t[53] = (x[12] & x[24]);
  assign t[54] = (x[15] & x[26]);
  assign t[55] = (x[15] & x[28]);
  assign t[56] = (x[9] & x[30]);
  assign t[57] = (x[12] & x[32]);
  assign t[58] = (x[15] & x[34]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind138(x, y);
 input [35:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[8];
  assign t[33] = t[46] ^ x[11];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[19];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[23];
  assign t[39] = t[52] ^ x[25];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[27];
  assign t[41] = t[54] ^ x[29];
  assign t[42] = t[55] ^ x[31];
  assign t[43] = t[56] ^ x[33];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = (x[6] & x[7]);
  assign t[46] = (x[9] & x[10]);
  assign t[47] = (x[12] & x[13]);
  assign t[48] = (x[15] & x[16]);
  assign t[49] = (x[9] & x[18]);
  assign t[4] = t[7];
  assign t[50] = (x[9] & x[20]);
  assign t[51] = (x[12] & x[22]);
  assign t[52] = (x[12] & x[24]);
  assign t[53] = (x[15] & x[26]);
  assign t[54] = (x[15] & x[28]);
  assign t[55] = (x[9] & x[30]);
  assign t[56] = (x[12] & x[32]);
  assign t[57] = (x[15] & x[34]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1_ind(x, y);
 input [366:0] x;
 output [138:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[171], x[170], x[169], x[147]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[171], x[170], x[169], x[174], x[173], x[172], x[147]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[159], x[158], x[157], x[147]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[156], x[155], x[154], x[147]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[153], x[152], x[151], x[159], x[158], x[157], x[147]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[165], x[164], x[163], x[147]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[168], x[167], x[166], x[147]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[150], x[149], x[148], x[147]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[165], x[164], x[163], x[162], x[161], x[160], x[147]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[140], x[139], x[146], x[145], x[144], x[143], x[142], x[141], x[138], x[171], x[170], x[169], x[177], x[147], x[176], x[175]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[146], x[145], x[171], x[170], x[169], x[140], x[139], x[144], x[143], x[138], x[180], x[147], x[179], x[178]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[144], x[143], x[140], x[139], x[146], x[145], x[142], x[141], x[138], x[171], x[170], x[169], x[183], x[147], x[182], x[181]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[144], x[143], x[140], x[139], x[146], x[145], x[171], x[170], x[169], x[142], x[141], x[138], x[186], x[147], x[185], x[184]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[113], x[112], x[119], x[118], x[117], x[116], x[171], x[170], x[169], x[115], x[114], x[111], x[189], x[147], x[188], x[187]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[119], x[118], x[171], x[170], x[169], x[113], x[112], x[117], x[116], x[111], x[192], x[147], x[191], x[190]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[117], x[116], x[113], x[112], x[119], x[118], x[171], x[170], x[169], x[115], x[114], x[111], x[195], x[147], x[194], x[193]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[117], x[116], x[113], x[112], x[119], x[118], x[171], x[170], x[169], x[115], x[114], x[111], x[198], x[147], x[197], x[196]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[122], x[121], x[128], x[127], x[126], x[125], x[171], x[170], x[169], x[124], x[123], x[120], x[201], x[147], x[200], x[199]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[128], x[127], x[171], x[170], x[169], x[122], x[121], x[126], x[125], x[120], x[204], x[147], x[203], x[202]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[126], x[125], x[122], x[121], x[128], x[127], x[171], x[170], x[169], x[124], x[123], x[120], x[207], x[147], x[206], x[205]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[126], x[125], x[122], x[121], x[128], x[127], x[171], x[170], x[169], x[124], x[123], x[120], x[210], x[147], x[209], x[208]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[131], x[130], x[137], x[136], x[135], x[134], x[171], x[170], x[169], x[133], x[132], x[129], x[213], x[147], x[212], x[211]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[137], x[136], x[171], x[170], x[169], x[131], x[130], x[135], x[134], x[129], x[216], x[147], x[215], x[214]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[135], x[134], x[131], x[130], x[137], x[136], x[171], x[170], x[169], x[133], x[132], x[129], x[219], x[147], x[218], x[217]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[135], x[134], x[131], x[130], x[137], x[136], x[171], x[170], x[169], x[133], x[132], x[129], x[222], x[147], x[221], x[220]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[77], x[76], x[83], x[82], x[81], x[80], x[171], x[170], x[169], x[79], x[78], x[75], x[225], x[147], x[224], x[223]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[83], x[82], x[171], x[170], x[169], x[77], x[76], x[81], x[80], x[75], x[228], x[147], x[227], x[226]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[81], x[80], x[77], x[76], x[83], x[82], x[171], x[170], x[169], x[79], x[78], x[75], x[231], x[147], x[230], x[229]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[81], x[80], x[77], x[76], x[83], x[82], x[171], x[170], x[169], x[79], x[78], x[75], x[234], x[147], x[233], x[232]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[104], x[103], x[110], x[109], x[108], x[107], x[171], x[170], x[169], x[106], x[105], x[102], x[237], x[147], x[236], x[235]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[110], x[109], x[171], x[170], x[169], x[104], x[103], x[108], x[107], x[102], x[240], x[147], x[239], x[238]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[108], x[107], x[104], x[103], x[110], x[109], x[106], x[105], x[102], x[171], x[170], x[169], x[243], x[147], x[242], x[241]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[108], x[107], x[104], x[103], x[110], x[109], x[106], x[105], x[102], x[171], x[170], x[169], x[246], x[147], x[245], x[244]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[95], x[94], x[101], x[100], x[99], x[98], x[97], x[96], x[93], x[171], x[170], x[169], x[249], x[147], x[248], x[247]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[101], x[100], x[95], x[94], x[99], x[98], x[93], x[171], x[170], x[169], x[252], x[147], x[251], x[250]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[99], x[98], x[95], x[94], x[101], x[100], x[97], x[96], x[93], x[171], x[170], x[169], x[255], x[147], x[254], x[253]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[99], x[98], x[95], x[94], x[101], x[100], x[97], x[96], x[93], x[171], x[170], x[169], x[258], x[147], x[257], x[256]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[86], x[85], x[92], x[91], x[90], x[89], x[171], x[170], x[169], x[88], x[87], x[84], x[261], x[147], x[260], x[259]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[92], x[91], x[171], x[170], x[169], x[86], x[85], x[90], x[89], x[84], x[264], x[147], x[263], x[262]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[90], x[89], x[86], x[85], x[92], x[91], x[171], x[170], x[169], x[88], x[87], x[84], x[267], x[147], x[266], x[265]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[90], x[89], x[86], x[85], x[92], x[91], x[171], x[170], x[169], x[88], x[87], x[84], x[270], x[147], x[269], x[268]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[41], x[40], x[140], x[139], x[47], x[46], x[45], x[44], x[146], x[145], x[144], x[143], x[43], x[42], x[39], x[142], x[141], x[138], x[171], x[170], x[169], x[273], x[177], x[147], x[272], x[271]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[47], x[46], x[146], x[145], x[41], x[40], x[45], x[44], x[39], x[140], x[139], x[144], x[143], x[138], x[276], x[180], x[171], x[170], x[169], x[147], x[275], x[274]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[45], x[44], x[144], x[143], x[41], x[40], x[47], x[46], x[140], x[139], x[146], x[145], x[43], x[42], x[39], x[142], x[141], x[138], x[171], x[170], x[169], x[279], x[183], x[147], x[278], x[277]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[45], x[44], x[144], x[143], x[41], x[40], x[47], x[46], x[140], x[139], x[146], x[145], x[43], x[42], x[39], x[142], x[141], x[138], x[171], x[170], x[169], x[282], x[186], x[147], x[281], x[280]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[68], x[67], x[113], x[112], x[74], x[73], x[72], x[71], x[119], x[118], x[117], x[116], x[70], x[69], x[66], x[115], x[114], x[111], x[285], x[189], x[171], x[170], x[169], x[147], x[284], x[283]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[74], x[73], x[119], x[118], x[68], x[67], x[72], x[71], x[66], x[113], x[112], x[117], x[116], x[111], x[171], x[170], x[169], x[288], x[192], x[147], x[287], x[286]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[72], x[71], x[117], x[116], x[68], x[67], x[74], x[73], x[113], x[112], x[119], x[118], x[70], x[69], x[66], x[115], x[114], x[111], x[171], x[170], x[169], x[291], x[195], x[147], x[290], x[289]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[72], x[71], x[117], x[116], x[68], x[67], x[74], x[73], x[113], x[112], x[119], x[118], x[70], x[69], x[66], x[115], x[114], x[111], x[294], x[198], x[171], x[170], x[169], x[147], x[293], x[292]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[59], x[58], x[122], x[121], x[65], x[64], x[63], x[62], x[128], x[127], x[126], x[125], x[61], x[60], x[57], x[171], x[170], x[169], x[124], x[123], x[120], x[297], x[201], x[153], x[152], x[151], x[147], x[296], x[295]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[65], x[64], x[128], x[127], x[59], x[58], x[63], x[62], x[57], x[171], x[170], x[169], x[122], x[121], x[126], x[125], x[120], x[300], x[204], x[159], x[158], x[157], x[147], x[299], x[298]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[63], x[62], x[126], x[125], x[59], x[58], x[65], x[64], x[122], x[121], x[128], x[127], x[61], x[60], x[57], x[171], x[170], x[169], x[124], x[123], x[120], x[303], x[207], x[156], x[155], x[154], x[147], x[302], x[301]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[63], x[62], x[126], x[125], x[59], x[58], x[65], x[64], x[122], x[121], x[128], x[127], x[61], x[60], x[57], x[171], x[170], x[169], x[124], x[123], x[120], x[306], x[210], x[147], x[305], x[304]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[50], x[49], x[131], x[130], x[56], x[55], x[54], x[53], x[137], x[136], x[135], x[134], x[52], x[51], x[48], x[171], x[170], x[169], x[133], x[132], x[129], x[309], x[213], x[162], x[161], x[160], x[147], x[308], x[307]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[56], x[55], x[137], x[136], x[50], x[49], x[54], x[53], x[48], x[171], x[170], x[169], x[131], x[130], x[135], x[134], x[129], x[312], x[216], x[165], x[164], x[163], x[147], x[311], x[310]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[54], x[53], x[135], x[134], x[50], x[49], x[56], x[55], x[131], x[130], x[137], x[136], x[52], x[51], x[48], x[171], x[170], x[169], x[133], x[132], x[129], x[315], x[219], x[168], x[167], x[166], x[147], x[314], x[313]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[54], x[53], x[135], x[134], x[50], x[49], x[56], x[55], x[131], x[130], x[137], x[136], x[52], x[51], x[48], x[171], x[170], x[169], x[133], x[132], x[129], x[318], x[222], x[150], x[149], x[148], x[147], x[317], x[316]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[140], x[139], x[77], x[76], x[14], x[13], x[146], x[145], x[144], x[143], x[83], x[82], x[81], x[80], x[20], x[19], x[18], x[17], x[142], x[141], x[138], x[79], x[78], x[75], x[16], x[15], x[12], x[171], x[170], x[169], x[177], x[225], x[321], x[147], x[320], x[319]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[146], x[145], x[83], x[82], x[20], x[19], x[140], x[139], x[144], x[143], x[138], x[77], x[76], x[81], x[80], x[75], x[14], x[13], x[18], x[17], x[12], x[171], x[170], x[169], x[180], x[228], x[324], x[147], x[323], x[322]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[144], x[143], x[81], x[80], x[18], x[17], x[140], x[139], x[146], x[145], x[77], x[76], x[83], x[82], x[14], x[13], x[20], x[19], x[142], x[141], x[138], x[79], x[78], x[75], x[16], x[15], x[12], x[171], x[170], x[169], x[183], x[231], x[327], x[147], x[326], x[325]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[144], x[143], x[81], x[80], x[18], x[17], x[140], x[139], x[146], x[145], x[77], x[76], x[83], x[82], x[14], x[13], x[20], x[19], x[142], x[141], x[138], x[79], x[78], x[75], x[16], x[15], x[12], x[171], x[170], x[169], x[186], x[234], x[330], x[147], x[329], x[328]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[113], x[112], x[104], x[103], x[23], x[22], x[119], x[118], x[117], x[116], x[110], x[109], x[108], x[107], x[29], x[28], x[27], x[26], x[115], x[114], x[111], x[106], x[105], x[102], x[25], x[24], x[21], x[171], x[170], x[169], x[189], x[237], x[333], x[147], x[332], x[331]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[119], x[118], x[110], x[109], x[29], x[28], x[113], x[112], x[117], x[116], x[111], x[104], x[103], x[108], x[107], x[102], x[23], x[22], x[27], x[26], x[21], x[192], x[240], x[336], x[171], x[170], x[169], x[147], x[335], x[334]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[117], x[116], x[108], x[107], x[27], x[26], x[113], x[112], x[119], x[118], x[104], x[103], x[110], x[109], x[23], x[22], x[29], x[28], x[115], x[114], x[111], x[106], x[105], x[102], x[25], x[24], x[21], x[195], x[243], x[339], x[171], x[170], x[169], x[147], x[338], x[337]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[117], x[116], x[108], x[107], x[27], x[26], x[113], x[112], x[119], x[118], x[104], x[103], x[110], x[109], x[23], x[22], x[29], x[28], x[115], x[114], x[111], x[106], x[105], x[102], x[25], x[24], x[21], x[171], x[170], x[169], x[198], x[246], x[342], x[147], x[341], x[340]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[122], x[121], x[95], x[94], x[32], x[31], x[128], x[127], x[126], x[125], x[101], x[100], x[99], x[98], x[38], x[37], x[36], x[35], x[124], x[123], x[120], x[97], x[96], x[93], x[34], x[33], x[30], x[201], x[249], x[345], x[171], x[170], x[169], x[147], x[344], x[343]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[128], x[127], x[101], x[100], x[38], x[37], x[122], x[121], x[126], x[125], x[120], x[95], x[94], x[99], x[98], x[93], x[32], x[31], x[36], x[35], x[30], x[171], x[170], x[169], x[204], x[252], x[348], x[147], x[347], x[346]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[126], x[125], x[99], x[98], x[36], x[35], x[122], x[121], x[128], x[127], x[95], x[94], x[101], x[100], x[32], x[31], x[38], x[37], x[124], x[123], x[120], x[97], x[96], x[93], x[34], x[33], x[30], x[171], x[170], x[169], x[207], x[255], x[351], x[147], x[350], x[349]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[126], x[125], x[99], x[98], x[36], x[35], x[122], x[121], x[128], x[127], x[95], x[94], x[101], x[100], x[32], x[31], x[38], x[37], x[124], x[123], x[120], x[97], x[96], x[93], x[34], x[33], x[30], x[210], x[258], x[354], x[171], x[170], x[169], x[147], x[353], x[352]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[131], x[130], x[86], x[85], x[5], x[4], x[137], x[136], x[135], x[134], x[92], x[91], x[90], x[89], x[11], x[10], x[9], x[8], x[133], x[132], x[129], x[88], x[87], x[84], x[7], x[6], x[3], x[171], x[170], x[169], x[213], x[261], x[357], x[147], x[356], x[355]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[137], x[136], x[92], x[91], x[11], x[10], x[131], x[130], x[135], x[134], x[129], x[86], x[85], x[90], x[89], x[84], x[5], x[4], x[9], x[8], x[3], x[171], x[170], x[169], x[216], x[264], x[360], x[147], x[359], x[358]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[135], x[134], x[90], x[89], x[9], x[8], x[131], x[130], x[137], x[136], x[86], x[85], x[92], x[91], x[5], x[4], x[11], x[10], x[133], x[132], x[129], x[88], x[87], x[84], x[7], x[6], x[3], x[219], x[267], x[363], x[171], x[170], x[169], x[147], x[362], x[361]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[135], x[134], x[90], x[89], x[9], x[8], x[131], x[130], x[137], x[136], x[86], x[85], x[92], x[91], x[5], x[4], x[11], x[10], x[133], x[132], x[129], x[88], x[87], x[84], x[7], x[6], x[3], x[171], x[170], x[169], x[222], x[270], x[366], x[147], x[365], x[364]}), .y(y[138]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [21:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[11] = ~x[0] & t[18];
  assign t[12] = ~x[0] & t[19];
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[27] ^ x[3];
  assign t[21] = t[28] ^ x[6];
  assign t[22] = t[29] ^ x[9];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[18];
  assign t[26] = t[33] ^ x[21];
  assign t[27] = (~t[34] & t[35]);
  assign t[28] = (~t[36] & t[37]);
  assign t[29] = (~t[38] & t[39]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (~t[40] & t[41]);
  assign t[31] = (~t[42] & t[43]);
  assign t[32] = (~t[44] & t[45]);
  assign t[33] = (~t[46] & t[47]);
  assign t[34] = t[48] ^ x[2];
  assign t[35] = t[49] ^ x[3];
  assign t[36] = t[50] ^ x[5];
  assign t[37] = t[51] ^ x[6];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[11];
  assign t[41] = t[55] ^ x[12];
  assign t[42] = t[56] ^ x[14];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[18];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[51] = (x[4]);
  assign t[52] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[53] = (x[7]);
  assign t[54] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[10]);
  assign t[56] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[13]);
  assign t[58] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[16]);
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[19]);
  assign t[6] = ~x[0] & t[15];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [21:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[11] = ~x[0] & t[18];
  assign t[12] = ~x[0] & t[19];
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[27] ^ x[3];
  assign t[21] = t[28] ^ x[6];
  assign t[22] = t[29] ^ x[9];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[18];
  assign t[26] = t[33] ^ x[21];
  assign t[27] = (~t[34] & t[35]);
  assign t[28] = (~t[36] & t[37]);
  assign t[29] = (~t[38] & t[39]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (~t[40] & t[41]);
  assign t[31] = (~t[42] & t[43]);
  assign t[32] = (~t[44] & t[45]);
  assign t[33] = (~t[46] & t[47]);
  assign t[34] = t[48] ^ x[2];
  assign t[35] = t[49] ^ x[3];
  assign t[36] = t[50] ^ x[5];
  assign t[37] = t[51] ^ x[6];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[11];
  assign t[41] = t[55] ^ x[12];
  assign t[42] = t[56] ^ x[14];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[18];
  assign t[46] = t[60] ^ x[20];
  assign t[47] = t[61] ^ x[21];
  assign t[48] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[51] = (x[4]);
  assign t[52] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[53] = (x[7]);
  assign t[54] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[10]);
  assign t[56] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[13]);
  assign t[58] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[16]);
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[19]);
  assign t[6] = ~x[0] & t[15];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[14] = (x[1]);
  assign t[15] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[16] = (x[4]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (~t[9] & t[10]);
  assign t[8] = (~t[11] & t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[14] = (x[1]);
  assign t[15] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[16] = (x[4]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (~t[9] & t[10]);
  assign t[8] = (~t[11] & t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind31(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind34(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind36(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind37(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind38(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind39(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[14] = (x[1]);
  assign t[15] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[16] = (x[4]);
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = ~x[0] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (~t[9] & t[10]);
  assign t[8] = (~t[11] & t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind41(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind42(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind43(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind44(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[14] = (x[1]);
  assign t[15] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[16] = (x[4]);
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = ~x[0] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (~t[9] & t[10]);
  assign t[8] = (~t[11] & t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~x[0] & t[2];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[3];
  assign t[7] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind46(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind47(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind48(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind49(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~x[0] & t[2];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[2];
  assign t[6] = t[8] ^ x[3];
  assign t[7] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [6:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[1]);
  assign t[16] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[4]);
  assign t[1] = ~t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = ~x[0] & t[5];
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[6];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind51(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind52(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind53(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind54(x, y);
 input [6:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[1]);
  assign t[16] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[4]);
  assign t[1] = ~t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = ~x[0] & t[5];
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[6];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[42]);
  assign t[12] = ~(t[40] | t[41]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[17] ? x[17] : x[16];
  assign t[16] = x[2] ? x[18] : t[18];
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[4]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[9]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[8]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[9] & t[11]);
  assign t[29] = ~(t[30] & t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[8]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[17] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[6] | t[39];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[6];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~x[2] & t[38];
  assign t[50] = (~t[55] & t[57]);
  assign t[51] = (~t[55] & t[58]);
  assign t[52] = (~t[55] & t[59]);
  assign t[53] = t[60] ^ x[5];
  assign t[54] = t[61] ^ x[6];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[4]);
  assign t[62] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[63] = (x[8]);
  assign t[64] = (x[9]);
  assign t[65] = (x[10]);
  assign t[66] = (x[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[39] | t[10]);
  assign t[8] = ~(t[40]);
  assign t[9] = ~(t[41]);
  assign y = (t[0] & ~t[13] & ~t[23] & ~t[32]) | (~t[0] & t[13] & ~t[23] & ~t[32]) | (~t[0] & ~t[13] & t[23] & ~t[32]) | (~t[0] & ~t[13] & ~t[23] & t[32]) | (t[0] & t[13] & t[23] & ~t[32]) | (t[0] & t[13] & ~t[23] & t[32]) | (t[0] & ~t[13] & t[23] & t[32]) | (~t[0] & t[13] & t[23] & t[32]);
endmodule

module R2ind56(x, y);
 input [15:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[13];
  assign t[22] = t[27] ^ x[14];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = (~t[29] & t[34]);
  assign t[28] = (~t[29] & t[35]);
  assign t[29] = t[36] ^ x[8];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[9];
  assign t[31] = t[38] ^ x[11];
  assign t[32] = t[39] ^ x[12];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[14];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[37] = (x[5]);
  assign t[38] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[4]);
  assign t[42] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [15:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[4]);
  assign t[37] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[38] = (x[8]);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[9]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [15:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[4]);
  assign t[37] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[38] = (x[8]);
  assign t[39] = (x[9]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[40]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[42]);
  assign t[14] = ~(t[40] | t[41]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[17] : x[16];
  assign t[18] = x[2] ? x[18] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[11]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[4] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[7] | t[38];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[9];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[6]);
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = (~t[53] & t[58]);
  assign t[52] = (~t[53] & t[59]);
  assign t[53] = t[60] ^ x[8];
  assign t[54] = t[61] ^ x[9];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[61] = (x[5]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[6]);
  assign t[65] = (x[7]);
  assign t[66] = (x[4]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[38] | t[12]);
  assign t[9] = ~x[2] & t[39];
  assign y = (t[0] & ~t[15] & ~t[23] & ~t[32]) | (~t[0] & t[15] & ~t[23] & ~t[32]) | (~t[0] & ~t[15] & t[23] & ~t[32]) | (~t[0] & ~t[15] & ~t[23] & t[32]) | (t[0] & t[15] & t[23] & ~t[32]) | (t[0] & t[15] & ~t[23] & t[32]) | (t[0] & ~t[15] & t[23] & t[32]) | (~t[0] & t[15] & t[23] & t[32]);
endmodule

module R2ind61(x, y);
 input [15:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[13];
  assign t[22] = t[27] ^ x[14];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = (~t[29] & t[34]);
  assign t[28] = (~t[29] & t[35]);
  assign t[29] = t[36] ^ x[8];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[9];
  assign t[31] = t[38] ^ x[11];
  assign t[32] = t[39] ^ x[12];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[14];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[37] = (x[5]);
  assign t[38] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[4]);
  assign t[42] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[4]);
  assign t[43] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[6]);
  assign t[42] = (x[7]);
  assign t[43] = (x[4]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[40]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[42]);
  assign t[14] = ~(t[40] | t[41]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[17] : x[16];
  assign t[18] = x[2] ? x[18] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[11]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[4] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[7] | t[38];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[9];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[6]);
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = (~t[53] & t[58]);
  assign t[52] = (~t[53] & t[59]);
  assign t[53] = t[60] ^ x[8];
  assign t[54] = t[61] ^ x[9];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[61] = (x[5]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[6]);
  assign t[65] = (x[7]);
  assign t[66] = (x[4]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[38] | t[12]);
  assign t[9] = ~x[2] & t[39];
  assign y = (t[0] & ~t[15] & ~t[23] & ~t[32]) | (~t[0] & t[15] & ~t[23] & ~t[32]) | (~t[0] & ~t[15] & t[23] & ~t[32]) | (~t[0] & ~t[15] & ~t[23] & t[32]) | (t[0] & t[15] & t[23] & ~t[32]) | (t[0] & t[15] & ~t[23] & t[32]) | (t[0] & ~t[15] & t[23] & t[32]) | (~t[0] & t[15] & t[23] & t[32]);
endmodule

module R2ind66(x, y);
 input [15:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[13];
  assign t[22] = t[27] ^ x[14];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = (~t[29] & t[34]);
  assign t[28] = (~t[29] & t[35]);
  assign t[29] = t[36] ^ x[8];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[9];
  assign t[31] = t[38] ^ x[11];
  assign t[32] = t[39] ^ x[12];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[14];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[37] = (x[5]);
  assign t[38] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[4]);
  assign t[42] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[4]);
  assign t[43] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[6]);
  assign t[42] = (x[7]);
  assign t[43] = (x[4]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[40]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[42]);
  assign t[14] = ~(t[40] | t[41]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[17] : x[16];
  assign t[18] = x[2] ? x[18] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[11]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[4] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[7] | t[38];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[9];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[6]);
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = (~t[53] & t[58]);
  assign t[52] = (~t[53] & t[59]);
  assign t[53] = t[60] ^ x[8];
  assign t[54] = t[61] ^ x[9];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[61] = (x[5]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[6]);
  assign t[65] = (x[7]);
  assign t[66] = (x[4]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[38] | t[12]);
  assign t[9] = ~x[2] & t[39];
  assign y = (t[0] & ~t[15] & ~t[23] & ~t[32]) | (~t[0] & t[15] & ~t[23] & ~t[32]) | (~t[0] & ~t[15] & t[23] & ~t[32]) | (~t[0] & ~t[15] & ~t[23] & t[32]) | (t[0] & t[15] & t[23] & ~t[32]) | (t[0] & t[15] & ~t[23] & t[32]) | (t[0] & ~t[15] & t[23] & t[32]) | (~t[0] & t[15] & t[23] & t[32]);
endmodule

module R2ind71(x, y);
 input [15:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[13];
  assign t[22] = t[27] ^ x[14];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = (~t[29] & t[34]);
  assign t[28] = (~t[29] & t[35]);
  assign t[29] = t[36] ^ x[8];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[9];
  assign t[31] = t[38] ^ x[11];
  assign t[32] = t[39] ^ x[12];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[14];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[37] = (x[5]);
  assign t[38] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[4]);
  assign t[42] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[4]);
  assign t[43] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[6]);
  assign t[42] = (x[7]);
  assign t[43] = (x[4]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[40]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[42]);
  assign t[14] = ~(t[40] | t[41]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[17] : x[16];
  assign t[18] = x[2] ? x[18] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[11]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[4] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[7] | t[38];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[9];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[6]);
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = (~t[53] & t[58]);
  assign t[52] = (~t[53] & t[59]);
  assign t[53] = t[60] ^ x[8];
  assign t[54] = t[61] ^ x[9];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[61] = (x[5]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[6]);
  assign t[65] = (x[7]);
  assign t[66] = (x[4]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[38] | t[12]);
  assign t[9] = ~x[2] & t[39];
  assign y = (t[0] & ~t[15] & ~t[23] & ~t[32]) | (~t[0] & t[15] & ~t[23] & ~t[32]) | (~t[0] & ~t[15] & t[23] & ~t[32]) | (~t[0] & ~t[15] & ~t[23] & t[32]) | (t[0] & t[15] & t[23] & ~t[32]) | (t[0] & t[15] & ~t[23] & t[32]) | (t[0] & ~t[15] & t[23] & t[32]) | (~t[0] & t[15] & t[23] & t[32]);
endmodule

module R2ind76(x, y);
 input [15:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[13];
  assign t[22] = t[27] ^ x[14];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = (~t[29] & t[34]);
  assign t[28] = (~t[29] & t[35]);
  assign t[29] = t[36] ^ x[8];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[9];
  assign t[31] = t[38] ^ x[11];
  assign t[32] = t[39] ^ x[12];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[14];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[37] = (x[5]);
  assign t[38] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[4]);
  assign t[42] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[4]);
  assign t[43] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[6]);
  assign t[42] = (x[7]);
  assign t[43] = (x[4]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[40]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[42]);
  assign t[14] = ~(t[40] | t[41]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[17] : x[16];
  assign t[18] = x[2] ? x[18] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[11]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[9] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[9] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[7] | t[38];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[9];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[6]);
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = (~t[53] & t[58]);
  assign t[52] = (~t[53] & t[59]);
  assign t[53] = t[60] ^ x[8];
  assign t[54] = t[61] ^ x[9];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[61] = (x[5]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[6]);
  assign t[65] = (x[7]);
  assign t[66] = (x[4]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[38] | t[12]);
  assign t[9] = ~x[2] & t[39];
  assign y = (t[0] & ~t[15] & ~t[23] & ~t[32]) | (~t[0] & t[15] & ~t[23] & ~t[32]) | (~t[0] & ~t[15] & t[23] & ~t[32]) | (~t[0] & ~t[15] & ~t[23] & t[32]) | (t[0] & t[15] & t[23] & ~t[32]) | (t[0] & t[15] & ~t[23] & t[32]) | (t[0] & ~t[15] & t[23] & t[32]) | (~t[0] & t[15] & t[23] & t[32]);
endmodule

module R2ind81(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[8]);
  assign t[11] = ~(t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[12];
  assign t[19] = t[24] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[5];
  assign t[28] = t[35] ^ x[6];
  assign t[29] = t[36] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[12];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[14];
  assign t[33] = t[40] ^ x[15];
  assign t[34] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[4]);
  assign t[36] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[37] = (x[8]);
  assign t[38] = (x[10]);
  assign t[39] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[9]);
  assign t[4] = ~x[2] & t[12];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = t[10] | t[13];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [15:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[4]);
  assign t[37] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[38] = (x[8]);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[9]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[6]);
  assign t[42] = (x[7]);
  assign t[43] = (x[4]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [24:0] x;
 output y;

 wire [64:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[40]);
  assign t[12] = ~(t[38] | t[39]);
  assign t[13] = ~(t[14] ^ t[15]);
  assign t[14] = ~t[16];
  assign t[15] = t[4] ? x[17] : x[16];
  assign t[16] = x[2] ? x[18] : t[17];
  assign t[17] = ~(t[18] & t[19]);
  assign t[18] = ~(t[38] & t[9]);
  assign t[19] = ~(t[40] & t[20]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] & t[8]);
  assign t[21] = ~(t[22] ^ t[23]);
  assign t[22] = ~t[24];
  assign t[23] = t[4] ? x[20] : x[19];
  assign t[24] = x[2] ? x[21] : t[25];
  assign t[25] = ~(t[26] & t[27]);
  assign t[26] = ~(t[9] & t[11]);
  assign t[27] = ~(t[28] & t[37]);
  assign t[28] = ~(t[29] & t[8]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] ^ t[32]);
  assign t[31] = ~t[33];
  assign t[32] = t[4] ? x[23] : x[22];
  assign t[33] = x[2] ? x[24] : t[34];
  assign t[34] = ~(t[26] & t[35]);
  assign t[35] = t[6] | t[37];
  assign t[36] = (t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = t[46] ^ x[6];
  assign t[42] = t[47] ^ x[12];
  assign t[43] = t[48] ^ x[13];
  assign t[44] = t[49] ^ x[14];
  assign t[45] = t[50] ^ x[15];
  assign t[46] = (~t[51] & t[52]);
  assign t[47] = (~t[53] & t[54]);
  assign t[48] = (~t[53] & t[55]);
  assign t[49] = (~t[53] & t[56]);
  assign t[4] = ~x[2] & t[36];
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = t[58] ^ x[5];
  assign t[52] = t[59] ^ x[6];
  assign t[53] = t[60] ^ x[11];
  assign t[54] = t[61] ^ x[12];
  assign t[55] = t[62] ^ x[13];
  assign t[56] = t[63] ^ x[14];
  assign t[57] = t[64] ^ x[15];
  assign t[58] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[61] = (x[8]);
  assign t[62] = (x[9]);
  assign t[63] = (x[10]);
  assign t[64] = (x[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[37] | t[10]);
  assign t[8] = ~(t[38]);
  assign t[9] = ~(t[39]);
  assign y = (t[0] & ~t[13] & ~t[21] & ~t[30]) | (~t[0] & t[13] & ~t[21] & ~t[30]) | (~t[0] & ~t[13] & t[21] & ~t[30]) | (~t[0] & ~t[13] & ~t[21] & t[30]) | (t[0] & t[13] & t[21] & ~t[30]) | (t[0] & t[13] & ~t[21] & t[30]) | (t[0] & ~t[13] & t[21] & t[30]) | (~t[0] & t[13] & t[21] & t[30]);
endmodule

module R2ind86(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[8]);
  assign t[11] = ~(t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[12];
  assign t[19] = t[24] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[5];
  assign t[28] = t[35] ^ x[6];
  assign t[29] = t[36] ^ x[11];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[12];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[14];
  assign t[33] = t[40] ^ x[15];
  assign t[34] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[4]);
  assign t[36] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[37] = (x[8]);
  assign t[38] = (x[10]);
  assign t[39] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[9]);
  assign t[4] = ~x[2] & t[12];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = t[10] | t[13];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [15:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[4]);
  assign t[37] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[38] = (x[8]);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[9]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [14:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[12];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = t[22] ^ x[14];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = ~t[3];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[25] & t[27]);
  assign t[22] = (~t[25] & t[28]);
  assign t[23] = t[29] ^ x[5];
  assign t[24] = t[30] ^ x[6];
  assign t[25] = t[31] ^ x[11];
  assign t[26] = t[32] ^ x[12];
  assign t[27] = t[33] ^ x[13];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (x[4]);
  assign t[31] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[32] = (x[9]);
  assign t[33] = (x[7]);
  assign t[34] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~x[2] & t[11];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[12] & t[8]);
  assign t[7] = ~(t[13] & t[9]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[14] & t[10]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [15:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[30] & t[31]);
  assign t[25] = (~t[30] & t[32]);
  assign t[26] = (~t[30] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[4]);
  assign t[37] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[38] = (x[8]);
  assign t[39] = (x[9]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[40]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[42]);
  assign t[14] = ~(t[40] | t[41]);
  assign t[15] = ~(t[16] ^ t[17]);
  assign t[16] = ~t[18];
  assign t[17] = t[4] ? x[17] : x[16];
  assign t[18] = x[2] ? x[18] : t[19];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[40] & t[11]);
  assign t[21] = ~(t[42] & t[22]);
  assign t[22] = ~(t[41] & t[10]);
  assign t[23] = ~(t[24] ^ t[25]);
  assign t[24] = ~t[26];
  assign t[25] = t[4] ? x[20] : x[19];
  assign t[26] = x[2] ? x[21] : t[27];
  assign t[27] = ~(t[28] & t[29]);
  assign t[28] = ~(t[11] & t[13]);
  assign t[29] = ~(t[30] & t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[31] & t[10]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[33] ^ t[34]);
  assign t[33] = ~t[35];
  assign t[34] = t[4] ? x[23] : x[22];
  assign t[35] = x[2] ? x[24] : t[36];
  assign t[36] = ~(t[28] & t[37]);
  assign t[37] = t[7] | t[38];
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[9];
  assign t[44] = t[49] ^ x[12];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[14];
  assign t[47] = t[52] ^ x[15];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[6]);
  assign t[50] = (~t[53] & t[57]);
  assign t[51] = (~t[53] & t[58]);
  assign t[52] = (~t[53] & t[59]);
  assign t[53] = t[60] ^ x[8];
  assign t[54] = t[61] ^ x[9];
  assign t[55] = t[62] ^ x[11];
  assign t[56] = t[63] ^ x[12];
  assign t[57] = t[64] ^ x[13];
  assign t[58] = t[65] ^ x[14];
  assign t[59] = t[66] ^ x[15];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[61] = (x[5]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[6]);
  assign t[65] = (x[7]);
  assign t[66] = (x[4]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[38] | t[12]);
  assign t[9] = ~x[2] & t[39];
  assign y = (t[0] & ~t[15] & ~t[23] & ~t[32]) | (~t[0] & t[15] & ~t[23] & ~t[32]) | (~t[0] & ~t[15] & t[23] & ~t[32]) | (~t[0] & ~t[15] & ~t[23] & t[32]) | (t[0] & t[15] & t[23] & ~t[32]) | (t[0] & t[15] & ~t[23] & t[32]) | (t[0] & ~t[15] & t[23] & t[32]) | (~t[0] & t[15] & t[23] & t[32]);
endmodule

module R2ind91(x, y);
 input [15:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[13];
  assign t[22] = t[27] ^ x[14];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = (~t[29] & t[34]);
  assign t[28] = (~t[29] & t[35]);
  assign t[29] = t[36] ^ x[8];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[9];
  assign t[31] = t[38] ^ x[11];
  assign t[32] = t[39] ^ x[12];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[14];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[37] = (x[5]);
  assign t[38] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[10]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[4]);
  assign t[42] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[4]);
  assign t[43] = (x[6]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [14:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[10];
  assign t[19] = t[23] ^ x[13];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[14];
  assign t[21] = (~t[25] & t[26]);
  assign t[22] = (~t[25] & t[27]);
  assign t[23] = (~t[28] & t[29]);
  assign t[24] = (~t[25] & t[30]);
  assign t[25] = t[31] ^ x[8];
  assign t[26] = t[32] ^ x[9];
  assign t[27] = t[33] ^ x[10];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[36] ^ x[14];
  assign t[31] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[32] = (x[6]);
  assign t[33] = (x[4]);
  assign t[34] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[11]);
  assign t[36] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [15:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = t[29] ^ x[15];
  assign t[25] = (~t[30] & t[31]);
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[30] & t[34]);
  assign t[28] = (~t[30] & t[35]);
  assign t[29] = (~t[30] & t[36]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[8];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = (x[4] & ~x[5] & ~x[6] & ~x[7]) | (~x[4] & x[5] & ~x[6] & ~x[7]) | (~x[4] & ~x[5] & x[6] & ~x[7]) | (~x[4] & ~x[5] & ~x[6] & x[7]) | (x[4] & x[5] & x[6] & ~x[7]) | (x[4] & x[5] & ~x[6] & x[7]) | (x[4] & ~x[5] & x[6] & x[7]) | (~x[4] & x[5] & x[6] & x[7]);
  assign t[38] = (x[5]);
  assign t[39] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[10]);
  assign t[41] = (x[6]);
  assign t[42] = (x[7]);
  assign t[43] = (x[4]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [37:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[112] ^ x[18];
  assign t[101] = t[113] ^ x[19];
  assign t[102] = t[114] ^ x[20];
  assign t[103] = t[115] ^ x[21];
  assign t[104] = t[116] ^ x[22];
  assign t[105] = t[117] ^ x[23];
  assign t[106] = t[118] ^ x[24];
  assign t[107] = t[119] ^ x[25];
  assign t[108] = (x[5] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0 & ~1'b0) | (x[5] & 1'b0 & ~1'b0 & 1'b0) | (x[5] & ~1'b0 & 1'b0 & 1'b0) | (~x[5] & 1'b0 & 1'b0 & 1'b0);
  assign t[109] = (x[5]);
  assign t[10] = ~x[2] & t[69];
  assign t[110] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[111] = (x[9]);
  assign t[112] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[113] = (x[15]);
  assign t[114] = (x[10]);
  assign t[115] = (x[11]);
  assign t[116] = (x[16]);
  assign t[117] = (x[17]);
  assign t[118] = (x[8]);
  assign t[119] = (x[14]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[70] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[71] | t[21]);
  assign t[16] = ~(t[72]);
  assign t[17] = ~(t[73]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[74]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[75]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[76]);
  assign t[23] = ~(t[72] | t[73]);
  assign t[24] = ~(t[77]);
  assign t[25] = ~(t[74] | t[75]);
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~t[29];
  assign t[28] = t[10] ? x[27] : x[26];
  assign t[29] = ~(t[30] ^ t[31]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~t[32];
  assign t[31] = x[2] ? x[28] : t[33];
  assign t[32] = x[2] ? x[29] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[72] & t[17]);
  assign t[36] = ~(t[76] & t[39]);
  assign t[37] = ~(t[74] & t[20]);
  assign t[38] = ~(t[77] & t[40]);
  assign t[39] = ~(t[73] & t[16]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[75] & t[19]);
  assign t[41] = ~(t[42] ^ t[43]);
  assign t[42] = ~t[44];
  assign t[43] = t[4] ? x[31] : x[30];
  assign t[44] = ~(t[45] ^ t[46]);
  assign t[45] = ~t[47];
  assign t[46] = x[2] ? x[32] : t[48];
  assign t[47] = x[2] ? x[33] : t[49];
  assign t[48] = ~(t[50] & t[51]);
  assign t[49] = ~(t[52] & t[53]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[17] & t[22]);
  assign t[51] = ~(t[54] & t[70]);
  assign t[52] = ~(t[20] & t[24]);
  assign t[53] = ~(t[55] & t[71]);
  assign t[54] = ~(t[56] & t[16]);
  assign t[55] = ~(t[57] & t[19]);
  assign t[56] = ~(t[76] & t[73]);
  assign t[57] = ~(t[77] & t[75]);
  assign t[58] = ~(t[59] ^ t[60]);
  assign t[59] = ~t[61];
  assign t[5] = ~t[8];
  assign t[60] = t[4] ? x[35] : x[34];
  assign t[61] = ~(t[62] ^ t[63]);
  assign t[62] = ~t[64];
  assign t[63] = x[2] ? x[36] : t[65];
  assign t[64] = x[2] ? x[37] : t[66];
  assign t[65] = ~(t[50] & t[67]);
  assign t[66] = ~(t[52] & t[68]);
  assign t[67] = t[12] | t[70];
  assign t[68] = t[14] | t[71];
  assign t[69] = (t[78]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (t[79]);
  assign t[71] = (t[80]);
  assign t[72] = (t[81]);
  assign t[73] = (t[82]);
  assign t[74] = (t[83]);
  assign t[75] = (t[84]);
  assign t[76] = (t[85]);
  assign t[77] = (t[86]);
  assign t[78] = t[87] ^ x[7];
  assign t[79] = t[88] ^ x[13];
  assign t[7] = ~(t[10]);
  assign t[80] = t[89] ^ x[19];
  assign t[81] = t[90] ^ x[20];
  assign t[82] = t[91] ^ x[21];
  assign t[83] = t[92] ^ x[22];
  assign t[84] = t[93] ^ x[23];
  assign t[85] = t[94] ^ x[24];
  assign t[86] = t[95] ^ x[25];
  assign t[87] = (~t[96] & t[97]);
  assign t[88] = (~t[98] & t[99]);
  assign t[89] = (~t[100] & t[101]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[90] = (~t[98] & t[102]);
  assign t[91] = (~t[98] & t[103]);
  assign t[92] = (~t[100] & t[104]);
  assign t[93] = (~t[100] & t[105]);
  assign t[94] = (~t[98] & t[106]);
  assign t[95] = (~t[100] & t[107]);
  assign t[96] = t[108] ^ x[6];
  assign t[97] = t[109] ^ x[7];
  assign t[98] = t[110] ^ x[12];
  assign t[99] = t[111] ^ x[13];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[26] & ~t[41] & ~t[58]) | (~t[0] & t[26] & ~t[41] & ~t[58]) | (~t[0] & ~t[26] & t[41] & ~t[58]) | (~t[0] & ~t[26] & ~t[41] & t[58]) | (t[0] & t[26] & t[41] & ~t[58]) | (t[0] & t[26] & ~t[41] & t[58]) | (t[0] & ~t[26] & t[41] & t[58]) | (~t[0] & t[26] & t[41] & t[58]);
endmodule

module R2ind96(x, y);
 input [25:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[24];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = t[18] | t[25];
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = t[21] | t[26];
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[22] | t[16]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[23] | t[19]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = t[42] ^ x[7];
  assign t[34] = t[43] ^ x[13];
  assign t[35] = t[44] ^ x[19];
  assign t[36] = t[45] ^ x[20];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[22];
  assign t[39] = t[48] ^ x[23];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[24];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = (~t[51] & t[52]);
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[53] & t[57]);
  assign t[46] = (~t[53] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = (~t[55] & t[60]);
  assign t[49] = (~t[53] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[55] & t[62]);
  assign t[51] = t[63] ^ x[6];
  assign t[52] = t[64] ^ x[7];
  assign t[53] = t[65] ^ x[12];
  assign t[54] = t[66] ^ x[13];
  assign t[55] = t[67] ^ x[18];
  assign t[56] = t[68] ^ x[19];
  assign t[57] = t[69] ^ x[20];
  assign t[58] = t[70] ^ x[21];
  assign t[59] = t[71] ^ x[22];
  assign t[5] = ~t[8];
  assign t[60] = t[72] ^ x[23];
  assign t[61] = t[73] ^ x[24];
  assign t[62] = t[74] ^ x[25];
  assign t[63] = (x[5] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0 & ~1'b0) | (x[5] & 1'b0 & ~1'b0 & 1'b0) | (x[5] & ~1'b0 & 1'b0 & 1'b0) | (~x[5] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[5]);
  assign t[65] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[66] = (x[9]);
  assign t[67] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[68] = (x[15]);
  assign t[69] = (x[11]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[8]);
  assign t[71] = (x[17]);
  assign t[72] = (x[14]);
  assign t[73] = (x[10]);
  assign t[74] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [25:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[27]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[32] & t[31]);
  assign t[25] = ~(t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[20];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[23];
  assign t[42] = t[51] ^ x[24];
  assign t[43] = t[52] ^ x[25];
  assign t[44] = (~t[53] & t[54]);
  assign t[45] = (~t[55] & t[56]);
  assign t[46] = (~t[57] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = (~t[55] & t[60]);
  assign t[49] = (~t[57] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[57] & t[62]);
  assign t[51] = (~t[55] & t[63]);
  assign t[52] = (~t[57] & t[64]);
  assign t[53] = t[65] ^ x[6];
  assign t[54] = t[66] ^ x[7];
  assign t[55] = t[67] ^ x[12];
  assign t[56] = t[68] ^ x[13];
  assign t[57] = t[69] ^ x[18];
  assign t[58] = t[70] ^ x[19];
  assign t[59] = t[71] ^ x[20];
  assign t[5] = ~t[8];
  assign t[60] = t[72] ^ x[21];
  assign t[61] = t[73] ^ x[22];
  assign t[62] = t[74] ^ x[23];
  assign t[63] = t[75] ^ x[24];
  assign t[64] = t[76] ^ x[25];
  assign t[65] = (x[5] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0 & ~1'b0) | (x[5] & 1'b0 & ~1'b0 & 1'b0) | (x[5] & ~1'b0 & 1'b0 & 1'b0) | (~x[5] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[5]);
  assign t[67] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[68] = (x[9]);
  assign t[69] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[15]);
  assign t[71] = (x[11]);
  assign t[72] = (x[8]);
  assign t[73] = (x[17]);
  assign t[74] = (x[14]);
  assign t[75] = (x[10]);
  assign t[76] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [23:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[25] & t[18]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[26] & t[19]);
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[23]);
  assign t[1] = ~t[3];
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = (t[33]);
  assign t[27] = t[34] ^ x[5];
  assign t[28] = t[35] ^ x[13];
  assign t[29] = t[36] ^ x[14];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[20];
  assign t[31] = t[38] ^ x[21];
  assign t[32] = t[39] ^ x[22];
  assign t[33] = t[40] ^ x[23];
  assign t[34] = (~t[41] & t[42]);
  assign t[35] = (~t[43] & t[44]);
  assign t[36] = (~t[43] & t[45]);
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[46] & t[48]);
  assign t[39] = (~t[43] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (~t[46] & t[50]);
  assign t[41] = t[51] ^ x[4];
  assign t[42] = t[52] ^ x[5];
  assign t[43] = t[53] ^ x[12];
  assign t[44] = t[54] ^ x[13];
  assign t[45] = t[55] ^ x[14];
  assign t[46] = t[56] ^ x[19];
  assign t[47] = t[57] ^ x[20];
  assign t[48] = t[58] ^ x[21];
  assign t[49] = t[59] ^ x[22];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[60] ^ x[23];
  assign t[51] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[3]);
  assign t[53] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[54] = (x[10]);
  assign t[55] = (x[8]);
  assign t[56] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[57] = (x[17]);
  assign t[58] = (x[15]);
  assign t[59] = (x[11]);
  assign t[5] = ~t[7];
  assign t[60] = (x[18]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [25:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[27] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[28] | t[21]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[20];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[23];
  assign t[42] = t[51] ^ x[24];
  assign t[43] = t[52] ^ x[25];
  assign t[44] = (~t[53] & t[54]);
  assign t[45] = (~t[55] & t[56]);
  assign t[46] = (~t[57] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = (~t[55] & t[60]);
  assign t[49] = (~t[57] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[57] & t[62]);
  assign t[51] = (~t[55] & t[63]);
  assign t[52] = (~t[57] & t[64]);
  assign t[53] = t[65] ^ x[6];
  assign t[54] = t[66] ^ x[7];
  assign t[55] = t[67] ^ x[12];
  assign t[56] = t[68] ^ x[13];
  assign t[57] = t[69] ^ x[18];
  assign t[58] = t[70] ^ x[19];
  assign t[59] = t[71] ^ x[20];
  assign t[5] = ~t[8];
  assign t[60] = t[72] ^ x[21];
  assign t[61] = t[73] ^ x[22];
  assign t[62] = t[74] ^ x[23];
  assign t[63] = t[75] ^ x[24];
  assign t[64] = t[76] ^ x[25];
  assign t[65] = (x[5] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0 & ~1'b0) | (x[5] & 1'b0 & ~1'b0 & 1'b0) | (x[5] & ~1'b0 & 1'b0 & 1'b0) | (~x[5] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[5]);
  assign t[67] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[68] = (x[9]);
  assign t[69] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[15]);
  assign t[71] = (x[10]);
  assign t[72] = (x[11]);
  assign t[73] = (x[16]);
  assign t[74] = (x[17]);
  assign t[75] = (x[8]);
  assign t[76] = (x[14]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [37:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[112] ^ x[18];
  assign t[101] = t[113] ^ x[19];
  assign t[102] = t[114] ^ x[20];
  assign t[103] = t[115] ^ x[21];
  assign t[104] = t[116] ^ x[22];
  assign t[105] = t[117] ^ x[23];
  assign t[106] = t[118] ^ x[24];
  assign t[107] = t[119] ^ x[25];
  assign t[108] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[109] = (x[3]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[110] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[111] = (x[9]);
  assign t[112] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[113] = (x[15]);
  assign t[114] = (x[10]);
  assign t[115] = (x[11]);
  assign t[116] = (x[16]);
  assign t[117] = (x[17]);
  assign t[118] = (x[8]);
  assign t[119] = (x[14]);
  assign t[11] = ~(t[70] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[71] | t[19]);
  assign t[14] = ~(t[72]);
  assign t[15] = ~(t[73]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[74]);
  assign t[18] = ~(t[75]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[76]);
  assign t[21] = ~(t[72] | t[73]);
  assign t[22] = ~(t[77]);
  assign t[23] = ~(t[74] | t[75]);
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~t[27];
  assign t[26] = t[28] ? x[27] : x[26];
  assign t[27] = ~(t[29] ^ t[30]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~t[32];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = x[2] ? x[28] : t[33];
  assign t[31] = ~(t[4]);
  assign t[32] = x[2] ? x[29] : t[34];
  assign t[33] = ~(t[35] & t[36]);
  assign t[34] = ~(t[37] & t[38]);
  assign t[35] = ~(t[72] & t[15]);
  assign t[36] = ~(t[76] & t[39]);
  assign t[37] = ~(t[74] & t[18]);
  assign t[38] = ~(t[77] & t[40]);
  assign t[39] = ~(t[73] & t[14]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[75] & t[17]);
  assign t[41] = ~(t[42] ^ t[43]);
  assign t[42] = ~t[44];
  assign t[43] = t[28] ? x[31] : x[30];
  assign t[44] = ~(t[45] ^ t[46]);
  assign t[45] = ~t[47];
  assign t[46] = x[2] ? x[32] : t[48];
  assign t[47] = x[2] ? x[33] : t[49];
  assign t[48] = ~(t[50] & t[51]);
  assign t[49] = ~(t[52] & t[53]);
  assign t[4] = ~x[2] & t[69];
  assign t[50] = ~(t[15] & t[20]);
  assign t[51] = ~(t[54] & t[70]);
  assign t[52] = ~(t[18] & t[22]);
  assign t[53] = ~(t[55] & t[71]);
  assign t[54] = ~(t[56] & t[14]);
  assign t[55] = ~(t[57] & t[17]);
  assign t[56] = ~(t[76] & t[73]);
  assign t[57] = ~(t[77] & t[75]);
  assign t[58] = ~(t[59] ^ t[60]);
  assign t[59] = ~t[61];
  assign t[5] = ~t[7];
  assign t[60] = t[4] ? x[35] : x[34];
  assign t[61] = ~(t[62] ^ t[63]);
  assign t[62] = ~t[64];
  assign t[63] = x[2] ? x[36] : t[65];
  assign t[64] = x[2] ? x[37] : t[66];
  assign t[65] = ~(t[50] & t[67]);
  assign t[66] = ~(t[52] & t[68]);
  assign t[67] = t[10] | t[70];
  assign t[68] = t[12] | t[71];
  assign t[69] = (t[78]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (t[79]);
  assign t[71] = (t[80]);
  assign t[72] = (t[81]);
  assign t[73] = (t[82]);
  assign t[74] = (t[83]);
  assign t[75] = (t[84]);
  assign t[76] = (t[85]);
  assign t[77] = (t[86]);
  assign t[78] = t[87] ^ x[5];
  assign t[79] = t[88] ^ x[13];
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[80] = t[89] ^ x[19];
  assign t[81] = t[90] ^ x[20];
  assign t[82] = t[91] ^ x[21];
  assign t[83] = t[92] ^ x[22];
  assign t[84] = t[93] ^ x[23];
  assign t[85] = t[94] ^ x[24];
  assign t[86] = t[95] ^ x[25];
  assign t[87] = (~t[96] & t[97]);
  assign t[88] = (~t[98] & t[99]);
  assign t[89] = (~t[100] & t[101]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[90] = (~t[98] & t[102]);
  assign t[91] = (~t[98] & t[103]);
  assign t[92] = (~t[100] & t[104]);
  assign t[93] = (~t[100] & t[105]);
  assign t[94] = (~t[98] & t[106]);
  assign t[95] = (~t[100] & t[107]);
  assign t[96] = t[108] ^ x[4];
  assign t[97] = t[109] ^ x[5];
  assign t[98] = t[110] ^ x[12];
  assign t[99] = t[111] ^ x[13];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0] & ~t[24] & ~t[41] & ~t[58]) | (~t[0] & t[24] & ~t[41] & ~t[58]) | (~t[0] & ~t[24] & t[41] & ~t[58]) | (~t[0] & ~t[24] & ~t[41] & t[58]) | (t[0] & t[24] & t[41] & ~t[58]) | (t[0] & t[24] & ~t[41] & t[58]) | (t[0] & ~t[24] & t[41] & t[58]) | (~t[0] & t[24] & t[41] & t[58]);
endmodule

module R2ind101(x, y);
 input [25:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = t[16] | t[23];
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[24];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[20] | t[14]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[21] | t[17]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29]);
  assign t[21] = ~(t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = t[40] ^ x[5];
  assign t[32] = t[41] ^ x[13];
  assign t[33] = t[42] ^ x[19];
  assign t[34] = t[43] ^ x[20];
  assign t[35] = t[44] ^ x[21];
  assign t[36] = t[45] ^ x[22];
  assign t[37] = t[46] ^ x[23];
  assign t[38] = t[47] ^ x[24];
  assign t[39] = t[48] ^ x[25];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (~t[49] & t[50]);
  assign t[41] = (~t[51] & t[52]);
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[51] & t[55]);
  assign t[44] = (~t[51] & t[56]);
  assign t[45] = (~t[53] & t[57]);
  assign t[46] = (~t[53] & t[58]);
  assign t[47] = (~t[51] & t[59]);
  assign t[48] = (~t[53] & t[60]);
  assign t[49] = t[61] ^ x[4];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[62] ^ x[5];
  assign t[51] = t[63] ^ x[12];
  assign t[52] = t[64] ^ x[13];
  assign t[53] = t[65] ^ x[18];
  assign t[54] = t[66] ^ x[19];
  assign t[55] = t[67] ^ x[20];
  assign t[56] = t[68] ^ x[21];
  assign t[57] = t[69] ^ x[22];
  assign t[58] = t[70] ^ x[23];
  assign t[59] = t[71] ^ x[24];
  assign t[5] = ~t[7];
  assign t[60] = t[72] ^ x[25];
  assign t[61] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[3]);
  assign t[63] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[64] = (x[9]);
  assign t[65] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[66] = (x[15]);
  assign t[67] = (x[11]);
  assign t[68] = (x[8]);
  assign t[69] = (x[17]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (x[14]);
  assign t[71] = (x[10]);
  assign t[72] = (x[16]);
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [25:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[27]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[32] & t[31]);
  assign t[25] = ~(t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[20];
  assign t[39] = t[48] ^ x[21];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[23];
  assign t[42] = t[51] ^ x[24];
  assign t[43] = t[52] ^ x[25];
  assign t[44] = (~t[53] & t[54]);
  assign t[45] = (~t[55] & t[56]);
  assign t[46] = (~t[57] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = (~t[55] & t[60]);
  assign t[49] = (~t[57] & t[61]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[57] & t[62]);
  assign t[51] = (~t[55] & t[63]);
  assign t[52] = (~t[57] & t[64]);
  assign t[53] = t[65] ^ x[6];
  assign t[54] = t[66] ^ x[7];
  assign t[55] = t[67] ^ x[12];
  assign t[56] = t[68] ^ x[13];
  assign t[57] = t[69] ^ x[18];
  assign t[58] = t[70] ^ x[19];
  assign t[59] = t[71] ^ x[20];
  assign t[5] = ~t[8];
  assign t[60] = t[72] ^ x[21];
  assign t[61] = t[73] ^ x[22];
  assign t[62] = t[74] ^ x[23];
  assign t[63] = t[75] ^ x[24];
  assign t[64] = t[76] ^ x[25];
  assign t[65] = (x[5] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0 & ~1'b0) | (x[5] & 1'b0 & ~1'b0 & 1'b0) | (x[5] & ~1'b0 & 1'b0 & 1'b0) | (~x[5] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[5]);
  assign t[67] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[68] = (x[9]);
  assign t[69] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[15]);
  assign t[71] = (x[11]);
  assign t[72] = (x[8]);
  assign t[73] = (x[17]);
  assign t[74] = (x[14]);
  assign t[75] = (x[10]);
  assign t[76] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [23:0] x;
 output y;

 wire [62:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[22];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25] & t[18]);
  assign t[15] = ~(t[26] & t[19]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[27] & t[20]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[28] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[25]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = (t[33]);
  assign t[27] = (t[34]);
  assign t[28] = (t[35]);
  assign t[29] = t[36] ^ x[7];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[13];
  assign t[31] = t[38] ^ x[14];
  assign t[32] = t[39] ^ x[20];
  assign t[33] = t[40] ^ x[21];
  assign t[34] = t[41] ^ x[22];
  assign t[35] = t[42] ^ x[23];
  assign t[36] = (~t[43] & t[44]);
  assign t[37] = (~t[45] & t[46]);
  assign t[38] = (~t[45] & t[47]);
  assign t[39] = (~t[48] & t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (~t[48] & t[50]);
  assign t[41] = (~t[45] & t[51]);
  assign t[42] = (~t[48] & t[52]);
  assign t[43] = t[53] ^ x[6];
  assign t[44] = t[54] ^ x[7];
  assign t[45] = t[55] ^ x[12];
  assign t[46] = t[56] ^ x[13];
  assign t[47] = t[57] ^ x[14];
  assign t[48] = t[58] ^ x[19];
  assign t[49] = t[59] ^ x[20];
  assign t[4] = ~(t[7]);
  assign t[50] = t[60] ^ x[21];
  assign t[51] = t[61] ^ x[22];
  assign t[52] = t[62] ^ x[23];
  assign t[53] = (x[5] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[5] & 1'b0 & ~1'b0 & ~1'b0) | (~x[5] & ~1'b0 & 1'b0 & ~1'b0) | (~x[5] & ~1'b0 & ~1'b0 & 1'b0) | (x[5] & 1'b0 & 1'b0 & ~1'b0) | (x[5] & 1'b0 & ~1'b0 & 1'b0) | (x[5] & ~1'b0 & 1'b0 & 1'b0) | (~x[5] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[5]);
  assign t[55] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[56] = (x[10]);
  assign t[57] = (x[8]);
  assign t[58] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[59] = (x[17]);
  assign t[5] = ~t[8];
  assign t[60] = (x[15]);
  assign t[61] = (x[11]);
  assign t[62] = (x[18]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [25:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[25] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[26] | t[19]);
  assign t[14] = ~(t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[27] | t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = t[42] ^ x[5];
  assign t[34] = t[43] ^ x[13];
  assign t[35] = t[44] ^ x[19];
  assign t[36] = t[45] ^ x[20];
  assign t[37] = t[46] ^ x[21];
  assign t[38] = t[47] ^ x[22];
  assign t[39] = t[48] ^ x[23];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[24];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = (~t[51] & t[52]);
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[53] & t[57]);
  assign t[46] = (~t[53] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = (~t[55] & t[60]);
  assign t[49] = (~t[53] & t[61]);
  assign t[4] = ~x[2] & t[24];
  assign t[50] = (~t[55] & t[62]);
  assign t[51] = t[63] ^ x[4];
  assign t[52] = t[64] ^ x[5];
  assign t[53] = t[65] ^ x[12];
  assign t[54] = t[66] ^ x[13];
  assign t[55] = t[67] ^ x[18];
  assign t[56] = t[68] ^ x[19];
  assign t[57] = t[69] ^ x[20];
  assign t[58] = t[70] ^ x[21];
  assign t[59] = t[71] ^ x[22];
  assign t[5] = ~t[7];
  assign t[60] = t[72] ^ x[23];
  assign t[61] = t[73] ^ x[24];
  assign t[62] = t[74] ^ x[25];
  assign t[63] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[3]);
  assign t[65] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[66] = (x[9]);
  assign t[67] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[68] = (x[15]);
  assign t[69] = (x[10]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (x[11]);
  assign t[71] = (x[16]);
  assign t[72] = (x[17]);
  assign t[73] = (x[8]);
  assign t[74] = (x[14]);
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [46:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (~t[112] & t[113]);
  assign t[101] = (~t[114] & t[115]);
  assign t[102] = (~t[116] & t[117]);
  assign t[103] = (~t[118] & t[119]);
  assign t[104] = (~t[114] & t[120]);
  assign t[105] = (~t[114] & t[121]);
  assign t[106] = (~t[118] & t[122]);
  assign t[107] = (~t[118] & t[123]);
  assign t[108] = (~t[114] & t[124]);
  assign t[109] = (~t[118] & t[125]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (~t[126] & t[127]);
  assign t[111] = (~t[128] & t[129]);
  assign t[112] = t[130] ^ x[4];
  assign t[113] = t[131] ^ x[5];
  assign t[114] = t[132] ^ x[12];
  assign t[115] = t[133] ^ x[13];
  assign t[116] = t[134] ^ x[15];
  assign t[117] = t[135] ^ x[16];
  assign t[118] = t[136] ^ x[21];
  assign t[119] = t[137] ^ x[22];
  assign t[11] = ~(t[15]);
  assign t[120] = t[138] ^ x[23];
  assign t[121] = t[139] ^ x[24];
  assign t[122] = t[140] ^ x[25];
  assign t[123] = t[141] ^ x[26];
  assign t[124] = t[142] ^ x[27];
  assign t[125] = t[143] ^ x[28];
  assign t[126] = t[144] ^ x[32];
  assign t[127] = t[145] ^ x[33];
  assign t[128] = t[146] ^ x[39];
  assign t[129] = t[147] ^ x[40];
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[3]);
  assign t[132] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[133] = (x[9]);
  assign t[134] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[135] = (x[14]);
  assign t[136] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[137] = (x[18]);
  assign t[138] = (x[10]);
  assign t[139] = (x[11]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = (x[19]);
  assign t[141] = (x[20]);
  assign t[142] = (x[8]);
  assign t[143] = (x[17]);
  assign t[144] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[145] = (x[31]);
  assign t[146] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[147] = (x[38]);
  assign t[14] = ~(t[77] | t[20]);
  assign t[15] = ~x[2] & t[78];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[79] | t[23]);
  assign t[18] = ~(t[80]);
  assign t[19] = ~(t[81]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[82]);
  assign t[22] = ~(t[83]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[84]);
  assign t[25] = ~(t[80] | t[81]);
  assign t[26] = ~(t[85]);
  assign t[27] = ~(t[82] | t[83]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[30] : x[29];
  assign t[33] = ~x[2] & t[86];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[34] : t[37];
  assign t[36] = x[2] ? x[35] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[80] & t[19]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[84] & t[43]);
  assign t[41] = ~(t[82] & t[22]);
  assign t[42] = ~(t[85] & t[44]);
  assign t[43] = ~(t[81] & t[18]);
  assign t[44] = ~(t[83] & t[21]);
  assign t[45] = ~(t[46] ^ t[47]);
  assign t[46] = t[48];
  assign t[47] = ~(t[49] ^ t[50]);
  assign t[48] = ~(t[51] ^ t[52]);
  assign t[49] = t[8] ? x[37] : x[36];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = ~x[2] & t[87];
  assign t[51] = ~t[53];
  assign t[52] = x[2] ? x[41] : t[54];
  assign t[53] = x[2] ? x[42] : t[55];
  assign t[54] = ~(t[56] & t[57]);
  assign t[55] = ~(t[58] & t[59]);
  assign t[56] = ~(t[19] & t[24]);
  assign t[57] = ~(t[60] & t[77]);
  assign t[58] = ~(t[22] & t[26]);
  assign t[59] = ~(t[61] & t[79]);
  assign t[5] = ~(~x[2] & ~t[76]);
  assign t[60] = ~(t[62] & t[18]);
  assign t[61] = ~(t[63] & t[21]);
  assign t[62] = ~(t[84] & t[81]);
  assign t[63] = ~(t[85] & t[83]);
  assign t[64] = ~(t[65] ^ t[66]);
  assign t[65] = t[67];
  assign t[66] = ~t[68];
  assign t[67] = ~(t[69] ^ t[70]);
  assign t[68] = t[8] ? x[44] : x[43];
  assign t[69] = ~t[71];
  assign t[6] = ~t[9];
  assign t[70] = x[2] ? x[45] : t[72];
  assign t[71] = x[2] ? x[46] : t[73];
  assign t[72] = ~(t[56] & t[74]);
  assign t[73] = ~(t[58] & t[75]);
  assign t[74] = t[13] | t[77];
  assign t[75] = t[16] | t[79];
  assign t[76] = (t[88]);
  assign t[77] = (t[89]);
  assign t[78] = (t[90]);
  assign t[79] = (t[91]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (t[92]);
  assign t[81] = (t[93]);
  assign t[82] = (t[94]);
  assign t[83] = (t[95]);
  assign t[84] = (t[96]);
  assign t[85] = (t[97]);
  assign t[86] = (t[98]);
  assign t[87] = (t[99]);
  assign t[88] = t[100] ^ x[5];
  assign t[89] = t[101] ^ x[13];
  assign t[8] = ~(t[11]);
  assign t[90] = t[102] ^ x[16];
  assign t[91] = t[103] ^ x[22];
  assign t[92] = t[104] ^ x[23];
  assign t[93] = t[105] ^ x[24];
  assign t[94] = t[106] ^ x[25];
  assign t[95] = t[107] ^ x[26];
  assign t[96] = t[108] ^ x[27];
  assign t[97] = t[109] ^ x[28];
  assign t[98] = t[110] ^ x[33];
  assign t[99] = t[111] ^ x[40];
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0] & ~t[28] & ~t[45] & ~t[64]) | (~t[0] & t[28] & ~t[45] & ~t[64]) | (~t[0] & ~t[28] & t[45] & ~t[64]) | (~t[0] & ~t[28] & ~t[45] & t[64]) | (t[0] & t[28] & t[45] & ~t[64]) | (t[0] & t[28] & ~t[45] & t[64]) | (t[0] & ~t[28] & t[45] & t[64]) | (~t[0] & t[28] & t[45] & t[64]);
endmodule

module R2ind106(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[25];
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = t[22] | t[27];
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[23] | t[17]);
  assign t[1] = t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[24] | t[20]);
  assign t[23] = ~(t[32]);
  assign t[24] = ~(t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[10];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[19];
  assign t[37] = t[46] ^ x[20];
  assign t[38] = t[47] ^ x[21];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[23];
  assign t[41] = t[50] ^ x[24];
  assign t[42] = t[51] ^ x[25];
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[56] & t[57]);
  assign t[46] = (~t[52] & t[58]);
  assign t[47] = (~t[52] & t[59]);
  assign t[48] = (~t[56] & t[60]);
  assign t[49] = (~t[56] & t[61]);
  assign t[4] = t[7] ? x[1] : x[0];
  assign t[50] = (~t[52] & t[62]);
  assign t[51] = (~t[56] & t[63]);
  assign t[52] = t[64] ^ x[9];
  assign t[53] = t[65] ^ x[10];
  assign t[54] = t[66] ^ x[12];
  assign t[55] = t[67] ^ x[13];
  assign t[56] = t[68] ^ x[18];
  assign t[57] = t[69] ^ x[19];
  assign t[58] = t[70] ^ x[20];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = ~t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[23];
  assign t[62] = t[74] ^ x[24];
  assign t[63] = t[75] ^ x[25];
  assign t[64] = (x[5] & ~x[6] & ~x[7] & ~x[8]) | (~x[5] & x[6] & ~x[7] & ~x[8]) | (~x[5] & ~x[6] & x[7] & ~x[8]) | (~x[5] & ~x[6] & ~x[7] & x[8]) | (x[5] & x[6] & x[7] & ~x[8]) | (x[5] & x[6] & ~x[7] & x[8]) | (x[5] & ~x[6] & x[7] & x[8]) | (~x[5] & x[6] & x[7] & x[8]);
  assign t[65] = (x[6]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[11]);
  assign t[68] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[69] = (x[15]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[8]);
  assign t[71] = (x[5]);
  assign t[72] = (x[17]);
  assign t[73] = (x[14]);
  assign t[74] = (x[7]);
  assign t[75] = (x[16]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [28:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[29]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[33] & t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] & t[34]);
  assign t[27] = ~(t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[13];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[22];
  assign t[42] = t[52] ^ x[23];
  assign t[43] = t[53] ^ x[24];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[26];
  assign t[46] = t[56] ^ x[27];
  assign t[47] = t[57] ^ x[28];
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = (~t[60] & t[66]);
  assign t[53] = (~t[60] & t[67]);
  assign t[54] = (~t[64] & t[68]);
  assign t[55] = (~t[64] & t[69]);
  assign t[56] = (~t[60] & t[70]);
  assign t[57] = (~t[64] & t[71]);
  assign t[58] = t[72] ^ x[4];
  assign t[59] = t[73] ^ x[5];
  assign t[5] = ~x[2] & t[28];
  assign t[60] = t[74] ^ x[12];
  assign t[61] = t[75] ^ x[13];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[16];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[22];
  assign t[66] = t[80] ^ x[23];
  assign t[67] = t[81] ^ x[24];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[26];
  assign t[6] = ~t[9];
  assign t[70] = t[84] ^ x[27];
  assign t[71] = t[85] ^ x[28];
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[75] = (x[9]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[18]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[11]);
  assign t[81] = (x[8]);
  assign t[82] = (x[20]);
  assign t[83] = (x[17]);
  assign t[84] = (x[10]);
  assign t[85] = (x[19]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [26:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~(t[26] & t[19]);
  assign t[15] = ~x[2] & t[27];
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29] & t[21]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[31] & t[23]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[28]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[13];
  assign t[34] = t[42] ^ x[14];
  assign t[35] = t[43] ^ x[17];
  assign t[36] = t[44] ^ x[23];
  assign t[37] = t[45] ^ x[24];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = t[47] ^ x[26];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = (~t[48] & t[49]);
  assign t[41] = (~t[50] & t[51]);
  assign t[42] = (~t[50] & t[52]);
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[55] & t[57]);
  assign t[46] = (~t[50] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = t[60] ^ x[4];
  assign t[49] = t[61] ^ x[5];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = t[62] ^ x[12];
  assign t[51] = t[63] ^ x[13];
  assign t[52] = t[64] ^ x[14];
  assign t[53] = t[65] ^ x[16];
  assign t[54] = t[66] ^ x[17];
  assign t[55] = t[67] ^ x[22];
  assign t[56] = t[68] ^ x[23];
  assign t[57] = t[69] ^ x[24];
  assign t[58] = t[70] ^ x[25];
  assign t[59] = t[71] ^ x[26];
  assign t[5] = ~x[2] & t[24];
  assign t[60] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[3]);
  assign t[62] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[63] = (x[10]);
  assign t[64] = (x[8]);
  assign t[65] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[15]);
  assign t[67] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[68] = (x[20]);
  assign t[69] = (x[18]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[21]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [28:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[29] | t[20]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[31] | t[23]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[13];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[22];
  assign t[42] = t[52] ^ x[23];
  assign t[43] = t[53] ^ x[24];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[26];
  assign t[46] = t[56] ^ x[27];
  assign t[47] = t[57] ^ x[28];
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = (~t[60] & t[66]);
  assign t[53] = (~t[60] & t[67]);
  assign t[54] = (~t[64] & t[68]);
  assign t[55] = (~t[64] & t[69]);
  assign t[56] = (~t[60] & t[70]);
  assign t[57] = (~t[64] & t[71]);
  assign t[58] = t[72] ^ x[4];
  assign t[59] = t[73] ^ x[5];
  assign t[5] = ~(~x[2] & ~t[28]);
  assign t[60] = t[74] ^ x[12];
  assign t[61] = t[75] ^ x[13];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[16];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[22];
  assign t[66] = t[80] ^ x[23];
  assign t[67] = t[81] ^ x[24];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[26];
  assign t[6] = ~t[9];
  assign t[70] = t[84] ^ x[27];
  assign t[71] = t[85] ^ x[28];
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[75] = (x[9]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[18]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[10]);
  assign t[81] = (x[11]);
  assign t[82] = (x[19]);
  assign t[83] = (x[20]);
  assign t[84] = (x[8]);
  assign t[85] = (x[17]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [49:0] x;
 output y;

 wire [155:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[113] ^ x[33];
  assign t[101] = t[114] ^ x[40];
  assign t[102] = t[115] ^ x[47];
  assign t[103] = (~t[116] & t[117]);
  assign t[104] = (~t[118] & t[119]);
  assign t[105] = (~t[120] & t[121]);
  assign t[106] = (~t[122] & t[123]);
  assign t[107] = (~t[118] & t[124]);
  assign t[108] = (~t[118] & t[125]);
  assign t[109] = (~t[122] & t[126]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (~t[122] & t[127]);
  assign t[111] = (~t[118] & t[128]);
  assign t[112] = (~t[122] & t[129]);
  assign t[113] = (~t[130] & t[131]);
  assign t[114] = (~t[132] & t[133]);
  assign t[115] = (~t[134] & t[135]);
  assign t[116] = t[136] ^ x[4];
  assign t[117] = t[137] ^ x[5];
  assign t[118] = t[138] ^ x[12];
  assign t[119] = t[139] ^ x[13];
  assign t[11] = ~(t[15]);
  assign t[120] = t[140] ^ x[15];
  assign t[121] = t[141] ^ x[16];
  assign t[122] = t[142] ^ x[21];
  assign t[123] = t[143] ^ x[22];
  assign t[124] = t[144] ^ x[23];
  assign t[125] = t[145] ^ x[24];
  assign t[126] = t[146] ^ x[25];
  assign t[127] = t[147] ^ x[26];
  assign t[128] = t[148] ^ x[27];
  assign t[129] = t[149] ^ x[28];
  assign t[12] = ~(t[16] | t[17]);
  assign t[130] = t[150] ^ x[32];
  assign t[131] = t[151] ^ x[33];
  assign t[132] = t[152] ^ x[39];
  assign t[133] = t[153] ^ x[40];
  assign t[134] = t[154] ^ x[46];
  assign t[135] = t[155] ^ x[47];
  assign t[136] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[137] = (x[3]);
  assign t[138] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[140] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[141] = (x[14]);
  assign t[142] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[143] = (x[18]);
  assign t[144] = (x[10]);
  assign t[145] = (x[11]);
  assign t[146] = (x[19]);
  assign t[147] = (x[20]);
  assign t[148] = (x[8]);
  assign t[149] = (x[17]);
  assign t[14] = ~(t[78] | t[20]);
  assign t[150] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[151] = (x[31]);
  assign t[152] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[38]);
  assign t[154] = (x[45] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0 & ~1'b0) | (x[45] & 1'b0 & ~1'b0 & 1'b0) | (x[45] & ~1'b0 & 1'b0 & 1'b0) | (~x[45] & 1'b0 & 1'b0 & 1'b0);
  assign t[155] = (x[45]);
  assign t[15] = ~x[2] & t[79];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[80] | t[23]);
  assign t[18] = ~(t[81]);
  assign t[19] = ~(t[82]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[83]);
  assign t[22] = ~(t[84]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[85]);
  assign t[25] = ~(t[81] | t[82]);
  assign t[26] = ~(t[86]);
  assign t[27] = ~(t[83] | t[84]);
  assign t[28] = ~(t[29] ^ t[30]);
  assign t[29] = t[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[32] ^ t[33]);
  assign t[31] = ~(t[34] ^ t[35]);
  assign t[32] = t[8] ? x[30] : x[29];
  assign t[33] = ~x[2] & t[87];
  assign t[34] = ~t[36];
  assign t[35] = x[2] ? x[34] : t[37];
  assign t[36] = x[2] ? x[35] : t[38];
  assign t[37] = ~(t[39] & t[40]);
  assign t[38] = ~(t[41] & t[42]);
  assign t[39] = ~(t[81] & t[19]);
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = ~(t[85] & t[43]);
  assign t[41] = ~(t[83] & t[22]);
  assign t[42] = ~(t[86] & t[44]);
  assign t[43] = ~(t[82] & t[18]);
  assign t[44] = ~(t[84] & t[21]);
  assign t[45] = ~(t[46] ^ t[47]);
  assign t[46] = t[48];
  assign t[47] = ~(t[49] ^ t[50]);
  assign t[48] = ~(t[51] ^ t[52]);
  assign t[49] = t[8] ? x[37] : x[36];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = ~x[2] & t[88];
  assign t[51] = ~t[53];
  assign t[52] = x[2] ? x[41] : t[54];
  assign t[53] = x[2] ? x[42] : t[55];
  assign t[54] = ~(t[56] & t[57]);
  assign t[55] = ~(t[58] & t[59]);
  assign t[56] = ~(t[19] & t[24]);
  assign t[57] = ~(t[60] & t[78]);
  assign t[58] = ~(t[22] & t[26]);
  assign t[59] = ~(t[61] & t[80]);
  assign t[5] = ~(~x[2] & ~t[77]);
  assign t[60] = ~(t[62] & t[18]);
  assign t[61] = ~(t[63] & t[21]);
  assign t[62] = ~(t[85] & t[82]);
  assign t[63] = ~(t[86] & t[84]);
  assign t[64] = ~(t[65] ^ t[66]);
  assign t[65] = t[67];
  assign t[66] = ~(t[68] ^ t[69]);
  assign t[67] = ~(t[70] ^ t[71]);
  assign t[68] = t[8] ? x[44] : x[43];
  assign t[69] = ~x[2] & t[89];
  assign t[6] = ~t[9];
  assign t[70] = ~t[72];
  assign t[71] = x[2] ? x[48] : t[73];
  assign t[72] = x[2] ? x[49] : t[74];
  assign t[73] = ~(t[56] & t[75]);
  assign t[74] = ~(t[58] & t[76]);
  assign t[75] = t[13] | t[78];
  assign t[76] = t[16] | t[80];
  assign t[77] = (t[90]);
  assign t[78] = (t[91]);
  assign t[79] = (t[92]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (t[93]);
  assign t[81] = (t[94]);
  assign t[82] = (t[95]);
  assign t[83] = (t[96]);
  assign t[84] = (t[97]);
  assign t[85] = (t[98]);
  assign t[86] = (t[99]);
  assign t[87] = (t[100]);
  assign t[88] = (t[101]);
  assign t[89] = (t[102]);
  assign t[8] = ~(t[11]);
  assign t[90] = t[103] ^ x[5];
  assign t[91] = t[104] ^ x[13];
  assign t[92] = t[105] ^ x[16];
  assign t[93] = t[106] ^ x[22];
  assign t[94] = t[107] ^ x[23];
  assign t[95] = t[108] ^ x[24];
  assign t[96] = t[109] ^ x[25];
  assign t[97] = t[110] ^ x[26];
  assign t[98] = t[111] ^ x[27];
  assign t[99] = t[112] ^ x[28];
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0] & ~t[28] & ~t[45] & ~t[64]) | (~t[0] & t[28] & ~t[45] & ~t[64]) | (~t[0] & ~t[28] & t[45] & ~t[64]) | (~t[0] & ~t[28] & ~t[45] & t[64]) | (t[0] & t[28] & t[45] & ~t[64]) | (t[0] & t[28] & ~t[45] & t[64]) | (t[0] & ~t[28] & t[45] & t[64]) | (~t[0] & t[28] & t[45] & t[64]);
endmodule

module R2ind111(x, y);
 input [28:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = t[20] | t[27];
  assign t[15] = ~x[2] & t[28];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = t[23] | t[29];
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[18]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[25] | t[21]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = t[46] ^ x[5];
  assign t[37] = t[47] ^ x[13];
  assign t[38] = t[48] ^ x[16];
  assign t[39] = t[49] ^ x[22];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[23];
  assign t[41] = t[51] ^ x[24];
  assign t[42] = t[52] ^ x[25];
  assign t[43] = t[53] ^ x[26];
  assign t[44] = t[54] ^ x[27];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = (~t[56] & t[57]);
  assign t[47] = (~t[58] & t[59]);
  assign t[48] = (~t[60] & t[61]);
  assign t[49] = (~t[62] & t[63]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (~t[58] & t[64]);
  assign t[51] = (~t[58] & t[65]);
  assign t[52] = (~t[62] & t[66]);
  assign t[53] = (~t[62] & t[67]);
  assign t[54] = (~t[58] & t[68]);
  assign t[55] = (~t[62] & t[69]);
  assign t[56] = t[70] ^ x[4];
  assign t[57] = t[71] ^ x[5];
  assign t[58] = t[72] ^ x[12];
  assign t[59] = t[73] ^ x[13];
  assign t[5] = ~x[2] & t[26];
  assign t[60] = t[74] ^ x[15];
  assign t[61] = t[75] ^ x[16];
  assign t[62] = t[76] ^ x[21];
  assign t[63] = t[77] ^ x[22];
  assign t[64] = t[78] ^ x[23];
  assign t[65] = t[79] ^ x[24];
  assign t[66] = t[80] ^ x[25];
  assign t[67] = t[81] ^ x[26];
  assign t[68] = t[82] ^ x[27];
  assign t[69] = t[83] ^ x[28];
  assign t[6] = ~t[9];
  assign t[70] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[3]);
  assign t[72] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[73] = (x[9]);
  assign t[74] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[14]);
  assign t[76] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[77] = (x[18]);
  assign t[78] = (x[11]);
  assign t[79] = (x[8]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[20]);
  assign t[81] = (x[17]);
  assign t[82] = (x[10]);
  assign t[83] = (x[19]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [28:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[29]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[33] & t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] & t[34]);
  assign t[27] = ~(t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[13];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[22];
  assign t[42] = t[52] ^ x[23];
  assign t[43] = t[53] ^ x[24];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[26];
  assign t[46] = t[56] ^ x[27];
  assign t[47] = t[57] ^ x[28];
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = (~t[60] & t[66]);
  assign t[53] = (~t[60] & t[67]);
  assign t[54] = (~t[64] & t[68]);
  assign t[55] = (~t[64] & t[69]);
  assign t[56] = (~t[60] & t[70]);
  assign t[57] = (~t[64] & t[71]);
  assign t[58] = t[72] ^ x[4];
  assign t[59] = t[73] ^ x[5];
  assign t[5] = ~x[2] & t[28];
  assign t[60] = t[74] ^ x[12];
  assign t[61] = t[75] ^ x[13];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[16];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[22];
  assign t[66] = t[80] ^ x[23];
  assign t[67] = t[81] ^ x[24];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[26];
  assign t[6] = ~t[9];
  assign t[70] = t[84] ^ x[27];
  assign t[71] = t[85] ^ x[28];
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[75] = (x[9]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[18]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[11]);
  assign t[81] = (x[8]);
  assign t[82] = (x[20]);
  assign t[83] = (x[17]);
  assign t[84] = (x[10]);
  assign t[85] = (x[19]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [26:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~(t[26] & t[19]);
  assign t[15] = ~x[2] & t[27];
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29] & t[21]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[31] & t[23]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[28]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[13];
  assign t[34] = t[42] ^ x[14];
  assign t[35] = t[43] ^ x[17];
  assign t[36] = t[44] ^ x[23];
  assign t[37] = t[45] ^ x[24];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = t[47] ^ x[26];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = (~t[48] & t[49]);
  assign t[41] = (~t[50] & t[51]);
  assign t[42] = (~t[50] & t[52]);
  assign t[43] = (~t[53] & t[54]);
  assign t[44] = (~t[55] & t[56]);
  assign t[45] = (~t[55] & t[57]);
  assign t[46] = (~t[50] & t[58]);
  assign t[47] = (~t[55] & t[59]);
  assign t[48] = t[60] ^ x[4];
  assign t[49] = t[61] ^ x[5];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = t[62] ^ x[12];
  assign t[51] = t[63] ^ x[13];
  assign t[52] = t[64] ^ x[14];
  assign t[53] = t[65] ^ x[16];
  assign t[54] = t[66] ^ x[17];
  assign t[55] = t[67] ^ x[22];
  assign t[56] = t[68] ^ x[23];
  assign t[57] = t[69] ^ x[24];
  assign t[58] = t[70] ^ x[25];
  assign t[59] = t[71] ^ x[26];
  assign t[5] = ~x[2] & t[24];
  assign t[60] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[3]);
  assign t[62] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[63] = (x[10]);
  assign t[64] = (x[8]);
  assign t[65] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[15]);
  assign t[67] = (x[18] & ~x[19] & ~x[20] & ~x[21]) | (~x[18] & x[19] & ~x[20] & ~x[21]) | (~x[18] & ~x[19] & x[20] & ~x[21]) | (~x[18] & ~x[19] & ~x[20] & x[21]) | (x[18] & x[19] & x[20] & ~x[21]) | (x[18] & x[19] & ~x[20] & x[21]) | (x[18] & ~x[19] & x[20] & x[21]) | (~x[18] & x[19] & x[20] & x[21]);
  assign t[68] = (x[20]);
  assign t[69] = (x[18]);
  assign t[6] = ~t[9];
  assign t[70] = (x[11]);
  assign t[71] = (x[21]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [28:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[29] | t[20]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[31] | t[23]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[13];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[16];
  assign t[41] = t[51] ^ x[22];
  assign t[42] = t[52] ^ x[23];
  assign t[43] = t[53] ^ x[24];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[26];
  assign t[46] = t[56] ^ x[27];
  assign t[47] = t[57] ^ x[28];
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = (~t[60] & t[66]);
  assign t[53] = (~t[60] & t[67]);
  assign t[54] = (~t[64] & t[68]);
  assign t[55] = (~t[64] & t[69]);
  assign t[56] = (~t[60] & t[70]);
  assign t[57] = (~t[64] & t[71]);
  assign t[58] = t[72] ^ x[4];
  assign t[59] = t[73] ^ x[5];
  assign t[5] = ~(~x[2] & ~t[28]);
  assign t[60] = t[74] ^ x[12];
  assign t[61] = t[75] ^ x[13];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[16];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[22];
  assign t[66] = t[80] ^ x[23];
  assign t[67] = t[81] ^ x[24];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[26];
  assign t[6] = ~t[9];
  assign t[70] = t[84] ^ x[27];
  assign t[71] = t[85] ^ x[28];
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[8] & ~x[9] & ~x[10] & ~x[11]) | (~x[8] & x[9] & ~x[10] & ~x[11]) | (~x[8] & ~x[9] & x[10] & ~x[11]) | (~x[8] & ~x[9] & ~x[10] & x[11]) | (x[8] & x[9] & x[10] & ~x[11]) | (x[8] & x[9] & ~x[10] & x[11]) | (x[8] & ~x[9] & x[10] & x[11]) | (~x[8] & x[9] & x[10] & x[11]);
  assign t[75] = (x[9]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[18]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[10]);
  assign t[81] = (x[11]);
  assign t[82] = (x[19]);
  assign t[83] = (x[20]);
  assign t[84] = (x[8]);
  assign t[85] = (x[17]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [50:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[113]);
  assign t[101] = (t[114]);
  assign t[102] = (t[115]);
  assign t[103] = (t[116]);
  assign t[104] = (t[117]);
  assign t[105] = (t[118]);
  assign t[106] = (t[119]);
  assign t[107] = (t[120]);
  assign t[108] = (t[121]);
  assign t[109] = t[122] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[123] ^ x[14];
  assign t[111] = t[124] ^ x[20];
  assign t[112] = t[125] ^ x[26];
  assign t[113] = t[126] ^ x[27];
  assign t[114] = t[127] ^ x[28];
  assign t[115] = t[128] ^ x[29];
  assign t[116] = t[129] ^ x[30];
  assign t[117] = t[130] ^ x[31];
  assign t[118] = t[131] ^ x[32];
  assign t[119] = t[132] ^ x[33];
  assign t[11] = ~x[2] & t[96];
  assign t[120] = t[133] ^ x[34];
  assign t[121] = t[134] ^ x[35];
  assign t[122] = (~t[135] & t[136]);
  assign t[123] = (~t[137] & t[138]);
  assign t[124] = (~t[139] & t[140]);
  assign t[125] = (~t[141] & t[142]);
  assign t[126] = (~t[137] & t[143]);
  assign t[127] = (~t[137] & t[144]);
  assign t[128] = (~t[139] & t[145]);
  assign t[129] = (~t[139] & t[146]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (~t[141] & t[147]);
  assign t[131] = (~t[141] & t[148]);
  assign t[132] = (~t[137] & t[149]);
  assign t[133] = (~t[139] & t[150]);
  assign t[134] = (~t[141] & t[151]);
  assign t[135] = t[152] ^ x[7];
  assign t[136] = t[153] ^ x[8];
  assign t[137] = t[154] ^ x[13];
  assign t[138] = t[155] ^ x[14];
  assign t[139] = t[156] ^ x[19];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[157] ^ x[20];
  assign t[141] = t[158] ^ x[25];
  assign t[142] = t[159] ^ x[26];
  assign t[143] = t[160] ^ x[27];
  assign t[144] = t[161] ^ x[28];
  assign t[145] = t[162] ^ x[29];
  assign t[146] = t[163] ^ x[30];
  assign t[147] = t[164] ^ x[31];
  assign t[148] = t[165] ^ x[32];
  assign t[149] = t[166] ^ x[33];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[167] ^ x[34];
  assign t[151] = t[168] ^ x[35];
  assign t[152] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[6]);
  assign t[154] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[155] = (x[10]);
  assign t[156] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[157] = (x[16]);
  assign t[158] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[159] = (x[22]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[11]);
  assign t[161] = (x[12]);
  assign t[162] = (x[17]);
  assign t[163] = (x[18]);
  assign t[164] = (x[23]);
  assign t[165] = (x[24]);
  assign t[166] = (x[9]);
  assign t[167] = (x[15]);
  assign t[168] = (x[21]);
  assign t[16] = ~(t[97] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[98] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[99] | t[29]);
  assign t[21] = ~(t[100]);
  assign t[22] = ~(t[101]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[103]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[104]);
  assign t[28] = ~(t[105]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[106]);
  assign t[31] = ~(t[100] | t[101]);
  assign t[32] = ~(t[107]);
  assign t[33] = ~(t[102] | t[103]);
  assign t[34] = ~(t[108]);
  assign t[35] = ~(t[104] | t[105]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[37] : x[36];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[38] : t[45];
  assign t[43] = x[2] ? x[39] : t[46];
  assign t[44] = x[2] ? x[40] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[100] & t[22]);
  assign t[49] = ~(t[106] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[102] & t[25]);
  assign t[51] = ~(t[107] & t[55]);
  assign t[52] = ~(t[104] & t[28]);
  assign t[53] = ~(t[108] & t[56]);
  assign t[54] = ~(t[101] & t[21]);
  assign t[55] = ~(t[103] & t[24]);
  assign t[56] = ~(t[105] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[4] ? x[42] : x[41];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[43] : t[66];
  assign t[64] = x[2] ? x[44] : t[67];
  assign t[65] = x[2] ? x[45] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = ~(t[75] & t[97]);
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = ~(t[76] & t[98]);
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = ~(t[77] & t[99]);
  assign t[75] = ~(t[78] & t[21]);
  assign t[76] = ~(t[79] & t[24]);
  assign t[77] = ~(t[80] & t[27]);
  assign t[78] = ~(t[106] & t[101]);
  assign t[79] = ~(t[107] & t[103]);
  assign t[7] = ~(t[11]);
  assign t[80] = ~(t[108] & t[105]);
  assign t[81] = ~(t[82] ^ t[83]);
  assign t[82] = ~t[84];
  assign t[83] = t[4] ? x[47] : x[46];
  assign t[84] = ~(t[85] ^ t[86]);
  assign t[85] = t[87];
  assign t[86] = ~(t[88] ^ t[89]);
  assign t[87] = x[2] ? x[48] : t[90];
  assign t[88] = x[2] ? x[49] : t[91];
  assign t[89] = x[2] ? x[50] : t[92];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = ~(t[69] & t[93]);
  assign t[91] = ~(t[71] & t[94]);
  assign t[92] = ~(t[73] & t[95]);
  assign t[93] = t[15] | t[97];
  assign t[94] = t[17] | t[98];
  assign t[95] = t[19] | t[99];
  assign t[96] = (t[109]);
  assign t[97] = (t[110]);
  assign t[98] = (t[111]);
  assign t[99] = (t[112]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57] & ~t[81]) | (~t[0] & t[36] & ~t[57] & ~t[81]) | (~t[0] & ~t[36] & t[57] & ~t[81]) | (~t[0] & ~t[36] & ~t[57] & t[81]) | (t[0] & t[36] & t[57] & ~t[81]) | (t[0] & t[36] & ~t[57] & t[81]) | (t[0] & ~t[36] & t[57] & t[81]) | (~t[0] & t[36] & t[57] & t[81]);
endmodule

module R2ind116(x, y);
 input [35:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[24]);
  assign t[102] = (x[21]);
  assign t[103] = (x[11]);
  assign t[104] = (x[17]);
  assign t[105] = (x[23]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[33];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[14];
  assign t[48] = t[61] ^ x[20];
  assign t[49] = t[62] ^ x[26];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[27];
  assign t[51] = t[64] ^ x[28];
  assign t[52] = t[65] ^ x[29];
  assign t[53] = t[66] ^ x[30];
  assign t[54] = t[67] ^ x[31];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[33];
  assign t[57] = t[70] ^ x[34];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = (~t[72] & t[73]);
  assign t[5] = t[8];
  assign t[60] = (~t[74] & t[75]);
  assign t[61] = (~t[76] & t[77]);
  assign t[62] = (~t[78] & t[79]);
  assign t[63] = (~t[74] & t[80]);
  assign t[64] = (~t[74] & t[81]);
  assign t[65] = (~t[76] & t[82]);
  assign t[66] = (~t[76] & t[83]);
  assign t[67] = (~t[78] & t[84]);
  assign t[68] = (~t[78] & t[85]);
  assign t[69] = (~t[74] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[76] & t[87]);
  assign t[71] = (~t[78] & t[88]);
  assign t[72] = t[89] ^ x[7];
  assign t[73] = t[90] ^ x[8];
  assign t[74] = t[91] ^ x[13];
  assign t[75] = t[92] ^ x[14];
  assign t[76] = t[93] ^ x[19];
  assign t[77] = t[94] ^ x[20];
  assign t[78] = t[95] ^ x[25];
  assign t[79] = t[96] ^ x[26];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[27];
  assign t[81] = t[98] ^ x[28];
  assign t[82] = t[99] ^ x[29];
  assign t[83] = t[100] ^ x[30];
  assign t[84] = t[101] ^ x[31];
  assign t[85] = t[102] ^ x[32];
  assign t[86] = t[103] ^ x[33];
  assign t[87] = t[104] ^ x[34];
  assign t[88] = t[105] ^ x[35];
  assign t[89] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[6]);
  assign t[91] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[92] = (x[10]);
  assign t[93] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[94] = (x[16]);
  assign t[95] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[96] = (x[22]);
  assign t[97] = (x[12]);
  assign t[98] = (x[9]);
  assign t[99] = (x[18]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [35:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[12]);
  assign t[101] = (x[9]);
  assign t[102] = (x[18]);
  assign t[103] = (x[15]);
  assign t[104] = (x[24]);
  assign t[105] = (x[21]);
  assign t[106] = (x[11]);
  assign t[107] = (x[17]);
  assign t[108] = (x[23]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[36];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[38]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[45] & t[44]);
  assign t[35] = ~(t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[28];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[34];
  assign t[61] = t[74] ^ x[35];
  assign t[62] = (~t[75] & t[76]);
  assign t[63] = (~t[77] & t[78]);
  assign t[64] = (~t[79] & t[80]);
  assign t[65] = (~t[81] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[81] & t[87]);
  assign t[71] = (~t[81] & t[88]);
  assign t[72] = (~t[77] & t[89]);
  assign t[73] = (~t[79] & t[90]);
  assign t[74] = (~t[81] & t[91]);
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[8];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[19];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[25];
  assign t[82] = t[99] ^ x[26];
  assign t[83] = t[100] ^ x[27];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = t[108] ^ x[35];
  assign t[92] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[6]);
  assign t[94] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[95] = (x[10]);
  assign t[96] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[97] = (x[16]);
  assign t[98] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[99] = (x[22]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [32:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[14];
  assign t[42] = t[52] ^ x[15];
  assign t[43] = t[53] ^ x[21];
  assign t[44] = t[54] ^ x[22];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[29];
  assign t[47] = t[57] ^ x[30];
  assign t[48] = t[58] ^ x[31];
  assign t[49] = t[59] ^ x[32];
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[62] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = (~t[65] & t[67]);
  assign t[55] = (~t[68] & t[69]);
  assign t[56] = (~t[68] & t[70]);
  assign t[57] = (~t[62] & t[71]);
  assign t[58] = (~t[65] & t[72]);
  assign t[59] = (~t[68] & t[73]);
  assign t[5] = t[8];
  assign t[60] = t[74] ^ x[7];
  assign t[61] = t[75] ^ x[8];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[15];
  assign t[65] = t[79] ^ x[20];
  assign t[66] = t[80] ^ x[21];
  assign t[67] = t[81] ^ x[22];
  assign t[68] = t[82] ^ x[27];
  assign t[69] = t[83] ^ x[28];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[84] ^ x[29];
  assign t[71] = t[85] ^ x[30];
  assign t[72] = t[86] ^ x[31];
  assign t[73] = t[87] ^ x[32];
  assign t[74] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[6]);
  assign t[76] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[77] = (x[11]);
  assign t[78] = (x[9]);
  assign t[79] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[18]);
  assign t[81] = (x[16]);
  assign t[82] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[83] = (x[25]);
  assign t[84] = (x[23]);
  assign t[85] = (x[12]);
  assign t[86] = (x[19]);
  assign t[87] = (x[26]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [35:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[11]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[18]);
  assign t[104] = (x[23]);
  assign t[105] = (x[24]);
  assign t[106] = (x[9]);
  assign t[107] = (x[15]);
  assign t[108] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[36];
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[28];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[34];
  assign t[61] = t[74] ^ x[35];
  assign t[62] = (~t[75] & t[76]);
  assign t[63] = (~t[77] & t[78]);
  assign t[64] = (~t[79] & t[80]);
  assign t[65] = (~t[81] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[81] & t[87]);
  assign t[71] = (~t[81] & t[88]);
  assign t[72] = (~t[77] & t[89]);
  assign t[73] = (~t[79] & t[90]);
  assign t[74] = (~t[81] & t[91]);
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[8];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[19];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[25];
  assign t[82] = t[99] ^ x[26];
  assign t[83] = t[100] ^ x[27];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = t[108] ^ x[35];
  assign t[92] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[6]);
  assign t[94] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[95] = (x[10]);
  assign t[96] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[97] = (x[16]);
  assign t[98] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[99] = (x[22]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [50:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[113]);
  assign t[101] = (t[114]);
  assign t[102] = (t[115]);
  assign t[103] = (t[116]);
  assign t[104] = (t[117]);
  assign t[105] = (t[118]);
  assign t[106] = (t[119]);
  assign t[107] = (t[120]);
  assign t[108] = (t[121]);
  assign t[109] = t[122] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[123] ^ x[14];
  assign t[111] = t[124] ^ x[20];
  assign t[112] = t[125] ^ x[26];
  assign t[113] = t[126] ^ x[27];
  assign t[114] = t[127] ^ x[28];
  assign t[115] = t[128] ^ x[29];
  assign t[116] = t[129] ^ x[30];
  assign t[117] = t[130] ^ x[31];
  assign t[118] = t[131] ^ x[32];
  assign t[119] = t[132] ^ x[33];
  assign t[11] = ~x[2] & t[96];
  assign t[120] = t[133] ^ x[34];
  assign t[121] = t[134] ^ x[35];
  assign t[122] = (~t[135] & t[136]);
  assign t[123] = (~t[137] & t[138]);
  assign t[124] = (~t[139] & t[140]);
  assign t[125] = (~t[141] & t[142]);
  assign t[126] = (~t[137] & t[143]);
  assign t[127] = (~t[137] & t[144]);
  assign t[128] = (~t[139] & t[145]);
  assign t[129] = (~t[139] & t[146]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (~t[141] & t[147]);
  assign t[131] = (~t[141] & t[148]);
  assign t[132] = (~t[137] & t[149]);
  assign t[133] = (~t[139] & t[150]);
  assign t[134] = (~t[141] & t[151]);
  assign t[135] = t[152] ^ x[7];
  assign t[136] = t[153] ^ x[8];
  assign t[137] = t[154] ^ x[13];
  assign t[138] = t[155] ^ x[14];
  assign t[139] = t[156] ^ x[19];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[157] ^ x[20];
  assign t[141] = t[158] ^ x[25];
  assign t[142] = t[159] ^ x[26];
  assign t[143] = t[160] ^ x[27];
  assign t[144] = t[161] ^ x[28];
  assign t[145] = t[162] ^ x[29];
  assign t[146] = t[163] ^ x[30];
  assign t[147] = t[164] ^ x[31];
  assign t[148] = t[165] ^ x[32];
  assign t[149] = t[166] ^ x[33];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[167] ^ x[34];
  assign t[151] = t[168] ^ x[35];
  assign t[152] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[6]);
  assign t[154] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[155] = (x[10]);
  assign t[156] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[157] = (x[16]);
  assign t[158] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[159] = (x[22]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[11]);
  assign t[161] = (x[12]);
  assign t[162] = (x[17]);
  assign t[163] = (x[18]);
  assign t[164] = (x[23]);
  assign t[165] = (x[24]);
  assign t[166] = (x[9]);
  assign t[167] = (x[15]);
  assign t[168] = (x[21]);
  assign t[16] = ~(t[97] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[98] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[99] | t[29]);
  assign t[21] = ~(t[100]);
  assign t[22] = ~(t[101]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[103]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[104]);
  assign t[28] = ~(t[105]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[106]);
  assign t[31] = ~(t[100] | t[101]);
  assign t[32] = ~(t[107]);
  assign t[33] = ~(t[102] | t[103]);
  assign t[34] = ~(t[108]);
  assign t[35] = ~(t[104] | t[105]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[11] ? x[37] : x[36];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[38] : t[45];
  assign t[43] = x[2] ? x[39] : t[46];
  assign t[44] = x[2] ? x[40] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[100] & t[22]);
  assign t[49] = ~(t[106] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[102] & t[25]);
  assign t[51] = ~(t[107] & t[55]);
  assign t[52] = ~(t[104] & t[28]);
  assign t[53] = ~(t[108] & t[56]);
  assign t[54] = ~(t[101] & t[21]);
  assign t[55] = ~(t[103] & t[24]);
  assign t[56] = ~(t[105] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[11] ? x[42] : x[41];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[43] : t[66];
  assign t[64] = x[2] ? x[44] : t[67];
  assign t[65] = x[2] ? x[45] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = ~(t[75] & t[97]);
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = ~(t[76] & t[98]);
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = ~(t[77] & t[99]);
  assign t[75] = ~(t[78] & t[21]);
  assign t[76] = ~(t[79] & t[24]);
  assign t[77] = ~(t[80] & t[27]);
  assign t[78] = ~(t[106] & t[101]);
  assign t[79] = ~(t[107] & t[103]);
  assign t[7] = ~(t[11]);
  assign t[80] = ~(t[108] & t[105]);
  assign t[81] = ~(t[82] ^ t[83]);
  assign t[82] = ~t[84];
  assign t[83] = t[4] ? x[47] : x[46];
  assign t[84] = ~(t[85] ^ t[86]);
  assign t[85] = t[87];
  assign t[86] = ~(t[88] ^ t[89]);
  assign t[87] = x[2] ? x[48] : t[90];
  assign t[88] = x[2] ? x[49] : t[91];
  assign t[89] = x[2] ? x[50] : t[92];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = ~(t[69] & t[93]);
  assign t[91] = ~(t[71] & t[94]);
  assign t[92] = ~(t[73] & t[95]);
  assign t[93] = t[15] | t[97];
  assign t[94] = t[17] | t[98];
  assign t[95] = t[19] | t[99];
  assign t[96] = (t[109]);
  assign t[97] = (t[110]);
  assign t[98] = (t[111]);
  assign t[99] = (t[112]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57] & ~t[81]) | (~t[0] & t[36] & ~t[57] & ~t[81]) | (~t[0] & ~t[36] & t[57] & ~t[81]) | (~t[0] & ~t[36] & ~t[57] & t[81]) | (t[0] & t[36] & t[57] & ~t[81]) | (t[0] & t[36] & ~t[57] & t[81]) | (t[0] & ~t[36] & t[57] & t[81]) | (~t[0] & t[36] & t[57] & t[81]);
endmodule

module R2ind121(x, y);
 input [35:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[24]);
  assign t[102] = (x[21]);
  assign t[103] = (x[11]);
  assign t[104] = (x[17]);
  assign t[105] = (x[23]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[33];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[14];
  assign t[48] = t[61] ^ x[20];
  assign t[49] = t[62] ^ x[26];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[27];
  assign t[51] = t[64] ^ x[28];
  assign t[52] = t[65] ^ x[29];
  assign t[53] = t[66] ^ x[30];
  assign t[54] = t[67] ^ x[31];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[33];
  assign t[57] = t[70] ^ x[34];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = (~t[72] & t[73]);
  assign t[5] = t[8];
  assign t[60] = (~t[74] & t[75]);
  assign t[61] = (~t[76] & t[77]);
  assign t[62] = (~t[78] & t[79]);
  assign t[63] = (~t[74] & t[80]);
  assign t[64] = (~t[74] & t[81]);
  assign t[65] = (~t[76] & t[82]);
  assign t[66] = (~t[76] & t[83]);
  assign t[67] = (~t[78] & t[84]);
  assign t[68] = (~t[78] & t[85]);
  assign t[69] = (~t[74] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[76] & t[87]);
  assign t[71] = (~t[78] & t[88]);
  assign t[72] = t[89] ^ x[7];
  assign t[73] = t[90] ^ x[8];
  assign t[74] = t[91] ^ x[13];
  assign t[75] = t[92] ^ x[14];
  assign t[76] = t[93] ^ x[19];
  assign t[77] = t[94] ^ x[20];
  assign t[78] = t[95] ^ x[25];
  assign t[79] = t[96] ^ x[26];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[27];
  assign t[81] = t[98] ^ x[28];
  assign t[82] = t[99] ^ x[29];
  assign t[83] = t[100] ^ x[30];
  assign t[84] = t[101] ^ x[31];
  assign t[85] = t[102] ^ x[32];
  assign t[86] = t[103] ^ x[33];
  assign t[87] = t[104] ^ x[34];
  assign t[88] = t[105] ^ x[35];
  assign t[89] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[6]);
  assign t[91] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[92] = (x[10]);
  assign t[93] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[94] = (x[16]);
  assign t[95] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[96] = (x[22]);
  assign t[97] = (x[12]);
  assign t[98] = (x[9]);
  assign t[99] = (x[18]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [35:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[18]);
  assign t[101] = (x[15]);
  assign t[102] = (x[24]);
  assign t[103] = (x[21]);
  assign t[104] = (x[11]);
  assign t[105] = (x[17]);
  assign t[106] = (x[23]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = ~(t[21] & t[35]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[36]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[39] & t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[20];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[26];
  assign t[51] = t[64] ^ x[27];
  assign t[52] = t[65] ^ x[28];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[30];
  assign t[55] = t[68] ^ x[31];
  assign t[56] = t[69] ^ x[32];
  assign t[57] = t[70] ^ x[33];
  assign t[58] = t[71] ^ x[34];
  assign t[59] = t[72] ^ x[35];
  assign t[5] = t[7];
  assign t[60] = (~t[73] & t[74]);
  assign t[61] = (~t[75] & t[76]);
  assign t[62] = (~t[77] & t[78]);
  assign t[63] = (~t[79] & t[80]);
  assign t[64] = (~t[75] & t[81]);
  assign t[65] = (~t[75] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (~t[75] & t[87]);
  assign t[71] = (~t[77] & t[88]);
  assign t[72] = (~t[79] & t[89]);
  assign t[73] = t[90] ^ x[4];
  assign t[74] = t[91] ^ x[5];
  assign t[75] = t[92] ^ x[13];
  assign t[76] = t[93] ^ x[14];
  assign t[77] = t[94] ^ x[19];
  assign t[78] = t[95] ^ x[20];
  assign t[79] = t[96] ^ x[25];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[97] ^ x[26];
  assign t[81] = t[98] ^ x[27];
  assign t[82] = t[99] ^ x[28];
  assign t[83] = t[100] ^ x[29];
  assign t[84] = t[101] ^ x[30];
  assign t[85] = t[102] ^ x[31];
  assign t[86] = t[103] ^ x[32];
  assign t[87] = t[104] ^ x[33];
  assign t[88] = t[105] ^ x[34];
  assign t[89] = t[106] ^ x[35];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[3]);
  assign t[92] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[93] = (x[10]);
  assign t[94] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[95] = (x[16]);
  assign t[96] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[97] = (x[22]);
  assign t[98] = (x[12]);
  assign t[99] = (x[9]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [32:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[29] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[35] & t[25]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[36] & t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = ~(t[37] & t[27]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[31]);
  assign t[27] = ~(t[33]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[14];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[15];
  assign t[41] = t[51] ^ x[21];
  assign t[42] = t[52] ^ x[22];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[29];
  assign t[45] = t[55] ^ x[30];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[32];
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~x[2] & t[28];
  assign t[50] = (~t[60] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[63] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[66] & t[68]);
  assign t[55] = (~t[60] & t[69]);
  assign t[56] = (~t[63] & t[70]);
  assign t[57] = (~t[66] & t[71]);
  assign t[58] = t[72] ^ x[4];
  assign t[59] = t[73] ^ x[5];
  assign t[5] = t[7];
  assign t[60] = t[74] ^ x[13];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[20];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[22];
  assign t[66] = t[80] ^ x[27];
  assign t[67] = t[81] ^ x[28];
  assign t[68] = t[82] ^ x[29];
  assign t[69] = t[83] ^ x[30];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[84] ^ x[31];
  assign t[71] = t[85] ^ x[32];
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[75] = (x[11]);
  assign t[76] = (x[9]);
  assign t[77] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[78] = (x[18]);
  assign t[79] = (x[16]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[81] = (x[25]);
  assign t[82] = (x[23]);
  assign t[83] = (x[12]);
  assign t[84] = (x[19]);
  assign t[85] = (x[26]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [35:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[11]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[18]);
  assign t[104] = (x[23]);
  assign t[105] = (x[24]);
  assign t[106] = (x[9]);
  assign t[107] = (x[15]);
  assign t[108] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[36];
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[28];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[34];
  assign t[61] = t[74] ^ x[35];
  assign t[62] = (~t[75] & t[76]);
  assign t[63] = (~t[77] & t[78]);
  assign t[64] = (~t[79] & t[80]);
  assign t[65] = (~t[81] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[81] & t[87]);
  assign t[71] = (~t[81] & t[88]);
  assign t[72] = (~t[77] & t[89]);
  assign t[73] = (~t[79] & t[90]);
  assign t[74] = (~t[81] & t[91]);
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[8];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[19];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[25];
  assign t[82] = t[99] ^ x[26];
  assign t[83] = t[100] ^ x[27];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = t[108] ^ x[35];
  assign t[92] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[6]);
  assign t[94] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[95] = (x[10]);
  assign t[96] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[97] = (x[16]);
  assign t[98] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[99] = (x[22]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [50:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[113]);
  assign t[101] = (t[114]);
  assign t[102] = (t[115]);
  assign t[103] = (t[116]);
  assign t[104] = (t[117]);
  assign t[105] = (t[118]);
  assign t[106] = (t[119]);
  assign t[107] = (t[120]);
  assign t[108] = (t[121]);
  assign t[109] = t[122] ^ x[5];
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = t[123] ^ x[14];
  assign t[111] = t[124] ^ x[20];
  assign t[112] = t[125] ^ x[26];
  assign t[113] = t[126] ^ x[27];
  assign t[114] = t[127] ^ x[28];
  assign t[115] = t[128] ^ x[29];
  assign t[116] = t[129] ^ x[30];
  assign t[117] = t[130] ^ x[31];
  assign t[118] = t[131] ^ x[32];
  assign t[119] = t[132] ^ x[33];
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = t[133] ^ x[34];
  assign t[121] = t[134] ^ x[35];
  assign t[122] = (~t[135] & t[136]);
  assign t[123] = (~t[137] & t[138]);
  assign t[124] = (~t[139] & t[140]);
  assign t[125] = (~t[141] & t[142]);
  assign t[126] = (~t[137] & t[143]);
  assign t[127] = (~t[137] & t[144]);
  assign t[128] = (~t[139] & t[145]);
  assign t[129] = (~t[139] & t[146]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[130] = (~t[141] & t[147]);
  assign t[131] = (~t[141] & t[148]);
  assign t[132] = (~t[137] & t[149]);
  assign t[133] = (~t[139] & t[150]);
  assign t[134] = (~t[141] & t[151]);
  assign t[135] = t[152] ^ x[4];
  assign t[136] = t[153] ^ x[5];
  assign t[137] = t[154] ^ x[13];
  assign t[138] = t[155] ^ x[14];
  assign t[139] = t[156] ^ x[19];
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = t[157] ^ x[20];
  assign t[141] = t[158] ^ x[25];
  assign t[142] = t[159] ^ x[26];
  assign t[143] = t[160] ^ x[27];
  assign t[144] = t[161] ^ x[28];
  assign t[145] = t[162] ^ x[29];
  assign t[146] = t[163] ^ x[30];
  assign t[147] = t[164] ^ x[31];
  assign t[148] = t[165] ^ x[32];
  assign t[149] = t[166] ^ x[33];
  assign t[14] = ~(t[97] | t[21]);
  assign t[150] = t[167] ^ x[34];
  assign t[151] = t[168] ^ x[35];
  assign t[152] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[3]);
  assign t[154] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[155] = (x[10]);
  assign t[156] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[157] = (x[16]);
  assign t[158] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[159] = (x[22]);
  assign t[15] = ~(t[22] | t[23]);
  assign t[160] = (x[11]);
  assign t[161] = (x[12]);
  assign t[162] = (x[17]);
  assign t[163] = (x[18]);
  assign t[164] = (x[23]);
  assign t[165] = (x[24]);
  assign t[166] = (x[9]);
  assign t[167] = (x[15]);
  assign t[168] = (x[21]);
  assign t[16] = ~(t[98] | t[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[18] = ~(t[99] | t[27]);
  assign t[19] = ~(t[100]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[101]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[102]);
  assign t[23] = ~(t[103]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[104]);
  assign t[26] = ~(t[105]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[106]);
  assign t[29] = ~(t[100] | t[101]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[107]);
  assign t[31] = ~(t[102] | t[103]);
  assign t[32] = ~(t[108]);
  assign t[33] = ~(t[104] | t[105]);
  assign t[34] = ~(t[35] ^ t[36]);
  assign t[35] = ~t[37];
  assign t[36] = t[38] ? x[37] : x[36];
  assign t[37] = ~(t[39] ^ t[40]);
  assign t[38] = ~(t[41]);
  assign t[39] = t[42];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[43] ^ t[44]);
  assign t[41] = ~(t[4]);
  assign t[42] = x[2] ? x[38] : t[45];
  assign t[43] = x[2] ? x[39] : t[46];
  assign t[44] = x[2] ? x[40] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[100] & t[20]);
  assign t[49] = ~(t[106] & t[54]);
  assign t[4] = ~x[2] & t[96];
  assign t[50] = ~(t[102] & t[23]);
  assign t[51] = ~(t[107] & t[55]);
  assign t[52] = ~(t[104] & t[26]);
  assign t[53] = ~(t[108] & t[56]);
  assign t[54] = ~(t[101] & t[19]);
  assign t[55] = ~(t[103] & t[22]);
  assign t[56] = ~(t[105] & t[25]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[38] ? x[42] : x[41];
  assign t[5] = t[7];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[43] : t[66];
  assign t[64] = x[2] ? x[44] : t[67];
  assign t[65] = x[2] ? x[45] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[20] & t[28]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = ~(t[75] & t[97]);
  assign t[71] = ~(t[23] & t[30]);
  assign t[72] = ~(t[76] & t[98]);
  assign t[73] = ~(t[26] & t[32]);
  assign t[74] = ~(t[77] & t[99]);
  assign t[75] = ~(t[78] & t[19]);
  assign t[76] = ~(t[79] & t[22]);
  assign t[77] = ~(t[80] & t[25]);
  assign t[78] = ~(t[106] & t[101]);
  assign t[79] = ~(t[107] & t[103]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = ~(t[108] & t[105]);
  assign t[81] = ~(t[82] ^ t[83]);
  assign t[82] = ~t[84];
  assign t[83] = t[4] ? x[47] : x[46];
  assign t[84] = ~(t[85] ^ t[86]);
  assign t[85] = t[87];
  assign t[86] = ~(t[88] ^ t[89]);
  assign t[87] = x[2] ? x[48] : t[90];
  assign t[88] = x[2] ? x[49] : t[91];
  assign t[89] = x[2] ? x[50] : t[92];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = ~(t[69] & t[93]);
  assign t[91] = ~(t[71] & t[94]);
  assign t[92] = ~(t[73] & t[95]);
  assign t[93] = t[13] | t[97];
  assign t[94] = t[15] | t[98];
  assign t[95] = t[17] | t[99];
  assign t[96] = (t[109]);
  assign t[97] = (t[110]);
  assign t[98] = (t[111]);
  assign t[99] = (t[112]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0] & ~t[34] & ~t[57] & ~t[81]) | (~t[0] & t[34] & ~t[57] & ~t[81]) | (~t[0] & ~t[34] & t[57] & ~t[81]) | (~t[0] & ~t[34] & ~t[57] & t[81]) | (t[0] & t[34] & t[57] & ~t[81]) | (t[0] & t[34] & ~t[57] & t[81]) | (t[0] & ~t[34] & t[57] & t[81]) | (~t[0] & t[34] & t[57] & t[81]);
endmodule

module R2ind126(x, y);
 input [35:0] x;
 output y;

 wire [103:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[21]);
  assign t[101] = (x[11]);
  assign t[102] = (x[17]);
  assign t[103] = (x[23]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = t[21] | t[32];
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = t[24] | t[33];
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] | t[34];
  assign t[19] = ~(t[35]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[28] | t[19]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] | t[22]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[30] | t[25]);
  assign t[28] = ~(t[41]);
  assign t[29] = ~(t[42]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = t[57] ^ x[5];
  assign t[45] = t[58] ^ x[14];
  assign t[46] = t[59] ^ x[20];
  assign t[47] = t[60] ^ x[26];
  assign t[48] = t[61] ^ x[27];
  assign t[49] = t[62] ^ x[28];
  assign t[4] = ~x[2] & t[31];
  assign t[50] = t[63] ^ x[29];
  assign t[51] = t[64] ^ x[30];
  assign t[52] = t[65] ^ x[31];
  assign t[53] = t[66] ^ x[32];
  assign t[54] = t[67] ^ x[33];
  assign t[55] = t[68] ^ x[34];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = (~t[70] & t[71]);
  assign t[58] = (~t[72] & t[73]);
  assign t[59] = (~t[74] & t[75]);
  assign t[5] = t[7];
  assign t[60] = (~t[76] & t[77]);
  assign t[61] = (~t[72] & t[78]);
  assign t[62] = (~t[72] & t[79]);
  assign t[63] = (~t[74] & t[80]);
  assign t[64] = (~t[74] & t[81]);
  assign t[65] = (~t[76] & t[82]);
  assign t[66] = (~t[76] & t[83]);
  assign t[67] = (~t[72] & t[84]);
  assign t[68] = (~t[74] & t[85]);
  assign t[69] = (~t[76] & t[86]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[87] ^ x[4];
  assign t[71] = t[88] ^ x[5];
  assign t[72] = t[89] ^ x[13];
  assign t[73] = t[90] ^ x[14];
  assign t[74] = t[91] ^ x[19];
  assign t[75] = t[92] ^ x[20];
  assign t[76] = t[93] ^ x[25];
  assign t[77] = t[94] ^ x[26];
  assign t[78] = t[95] ^ x[27];
  assign t[79] = t[96] ^ x[28];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[97] ^ x[29];
  assign t[81] = t[98] ^ x[30];
  assign t[82] = t[99] ^ x[31];
  assign t[83] = t[100] ^ x[32];
  assign t[84] = t[101] ^ x[33];
  assign t[85] = t[102] ^ x[34];
  assign t[86] = t[103] ^ x[35];
  assign t[87] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[3]);
  assign t[89] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = (x[10]);
  assign t[91] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[92] = (x[16]);
  assign t[93] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[94] = (x[22]);
  assign t[95] = (x[12]);
  assign t[96] = (x[9]);
  assign t[97] = (x[18]);
  assign t[98] = (x[15]);
  assign t[99] = (x[24]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [35:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[12]);
  assign t[101] = (x[9]);
  assign t[102] = (x[18]);
  assign t[103] = (x[15]);
  assign t[104] = (x[24]);
  assign t[105] = (x[21]);
  assign t[106] = (x[11]);
  assign t[107] = (x[17]);
  assign t[108] = (x[23]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[36];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[38]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[45] & t[44]);
  assign t[35] = ~(t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[28];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[34];
  assign t[61] = t[74] ^ x[35];
  assign t[62] = (~t[75] & t[76]);
  assign t[63] = (~t[77] & t[78]);
  assign t[64] = (~t[79] & t[80]);
  assign t[65] = (~t[81] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[81] & t[87]);
  assign t[71] = (~t[81] & t[88]);
  assign t[72] = (~t[77] & t[89]);
  assign t[73] = (~t[79] & t[90]);
  assign t[74] = (~t[81] & t[91]);
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[8];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[19];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[25];
  assign t[82] = t[99] ^ x[26];
  assign t[83] = t[100] ^ x[27];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = t[108] ^ x[35];
  assign t[92] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[6]);
  assign t[94] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[95] = (x[10]);
  assign t[96] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[97] = (x[16]);
  assign t[98] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[99] = (x[22]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [32:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[14];
  assign t[42] = t[52] ^ x[15];
  assign t[43] = t[53] ^ x[21];
  assign t[44] = t[54] ^ x[22];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[29];
  assign t[47] = t[57] ^ x[30];
  assign t[48] = t[58] ^ x[31];
  assign t[49] = t[59] ^ x[32];
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[62] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = (~t[65] & t[67]);
  assign t[55] = (~t[68] & t[69]);
  assign t[56] = (~t[68] & t[70]);
  assign t[57] = (~t[62] & t[71]);
  assign t[58] = (~t[65] & t[72]);
  assign t[59] = (~t[68] & t[73]);
  assign t[5] = t[8];
  assign t[60] = t[74] ^ x[7];
  assign t[61] = t[75] ^ x[8];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[15];
  assign t[65] = t[79] ^ x[20];
  assign t[66] = t[80] ^ x[21];
  assign t[67] = t[81] ^ x[22];
  assign t[68] = t[82] ^ x[27];
  assign t[69] = t[83] ^ x[28];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[84] ^ x[29];
  assign t[71] = t[85] ^ x[30];
  assign t[72] = t[86] ^ x[31];
  assign t[73] = t[87] ^ x[32];
  assign t[74] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[6]);
  assign t[76] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[77] = (x[11]);
  assign t[78] = (x[9]);
  assign t[79] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[18]);
  assign t[81] = (x[16]);
  assign t[82] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[83] = (x[25]);
  assign t[84] = (x[23]);
  assign t[85] = (x[12]);
  assign t[86] = (x[19]);
  assign t[87] = (x[26]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [35:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[17]);
  assign t[101] = (x[18]);
  assign t[102] = (x[23]);
  assign t[103] = (x[24]);
  assign t[104] = (x[9]);
  assign t[105] = (x[15]);
  assign t[106] = (x[21]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[14] = ~(t[35] | t[21]);
  assign t[15] = ~(t[22] | t[23]);
  assign t[16] = ~(t[36] | t[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[18] = ~(t[37] | t[27]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[44]);
  assign t[29] = ~(t[38] | t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[20];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[26];
  assign t[51] = t[64] ^ x[27];
  assign t[52] = t[65] ^ x[28];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[30];
  assign t[55] = t[68] ^ x[31];
  assign t[56] = t[69] ^ x[32];
  assign t[57] = t[70] ^ x[33];
  assign t[58] = t[71] ^ x[34];
  assign t[59] = t[72] ^ x[35];
  assign t[5] = t[7];
  assign t[60] = (~t[73] & t[74]);
  assign t[61] = (~t[75] & t[76]);
  assign t[62] = (~t[77] & t[78]);
  assign t[63] = (~t[79] & t[80]);
  assign t[64] = (~t[75] & t[81]);
  assign t[65] = (~t[75] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (~t[75] & t[87]);
  assign t[71] = (~t[77] & t[88]);
  assign t[72] = (~t[79] & t[89]);
  assign t[73] = t[90] ^ x[4];
  assign t[74] = t[91] ^ x[5];
  assign t[75] = t[92] ^ x[13];
  assign t[76] = t[93] ^ x[14];
  assign t[77] = t[94] ^ x[19];
  assign t[78] = t[95] ^ x[20];
  assign t[79] = t[96] ^ x[25];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[97] ^ x[26];
  assign t[81] = t[98] ^ x[27];
  assign t[82] = t[99] ^ x[28];
  assign t[83] = t[100] ^ x[29];
  assign t[84] = t[101] ^ x[30];
  assign t[85] = t[102] ^ x[31];
  assign t[86] = t[103] ^ x[32];
  assign t[87] = t[104] ^ x[33];
  assign t[88] = t[105] ^ x[34];
  assign t[89] = t[106] ^ x[35];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[3]);
  assign t[92] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[93] = (x[10]);
  assign t[94] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[95] = (x[16]);
  assign t[96] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[97] = (x[22]);
  assign t[98] = (x[11]);
  assign t[99] = (x[12]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [50:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (t[113]);
  assign t[101] = (t[114]);
  assign t[102] = (t[115]);
  assign t[103] = (t[116]);
  assign t[104] = (t[117]);
  assign t[105] = (t[118]);
  assign t[106] = (t[119]);
  assign t[107] = (t[120]);
  assign t[108] = (t[121]);
  assign t[109] = t[122] ^ x[8];
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = t[123] ^ x[14];
  assign t[111] = t[124] ^ x[20];
  assign t[112] = t[125] ^ x[26];
  assign t[113] = t[126] ^ x[27];
  assign t[114] = t[127] ^ x[28];
  assign t[115] = t[128] ^ x[29];
  assign t[116] = t[129] ^ x[30];
  assign t[117] = t[130] ^ x[31];
  assign t[118] = t[131] ^ x[32];
  assign t[119] = t[132] ^ x[33];
  assign t[11] = ~x[2] & t[96];
  assign t[120] = t[133] ^ x[34];
  assign t[121] = t[134] ^ x[35];
  assign t[122] = (~t[135] & t[136]);
  assign t[123] = (~t[137] & t[138]);
  assign t[124] = (~t[139] & t[140]);
  assign t[125] = (~t[141] & t[142]);
  assign t[126] = (~t[137] & t[143]);
  assign t[127] = (~t[137] & t[144]);
  assign t[128] = (~t[139] & t[145]);
  assign t[129] = (~t[139] & t[146]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (~t[141] & t[147]);
  assign t[131] = (~t[141] & t[148]);
  assign t[132] = (~t[137] & t[149]);
  assign t[133] = (~t[139] & t[150]);
  assign t[134] = (~t[141] & t[151]);
  assign t[135] = t[152] ^ x[7];
  assign t[136] = t[153] ^ x[8];
  assign t[137] = t[154] ^ x[13];
  assign t[138] = t[155] ^ x[14];
  assign t[139] = t[156] ^ x[19];
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = t[157] ^ x[20];
  assign t[141] = t[158] ^ x[25];
  assign t[142] = t[159] ^ x[26];
  assign t[143] = t[160] ^ x[27];
  assign t[144] = t[161] ^ x[28];
  assign t[145] = t[162] ^ x[29];
  assign t[146] = t[163] ^ x[30];
  assign t[147] = t[164] ^ x[31];
  assign t[148] = t[165] ^ x[32];
  assign t[149] = t[166] ^ x[33];
  assign t[14] = ~(t[19] | t[20]);
  assign t[150] = t[167] ^ x[34];
  assign t[151] = t[168] ^ x[35];
  assign t[152] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[6]);
  assign t[154] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[155] = (x[10]);
  assign t[156] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[157] = (x[16]);
  assign t[158] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[159] = (x[22]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (x[11]);
  assign t[161] = (x[12]);
  assign t[162] = (x[17]);
  assign t[163] = (x[18]);
  assign t[164] = (x[23]);
  assign t[165] = (x[24]);
  assign t[166] = (x[9]);
  assign t[167] = (x[15]);
  assign t[168] = (x[21]);
  assign t[16] = ~(t[97] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[98] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[99] | t[29]);
  assign t[21] = ~(t[100]);
  assign t[22] = ~(t[101]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[103]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[104]);
  assign t[28] = ~(t[105]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[106]);
  assign t[31] = ~(t[100] | t[101]);
  assign t[32] = ~(t[107]);
  assign t[33] = ~(t[102] | t[103]);
  assign t[34] = ~(t[108]);
  assign t[35] = ~(t[104] | t[105]);
  assign t[36] = ~(t[37] ^ t[38]);
  assign t[37] = ~t[39];
  assign t[38] = t[4] ? x[37] : x[36];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[42];
  assign t[41] = ~(t[43] ^ t[44]);
  assign t[42] = x[2] ? x[38] : t[45];
  assign t[43] = x[2] ? x[39] : t[46];
  assign t[44] = x[2] ? x[40] : t[47];
  assign t[45] = ~(t[48] & t[49]);
  assign t[46] = ~(t[50] & t[51]);
  assign t[47] = ~(t[52] & t[53]);
  assign t[48] = ~(t[100] & t[22]);
  assign t[49] = ~(t[106] & t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = ~(t[102] & t[25]);
  assign t[51] = ~(t[107] & t[55]);
  assign t[52] = ~(t[104] & t[28]);
  assign t[53] = ~(t[108] & t[56]);
  assign t[54] = ~(t[101] & t[21]);
  assign t[55] = ~(t[103] & t[24]);
  assign t[56] = ~(t[105] & t[27]);
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = t[11] ? x[42] : x[41];
  assign t[5] = t[8];
  assign t[60] = ~(t[61] ^ t[62]);
  assign t[61] = t[63];
  assign t[62] = ~(t[64] ^ t[65]);
  assign t[63] = x[2] ? x[43] : t[66];
  assign t[64] = x[2] ? x[44] : t[67];
  assign t[65] = x[2] ? x[45] : t[68];
  assign t[66] = ~(t[69] & t[70]);
  assign t[67] = ~(t[71] & t[72]);
  assign t[68] = ~(t[73] & t[74]);
  assign t[69] = ~(t[22] & t[30]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = ~(t[75] & t[97]);
  assign t[71] = ~(t[25] & t[32]);
  assign t[72] = ~(t[76] & t[98]);
  assign t[73] = ~(t[28] & t[34]);
  assign t[74] = ~(t[77] & t[99]);
  assign t[75] = ~(t[78] & t[21]);
  assign t[76] = ~(t[79] & t[24]);
  assign t[77] = ~(t[80] & t[27]);
  assign t[78] = ~(t[106] & t[101]);
  assign t[79] = ~(t[107] & t[103]);
  assign t[7] = ~(t[11]);
  assign t[80] = ~(t[108] & t[105]);
  assign t[81] = ~(t[82] ^ t[83]);
  assign t[82] = ~t[84];
  assign t[83] = t[4] ? x[47] : x[46];
  assign t[84] = ~(t[85] ^ t[86]);
  assign t[85] = t[87];
  assign t[86] = ~(t[88] ^ t[89]);
  assign t[87] = x[2] ? x[48] : t[90];
  assign t[88] = x[2] ? x[49] : t[91];
  assign t[89] = x[2] ? x[50] : t[92];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = ~(t[69] & t[93]);
  assign t[91] = ~(t[71] & t[94]);
  assign t[92] = ~(t[73] & t[95]);
  assign t[93] = t[15] | t[97];
  assign t[94] = t[17] | t[98];
  assign t[95] = t[19] | t[99];
  assign t[96] = (t[109]);
  assign t[97] = (t[110]);
  assign t[98] = (t[111]);
  assign t[99] = (t[112]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0] & ~t[36] & ~t[57] & ~t[81]) | (~t[0] & t[36] & ~t[57] & ~t[81]) | (~t[0] & ~t[36] & t[57] & ~t[81]) | (~t[0] & ~t[36] & ~t[57] & t[81]) | (t[0] & t[36] & t[57] & ~t[81]) | (t[0] & t[36] & ~t[57] & t[81]) | (t[0] & ~t[36] & t[57] & t[81]) | (~t[0] & t[36] & t[57] & t[81]);
endmodule

module R2ind131(x, y);
 input [35:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[24]);
  assign t[102] = (x[21]);
  assign t[103] = (x[11]);
  assign t[104] = (x[17]);
  assign t[105] = (x[23]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[33];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[14];
  assign t[48] = t[61] ^ x[20];
  assign t[49] = t[62] ^ x[26];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[27];
  assign t[51] = t[64] ^ x[28];
  assign t[52] = t[65] ^ x[29];
  assign t[53] = t[66] ^ x[30];
  assign t[54] = t[67] ^ x[31];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[33];
  assign t[57] = t[70] ^ x[34];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = (~t[72] & t[73]);
  assign t[5] = t[8];
  assign t[60] = (~t[74] & t[75]);
  assign t[61] = (~t[76] & t[77]);
  assign t[62] = (~t[78] & t[79]);
  assign t[63] = (~t[74] & t[80]);
  assign t[64] = (~t[74] & t[81]);
  assign t[65] = (~t[76] & t[82]);
  assign t[66] = (~t[76] & t[83]);
  assign t[67] = (~t[78] & t[84]);
  assign t[68] = (~t[78] & t[85]);
  assign t[69] = (~t[74] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[76] & t[87]);
  assign t[71] = (~t[78] & t[88]);
  assign t[72] = t[89] ^ x[7];
  assign t[73] = t[90] ^ x[8];
  assign t[74] = t[91] ^ x[13];
  assign t[75] = t[92] ^ x[14];
  assign t[76] = t[93] ^ x[19];
  assign t[77] = t[94] ^ x[20];
  assign t[78] = t[95] ^ x[25];
  assign t[79] = t[96] ^ x[26];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[27];
  assign t[81] = t[98] ^ x[28];
  assign t[82] = t[99] ^ x[29];
  assign t[83] = t[100] ^ x[30];
  assign t[84] = t[101] ^ x[31];
  assign t[85] = t[102] ^ x[32];
  assign t[86] = t[103] ^ x[33];
  assign t[87] = t[104] ^ x[34];
  assign t[88] = t[105] ^ x[35];
  assign t[89] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[6]);
  assign t[91] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[92] = (x[10]);
  assign t[93] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[94] = (x[16]);
  assign t[95] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[96] = (x[22]);
  assign t[97] = (x[12]);
  assign t[98] = (x[9]);
  assign t[99] = (x[18]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [35:0] x;
 output y;

 wire [106:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[18]);
  assign t[101] = (x[15]);
  assign t[102] = (x[24]);
  assign t[103] = (x[21]);
  assign t[104] = (x[11]);
  assign t[105] = (x[17]);
  assign t[106] = (x[23]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = ~(t[21] & t[35]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[36]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[39] & t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[20];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[26];
  assign t[51] = t[64] ^ x[27];
  assign t[52] = t[65] ^ x[28];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[30];
  assign t[55] = t[68] ^ x[31];
  assign t[56] = t[69] ^ x[32];
  assign t[57] = t[70] ^ x[33];
  assign t[58] = t[71] ^ x[34];
  assign t[59] = t[72] ^ x[35];
  assign t[5] = t[7];
  assign t[60] = (~t[73] & t[74]);
  assign t[61] = (~t[75] & t[76]);
  assign t[62] = (~t[77] & t[78]);
  assign t[63] = (~t[79] & t[80]);
  assign t[64] = (~t[75] & t[81]);
  assign t[65] = (~t[75] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (~t[75] & t[87]);
  assign t[71] = (~t[77] & t[88]);
  assign t[72] = (~t[79] & t[89]);
  assign t[73] = t[90] ^ x[4];
  assign t[74] = t[91] ^ x[5];
  assign t[75] = t[92] ^ x[13];
  assign t[76] = t[93] ^ x[14];
  assign t[77] = t[94] ^ x[19];
  assign t[78] = t[95] ^ x[20];
  assign t[79] = t[96] ^ x[25];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[97] ^ x[26];
  assign t[81] = t[98] ^ x[27];
  assign t[82] = t[99] ^ x[28];
  assign t[83] = t[100] ^ x[29];
  assign t[84] = t[101] ^ x[30];
  assign t[85] = t[102] ^ x[31];
  assign t[86] = t[103] ^ x[32];
  assign t[87] = t[104] ^ x[33];
  assign t[88] = t[105] ^ x[34];
  assign t[89] = t[106] ^ x[35];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[3]);
  assign t[92] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[93] = (x[10]);
  assign t[94] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[95] = (x[16]);
  assign t[96] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[97] = (x[22]);
  assign t[98] = (x[12]);
  assign t[99] = (x[9]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [32:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[14];
  assign t[42] = t[52] ^ x[15];
  assign t[43] = t[53] ^ x[21];
  assign t[44] = t[54] ^ x[22];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[29];
  assign t[47] = t[57] ^ x[30];
  assign t[48] = t[58] ^ x[31];
  assign t[49] = t[59] ^ x[32];
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[62] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = (~t[65] & t[67]);
  assign t[55] = (~t[68] & t[69]);
  assign t[56] = (~t[68] & t[70]);
  assign t[57] = (~t[62] & t[71]);
  assign t[58] = (~t[65] & t[72]);
  assign t[59] = (~t[68] & t[73]);
  assign t[5] = t[8];
  assign t[60] = t[74] ^ x[7];
  assign t[61] = t[75] ^ x[8];
  assign t[62] = t[76] ^ x[13];
  assign t[63] = t[77] ^ x[14];
  assign t[64] = t[78] ^ x[15];
  assign t[65] = t[79] ^ x[20];
  assign t[66] = t[80] ^ x[21];
  assign t[67] = t[81] ^ x[22];
  assign t[68] = t[82] ^ x[27];
  assign t[69] = t[83] ^ x[28];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[84] ^ x[29];
  assign t[71] = t[85] ^ x[30];
  assign t[72] = t[86] ^ x[31];
  assign t[73] = t[87] ^ x[32];
  assign t[74] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[6]);
  assign t[76] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[77] = (x[11]);
  assign t[78] = (x[9]);
  assign t[79] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[18]);
  assign t[81] = (x[16]);
  assign t[82] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[83] = (x[25]);
  assign t[84] = (x[23]);
  assign t[85] = (x[12]);
  assign t[86] = (x[19]);
  assign t[87] = (x[26]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [35:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[11]);
  assign t[101] = (x[12]);
  assign t[102] = (x[17]);
  assign t[103] = (x[18]);
  assign t[104] = (x[23]);
  assign t[105] = (x[24]);
  assign t[106] = (x[9]);
  assign t[107] = (x[15]);
  assign t[108] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[36];
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[14];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[28];
  assign t[55] = t[68] ^ x[29];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[31];
  assign t[58] = t[71] ^ x[32];
  assign t[59] = t[72] ^ x[33];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[34];
  assign t[61] = t[74] ^ x[35];
  assign t[62] = (~t[75] & t[76]);
  assign t[63] = (~t[77] & t[78]);
  assign t[64] = (~t[79] & t[80]);
  assign t[65] = (~t[81] & t[82]);
  assign t[66] = (~t[77] & t[83]);
  assign t[67] = (~t[77] & t[84]);
  assign t[68] = (~t[79] & t[85]);
  assign t[69] = (~t[79] & t[86]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (~t[81] & t[87]);
  assign t[71] = (~t[81] & t[88]);
  assign t[72] = (~t[77] & t[89]);
  assign t[73] = (~t[79] & t[90]);
  assign t[74] = (~t[81] & t[91]);
  assign t[75] = t[92] ^ x[7];
  assign t[76] = t[93] ^ x[8];
  assign t[77] = t[94] ^ x[13];
  assign t[78] = t[95] ^ x[14];
  assign t[79] = t[96] ^ x[19];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ x[20];
  assign t[81] = t[98] ^ x[25];
  assign t[82] = t[99] ^ x[26];
  assign t[83] = t[100] ^ x[27];
  assign t[84] = t[101] ^ x[28];
  assign t[85] = t[102] ^ x[29];
  assign t[86] = t[103] ^ x[30];
  assign t[87] = t[104] ^ x[31];
  assign t[88] = t[105] ^ x[32];
  assign t[89] = t[106] ^ x[33];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[107] ^ x[34];
  assign t[91] = t[108] ^ x[35];
  assign t[92] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[6]);
  assign t[94] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[95] = (x[10]);
  assign t[96] = (x[15] & ~x[16] & ~x[17] & ~x[18]) | (~x[15] & x[16] & ~x[17] & ~x[18]) | (~x[15] & ~x[16] & x[17] & ~x[18]) | (~x[15] & ~x[16] & ~x[17] & x[18]) | (x[15] & x[16] & x[17] & ~x[18]) | (x[15] & x[16] & ~x[17] & x[18]) | (x[15] & ~x[16] & x[17] & x[18]) | (~x[15] & x[16] & x[17] & x[18]);
  assign t[97] = (x[16]);
  assign t[98] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[99] = (x[22]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [369:0] x;
 output [134:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[18], x[17], x[16], x[6]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[18], x[17], x[16], x[6]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[15], x[14], x[13], x[6]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[15], x[14], x[13], x[6]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[12], x[11], x[10], x[18], x[17], x[16], x[6]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[12], x[11], x[10], x[18], x[17], x[16], x[6]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[24], x[23], x[22], x[6]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[24], x[23], x[22], x[6]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[27], x[26], x[25], x[6]}), .y(y[30]));
  R2ind31 R2ind31_inst(.y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.x({x[27], x[26], x[25], x[6]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[9], x[8], x[7], x[6]}), .y(y[35]));
  R2ind36 R2ind36_inst(.y(y[36]));
  R2ind37 R2ind37_inst(.y(y[37]));
  R2ind38 R2ind38_inst(.y(y[38]));
  R2ind39 R2ind39_inst(.x({x[9], x[8], x[7], x[6]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[6]}), .y(y[40]));
  R2ind41 R2ind41_inst(.y(y[41]));
  R2ind42 R2ind42_inst(.y(y[42]));
  R2ind43 R2ind43_inst(.y(y[43]));
  R2ind44 R2ind44_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[6]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[30], x[29], x[28], x[6]}), .y(y[45]));
  R2ind46 R2ind46_inst(.y(y[46]));
  R2ind47 R2ind47_inst(.y(y[47]));
  R2ind48 R2ind48_inst(.y(y[48]));
  R2ind49 R2ind49_inst(.x({x[30], x[29], x[28], x[6]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[30], x[29], x[28], x[33], x[32], x[31], x[6]}), .y(y[50]));
  R2ind51 R2ind51_inst(.y(y[51]));
  R2ind52 R2ind52_inst(.y(y[52]));
  R2ind53 R2ind53_inst(.y(y[53]));
  R2ind54 R2ind54_inst(.x({x[30], x[29], x[28], x[33], x[32], x[31], x[6]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[36], x[6], x[35], x[34]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[43], x[45], x[44], x[30], x[29], x[28], x[42], x[41], x[40], x[39], x[38], x[37], x[54], x[6], x[53], x[52]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[43], x[45], x[44], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[51], x[6], x[50], x[49]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[44], x[30], x[29], x[28], x[45], x[43], x[41], x[40], x[39], x[38], x[37], x[48], x[6], x[47], x[46]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[36], x[6], x[35], x[34]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[30], x[29], x[28], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[6], x[56], x[55]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[64], x[66], x[65], x[30], x[29], x[28], x[63], x[62], x[61], x[60], x[59], x[58], x[75], x[6], x[74], x[73]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[64], x[66], x[65], x[30], x[29], x[28], x[63], x[62], x[61], x[60], x[59], x[58], x[72], x[6], x[71], x[70]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[65], x[30], x[29], x[28], x[66], x[64], x[62], x[61], x[60], x[59], x[58], x[69], x[6], x[68], x[67]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[66], x[65], x[64], x[30], x[29], x[28], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[6], x[56], x[55]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[6], x[77], x[76]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[85], x[87], x[86], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[96], x[6], x[95], x[94]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[85], x[87], x[86], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[93], x[6], x[92], x[91]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[86], x[30], x[29], x[28], x[87], x[85], x[83], x[82], x[81], x[80], x[79], x[90], x[6], x[89], x[88]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[87], x[86], x[85], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[6], x[77], x[76]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[6], x[98], x[97]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[106], x[108], x[107], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[117], x[6], x[116], x[115]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[106], x[108], x[107], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[114], x[6], x[113], x[112]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[107], x[30], x[29], x[28], x[108], x[106], x[104], x[103], x[102], x[101], x[100], x[111], x[6], x[110], x[109]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[108], x[107], x[106], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[6], x[98], x[97]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[30], x[29], x[28], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[6], x[119], x[118]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[127], x[129], x[128], x[30], x[29], x[28], x[126], x[125], x[124], x[123], x[122], x[121], x[138], x[6], x[137], x[136]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[127], x[129], x[128], x[30], x[29], x[28], x[126], x[125], x[124], x[123], x[122], x[121], x[135], x[6], x[134], x[133]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[128], x[30], x[29], x[28], x[129], x[127], x[125], x[124], x[123], x[122], x[121], x[132], x[6], x[131], x[130]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[129], x[128], x[127], x[30], x[29], x[28], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[6], x[119], x[118]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[30], x[29], x[28], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[6], x[140], x[139]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[148], x[150], x[149], x[147], x[146], x[145], x[144], x[143], x[142], x[30], x[29], x[28], x[159], x[6], x[158], x[157]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[148], x[150], x[149], x[147], x[146], x[145], x[144], x[143], x[142], x[30], x[29], x[28], x[156], x[6], x[155], x[154]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[149], x[30], x[29], x[28], x[150], x[148], x[146], x[145], x[144], x[143], x[142], x[153], x[6], x[152], x[151]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[150], x[149], x[148], x[30], x[29], x[28], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[6], x[140], x[139]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[30], x[29], x[28], x[162], x[6], x[161], x[160]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[169], x[171], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[30], x[29], x[28], x[180], x[6], x[179], x[178]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[169], x[171], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[30], x[29], x[28], x[177], x[6], x[176], x[175]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[170], x[171], x[169], x[167], x[166], x[165], x[164], x[163], x[30], x[29], x[28], x[174], x[6], x[173], x[172]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[30], x[29], x[28], x[162], x[6], x[161], x[160]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[30], x[29], x[28], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[6], x[182], x[181]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[190], x[192], x[191], x[30], x[29], x[28], x[189], x[188], x[187], x[186], x[185], x[184], x[201], x[6], x[200], x[199]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[190], x[192], x[191], x[30], x[29], x[28], x[189], x[188], x[187], x[186], x[185], x[184], x[198], x[6], x[197], x[196]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[191], x[30], x[29], x[28], x[192], x[190], x[188], x[187], x[186], x[185], x[184], x[195], x[6], x[194], x[193]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[192], x[191], x[190], x[30], x[29], x[28], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[6], x[182], x[181]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[222], x[54], x[221], x[220], x[219], x[51], x[218], x[217], x[216], x[48], x[215], x[214], x[213], x[45], x[212], x[211], x[44], x[43], x[210], x[209], x[208], x[207], x[206], x[205], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[204], x[36], x[6], x[203], x[202]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[211], x[43], x[213], x[212], x[45], x[44], x[210], x[209], x[208], x[207], x[206], x[205], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[222], x[54], x[6], x[221], x[220]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[211], x[43], x[213], x[212], x[45], x[44], x[210], x[209], x[208], x[207], x[206], x[205], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[219], x[51], x[6], x[218], x[217]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[212], x[44], x[213], x[211], x[209], x[208], x[207], x[206], x[205], x[45], x[43], x[41], x[40], x[39], x[38], x[37], x[216], x[48], x[30], x[29], x[28], x[6], x[215], x[214]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[213], x[45], x[212], x[211], x[44], x[43], x[210], x[209], x[208], x[207], x[206], x[205], x[42], x[41], x[40], x[39], x[38], x[37], x[30], x[29], x[28], x[204], x[36], x[6], x[203], x[202]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[243], x[75], x[242], x[241], x[240], x[72], x[239], x[238], x[237], x[69], x[236], x[235], x[234], x[66], x[233], x[232], x[65], x[64], x[231], x[230], x[229], x[228], x[227], x[226], x[63], x[62], x[61], x[60], x[59], x[58], x[225], x[57], x[30], x[29], x[28], x[6], x[224], x[223]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[232], x[64], x[234], x[233], x[66], x[65], x[231], x[230], x[229], x[228], x[227], x[226], x[63], x[62], x[61], x[60], x[59], x[58], x[243], x[75], x[30], x[29], x[28], x[6], x[242], x[241]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[232], x[64], x[234], x[233], x[66], x[65], x[231], x[230], x[229], x[228], x[227], x[226], x[63], x[62], x[61], x[60], x[59], x[58], x[30], x[29], x[28], x[240], x[72], x[6], x[239], x[238]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[233], x[65], x[234], x[232], x[230], x[229], x[228], x[227], x[226], x[66], x[64], x[62], x[61], x[60], x[59], x[58], x[30], x[29], x[28], x[237], x[69], x[6], x[236], x[235]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[234], x[66], x[233], x[232], x[65], x[64], x[231], x[230], x[229], x[228], x[227], x[226], x[63], x[62], x[61], x[60], x[59], x[58], x[225], x[57], x[30], x[29], x[28], x[6], x[224], x[223]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[264], x[96], x[263], x[262], x[261], x[93], x[15], x[14], x[13], x[260], x[259], x[258], x[90], x[18], x[17], x[16], x[257], x[256], x[255], x[87], x[254], x[253], x[86], x[85], x[252], x[251], x[250], x[249], x[248], x[247], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[246], x[78], x[12], x[11], x[10], x[6], x[245], x[244]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[253], x[85], x[255], x[254], x[87], x[86], x[252], x[251], x[250], x[249], x[248], x[247], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[264], x[96], x[6], x[263], x[262]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[253], x[85], x[255], x[254], x[87], x[86], x[252], x[251], x[250], x[249], x[248], x[247], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[261], x[93], x[15], x[14], x[13], x[6], x[260], x[259]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[254], x[86], x[255], x[253], x[251], x[250], x[249], x[248], x[247], x[30], x[29], x[28], x[87], x[85], x[83], x[82], x[81], x[80], x[79], x[258], x[90], x[18], x[17], x[16], x[6], x[257], x[256]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[255], x[87], x[254], x[253], x[86], x[85], x[252], x[251], x[250], x[249], x[248], x[247], x[30], x[29], x[28], x[84], x[83], x[82], x[81], x[80], x[79], x[246], x[78], x[12], x[11], x[10], x[6], x[245], x[244]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[285], x[117], x[9], x[8], x[7], x[284], x[283], x[282], x[114], x[27], x[26], x[25], x[281], x[280], x[279], x[111], x[24], x[23], x[22], x[278], x[277], x[276], x[108], x[275], x[274], x[107], x[106], x[273], x[272], x[271], x[270], x[269], x[268], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[267], x[99], x[21], x[20], x[19], x[6], x[266], x[265]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[274], x[106], x[276], x[275], x[108], x[107], x[273], x[272], x[271], x[270], x[269], x[268], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[285], x[117], x[9], x[8], x[7], x[6], x[284], x[283]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[274], x[106], x[276], x[275], x[108], x[107], x[273], x[272], x[271], x[270], x[269], x[268], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[282], x[114], x[27], x[26], x[25], x[6], x[281], x[280]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[275], x[107], x[276], x[274], x[272], x[271], x[270], x[269], x[268], x[30], x[29], x[28], x[108], x[106], x[104], x[103], x[102], x[101], x[100], x[279], x[111], x[24], x[23], x[22], x[6], x[278], x[277]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[276], x[108], x[275], x[274], x[107], x[106], x[273], x[272], x[271], x[270], x[269], x[268], x[30], x[29], x[28], x[105], x[104], x[103], x[102], x[101], x[100], x[267], x[99], x[21], x[20], x[19], x[6], x[266], x[265]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[54], x[138], x[306], x[305], x[304], x[51], x[135], x[303], x[302], x[301], x[48], x[132], x[300], x[299], x[298], x[45], x[129], x[297], x[44], x[43], x[128], x[127], x[296], x[295], x[42], x[41], x[40], x[39], x[38], x[37], x[126], x[125], x[124], x[123], x[122], x[121], x[294], x[293], x[292], x[291], x[290], x[289], x[30], x[29], x[28], x[36], x[120], x[288], x[6], x[287], x[286]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[43], x[127], x[295], x[45], x[44], x[129], x[128], x[297], x[296], x[42], x[41], x[40], x[39], x[38], x[37], x[126], x[125], x[124], x[123], x[122], x[121], x[294], x[293], x[292], x[291], x[290], x[289], x[30], x[29], x[28], x[54], x[138], x[306], x[6], x[305], x[304]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[43], x[127], x[295], x[45], x[44], x[129], x[128], x[297], x[296], x[42], x[41], x[40], x[39], x[38], x[37], x[126], x[125], x[124], x[123], x[122], x[121], x[294], x[293], x[292], x[291], x[290], x[289], x[30], x[29], x[28], x[51], x[135], x[303], x[6], x[302], x[301]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[44], x[128], x[296], x[45], x[43], x[41], x[40], x[39], x[38], x[37], x[129], x[127], x[125], x[124], x[123], x[122], x[121], x[297], x[295], x[293], x[292], x[291], x[290], x[289], x[30], x[29], x[28], x[48], x[132], x[300], x[6], x[299], x[298]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[45], x[129], x[297], x[44], x[43], x[128], x[127], x[296], x[295], x[42], x[41], x[40], x[39], x[38], x[37], x[126], x[125], x[124], x[123], x[122], x[121], x[294], x[293], x[292], x[291], x[290], x[289], x[30], x[29], x[28], x[36], x[120], x[288], x[6], x[287], x[286]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[75], x[159], x[327], x[326], x[325], x[72], x[156], x[324], x[323], x[322], x[69], x[153], x[321], x[320], x[319], x[66], x[150], x[318], x[65], x[64], x[149], x[148], x[317], x[316], x[63], x[62], x[61], x[60], x[59], x[58], x[147], x[146], x[145], x[144], x[143], x[142], x[315], x[314], x[313], x[312], x[311], x[310], x[30], x[29], x[28], x[57], x[141], x[309], x[6], x[308], x[307]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[64], x[148], x[316], x[66], x[65], x[150], x[149], x[318], x[317], x[63], x[62], x[61], x[60], x[59], x[58], x[147], x[146], x[145], x[144], x[143], x[142], x[315], x[314], x[313], x[312], x[311], x[310], x[30], x[29], x[28], x[75], x[159], x[327], x[6], x[326], x[325]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[64], x[148], x[316], x[66], x[65], x[150], x[149], x[318], x[317], x[63], x[62], x[61], x[60], x[59], x[58], x[147], x[146], x[145], x[144], x[143], x[142], x[315], x[314], x[313], x[312], x[311], x[310], x[72], x[156], x[324], x[30], x[29], x[28], x[6], x[323], x[322]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[65], x[149], x[317], x[66], x[64], x[62], x[61], x[60], x[59], x[58], x[150], x[148], x[146], x[145], x[144], x[143], x[142], x[318], x[316], x[314], x[313], x[312], x[311], x[310], x[69], x[153], x[321], x[30], x[29], x[28], x[6], x[320], x[319]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[66], x[150], x[318], x[65], x[64], x[149], x[148], x[317], x[316], x[63], x[62], x[61], x[60], x[59], x[58], x[147], x[146], x[145], x[144], x[143], x[142], x[315], x[314], x[313], x[312], x[311], x[310], x[30], x[29], x[28], x[57], x[141], x[309], x[6], x[308], x[307]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[96], x[180], x[348], x[347], x[346], x[93], x[177], x[345], x[344], x[343], x[90], x[174], x[342], x[341], x[340], x[87], x[171], x[339], x[86], x[85], x[170], x[169], x[338], x[337], x[84], x[83], x[82], x[81], x[80], x[79], x[168], x[167], x[166], x[165], x[164], x[163], x[336], x[335], x[334], x[333], x[332], x[331], x[78], x[162], x[330], x[30], x[29], x[28], x[6], x[329], x[328]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[85], x[169], x[337], x[87], x[86], x[171], x[170], x[339], x[338], x[84], x[83], x[82], x[81], x[80], x[79], x[168], x[167], x[166], x[165], x[164], x[163], x[336], x[335], x[334], x[333], x[332], x[331], x[96], x[180], x[348], x[30], x[29], x[28], x[6], x[347], x[346]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[85], x[169], x[337], x[87], x[86], x[171], x[170], x[339], x[338], x[84], x[83], x[82], x[81], x[80], x[79], x[168], x[167], x[166], x[165], x[164], x[163], x[336], x[335], x[334], x[333], x[332], x[331], x[30], x[29], x[28], x[93], x[177], x[345], x[6], x[344], x[343]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[86], x[170], x[338], x[87], x[85], x[83], x[82], x[81], x[80], x[79], x[171], x[169], x[167], x[166], x[165], x[164], x[163], x[339], x[337], x[335], x[334], x[333], x[332], x[331], x[30], x[29], x[28], x[90], x[174], x[342], x[6], x[341], x[340]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[87], x[171], x[339], x[86], x[85], x[170], x[169], x[338], x[337], x[84], x[83], x[82], x[81], x[80], x[79], x[168], x[167], x[166], x[165], x[164], x[163], x[336], x[335], x[334], x[333], x[332], x[331], x[78], x[162], x[330], x[30], x[29], x[28], x[6], x[329], x[328]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[117], x[201], x[369], x[368], x[367], x[114], x[198], x[366], x[365], x[364], x[111], x[195], x[363], x[362], x[361], x[108], x[192], x[360], x[107], x[106], x[191], x[190], x[359], x[358], x[105], x[104], x[103], x[102], x[101], x[100], x[189], x[188], x[187], x[186], x[185], x[184], x[357], x[356], x[355], x[354], x[353], x[352], x[30], x[29], x[28], x[99], x[183], x[351], x[6], x[350], x[349]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[106], x[190], x[358], x[108], x[107], x[192], x[191], x[360], x[359], x[105], x[104], x[103], x[102], x[101], x[100], x[189], x[188], x[187], x[186], x[185], x[184], x[357], x[356], x[355], x[354], x[353], x[352], x[30], x[29], x[28], x[117], x[201], x[369], x[6], x[368], x[367]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[106], x[190], x[358], x[108], x[107], x[192], x[191], x[360], x[359], x[105], x[104], x[103], x[102], x[101], x[100], x[189], x[188], x[187], x[186], x[185], x[184], x[357], x[356], x[355], x[354], x[353], x[352], x[114], x[198], x[366], x[30], x[29], x[28], x[6], x[365], x[364]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[107], x[191], x[359], x[108], x[106], x[104], x[103], x[102], x[101], x[100], x[192], x[190], x[188], x[187], x[186], x[185], x[184], x[360], x[358], x[356], x[355], x[354], x[353], x[352], x[30], x[29], x[28], x[111], x[195], x[363], x[6], x[362], x[361]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[108], x[192], x[360], x[107], x[106], x[191], x[190], x[359], x[358], x[105], x[104], x[103], x[102], x[101], x[100], x[189], x[188], x[187], x[186], x[185], x[184], x[357], x[356], x[355], x[354], x[353], x[352], x[30], x[29], x[28], x[99], x[183], x[351], x[6], x[350], x[349]}), .y(y[134]));
endmodule

