/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [87:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_438 ;
    wire signal_441 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(1)) cell_176 ( .a ({X_s1[0], X_s0[0]}), .b ({signal_438, signal_192}) ) ;
    INV_X1 cell_177 ( .A ( 1'b1 ), .ZN ( signal_193 ) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_178 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[4], X_s0[4]}), .c ({signal_441, signal_194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[5], X_s0[5]}), .c ({signal_444, signal_195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .a ({X_s1[7], X_s0[7]}), .b ({X_s1[4], X_s0[4]}), .c ({signal_445, signal_196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .a ({X_s1[6], X_s0[6]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_446, signal_197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .a ({X_s1[3], X_s0[3]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_448, signal_198}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_183 ( .a ({signal_445, signal_196}), .b ({signal_449, signal_199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .a ({X_s1[6], X_s0[6]}), .b ({signal_445, signal_196}), .c ({signal_452, signal_202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_187 ( .a ({X_s1[2], X_s0[2]}), .b ({signal_444, signal_195}), .c ({signal_454, signal_203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_188 ( .a ({signal_444, signal_195}), .b ({signal_446, signal_197}), .c ({signal_455, signal_204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_189 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_446, signal_197}), .c ({signal_457, signal_205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_190 ( .a ({X_s1[4], X_s0[4]}), .b ({signal_448, signal_198}), .c ({signal_458, signal_206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_191 ( .a ({X_s1[5], X_s0[5]}), .b ({signal_446, signal_197}), .c ({signal_459, signal_207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_192 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_448, signal_198}), .c ({signal_460, signal_208}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_193 ( .a ({signal_455, signal_204}), .b ({signal_461, signal_209}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_194 ( .a ({signal_459, signal_207}), .b ({signal_462, signal_210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_201 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_459, signal_207}), .c ({signal_469, signal_217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_202 ( .a ({signal_454, signal_203}), .b ({signal_457, signal_205}), .c ({signal_470, signal_218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_203 ( .a ({X_s1[4], X_s0[4]}), .b ({signal_457, signal_205}), .c ({signal_471, signal_219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_204 ( .a ({X_s1[3], X_s0[3]}), .b ({signal_457, signal_205}), .c ({signal_472, signal_220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_205 ( .a ({X_s1[4], X_s0[4]}), .b ({signal_459, signal_207}), .c ({signal_473, signal_221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_206 ( .a ({signal_445, signal_196}), .b ({signal_460, signal_208}), .c ({signal_474, signal_222}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_208 ( .a ({signal_469, signal_217}), .b ({signal_476, signal_224}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_209 ( .a ({signal_470, signal_218}), .b ({signal_477, signal_225}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_210 ( .a ({signal_473, signal_221}), .b ({signal_478, signal_226}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_211 ( .a ({signal_474, signal_222}), .b ({signal_479, signal_227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_219 ( .a ({X_s1[2], X_s0[2]}), .b ({signal_472, signal_220}), .c ({signal_487, signal_235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_220 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_473, signal_221}), .c ({signal_488, signal_236}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_222 ( .a ({signal_487, signal_235}), .b ({signal_490, signal_238}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_223 ( .a ({signal_488, signal_236}), .b ({signal_491, signal_239}) ) ;

    /* cells in depth 1 */
    buf_clk cell_669 ( .C ( clk ), .D ( signal_193 ), .Q ( signal_1033 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .a ({signal_438, signal_192}), .b ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_450, signal_200}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .a ({1'b0, signal_193}), .b ({signal_441, signal_194}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_451, signal_201}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_195 ( .a ({signal_450, signal_200}), .b ({signal_463, signal_211}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_196 ( .a ({signal_451, signal_201}), .b ({signal_464, signal_212}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_197 ( .a ({1'b0, signal_193}), .b ({signal_454, signal_203}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_465, signal_213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_198 ( .a ({1'b0, signal_193}), .b ({signal_458, signal_206}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_466, signal_214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_199 ( .a ({1'b0, signal_193}), .b ({signal_449, signal_199}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_467, signal_215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_200 ( .a ({1'b0, signal_193}), .b ({signal_452, signal_202}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_468, signal_216}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_207 ( .a ({signal_465, signal_213}), .b ({signal_475, signal_223}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_212 ( .a ({signal_466, signal_214}), .b ({signal_480, signal_228}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_213 ( .a ({signal_467, signal_215}), .b ({signal_481, signal_229}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_214 ( .a ({signal_468, signal_216}), .b ({signal_482, signal_230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_215 ( .a ({1'b0, 1'b1}), .b ({signal_462, signal_210}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_483, signal_231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_216 ( .a ({1'b0, signal_193}), .b ({signal_471, signal_219}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_484, signal_232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_217 ( .a ({1'b0, signal_193}), .b ({signal_472, signal_220}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_485, signal_233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_218 ( .a ({1'b0, 1'b1}), .b ({signal_461, signal_209}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_486, signal_234}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_221 ( .a ({signal_483, signal_231}), .b ({signal_489, signal_237}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_224 ( .a ({signal_484, signal_232}), .b ({signal_492, signal_240}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_225 ( .a ({signal_485, signal_233}), .b ({signal_493, signal_241}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_226 ( .a ({signal_486, signal_234}), .b ({signal_494, signal_242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_228 ( .a ({1'b0, 1'b1}), .b ({signal_477, signal_225}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_496, signal_244}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_229 ( .a ({1'b0, 1'b1}), .b ({signal_478, signal_226}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_497, signal_245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_230 ( .a ({1'b0, 1'b1}), .b ({signal_476, signal_224}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_498, signal_246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_231 ( .a ({1'b0, 1'b1}), .b ({signal_479, signal_227}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_499, signal_247}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_232 ( .a ({signal_496, signal_244}), .b ({signal_500, signal_248}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_233 ( .a ({signal_497, signal_245}), .b ({signal_501, signal_249}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_234 ( .a ({signal_498, signal_246}), .b ({signal_502, signal_250}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_235 ( .a ({signal_499, signal_247}), .b ({signal_503, signal_251}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({1'b0, signal_193}), .b ({signal_491, signal_239}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_506, signal_254}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .a ({1'b0, 1'b1}), .b ({signal_490, signal_238}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_507, signal_255}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_241 ( .a ({signal_506, signal_254}), .b ({signal_509, signal_257}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_242 ( .a ({signal_507, signal_255}), .b ({signal_510, signal_258}) ) ;
    buf_clk cell_670 ( .C ( clk ), .D ( signal_1033 ), .Q ( signal_1034 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_671 ( .C ( clk ), .D ( signal_1034 ), .Q ( signal_1035 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_227 ( .a ({signal_475, signal_223}), .b ({signal_463, signal_211}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_495, signal_243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({signal_480, signal_228}), .b ({signal_489, signal_237}), .clk ( clk ), .r ( Fresh[17] ), .c ({signal_504, signal_252}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({signal_493, signal_241}), .b ({signal_494, signal_242}), .clk ( clk ), .r ( Fresh[18] ), .c ({signal_505, signal_253}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_240 ( .a ({signal_505, signal_253}), .b ({signal_508, signal_256}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({signal_481, signal_229}), .b ({signal_500, signal_248}), .clk ( clk ), .r ( Fresh[19] ), .c ({signal_511, signal_259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .a ({signal_492, signal_240}), .b ({signal_501, signal_249}), .clk ( clk ), .r ( Fresh[20] ), .c ({signal_512, signal_260}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .a ({signal_464, signal_212}), .b ({signal_502, signal_250}), .clk ( clk ), .r ( Fresh[21] ), .c ({signal_513, signal_261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .a ({signal_482, signal_230}), .b ({signal_503, signal_251}), .clk ( clk ), .r ( Fresh[22] ), .c ({signal_514, signal_262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .a ({signal_509, signal_257}), .b ({signal_510, signal_258}), .clk ( clk ), .r ( Fresh[23] ), .c ({signal_515, signal_263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .a ({signal_495, signal_243}), .b ({signal_514, signal_262}), .c ({signal_519, signal_267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .a ({signal_504, signal_252}), .b ({signal_514, signal_262}), .c ({signal_520, signal_268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .a ({signal_513, signal_261}), .b ({signal_505, signal_253}), .c ({signal_521, signal_269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .a ({signal_511, signal_259}), .b ({signal_512, signal_260}), .c ({signal_522, signal_270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .a ({signal_512, signal_260}), .b ({signal_505, signal_253}), .c ({signal_523, signal_271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .a ({signal_511, signal_259}), .b ({signal_513, signal_261}), .c ({signal_524, signal_272}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_257 ( .a ({signal_515, signal_263}), .b ({signal_525, signal_273}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_258 ( .a ({signal_520, signal_268}), .b ({signal_526, signal_274}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_259 ( .a ({signal_521, signal_269}), .b ({signal_527, signal_275}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_260 ( .a ({signal_523, signal_271}), .b ({signal_528, signal_276}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_261 ( .a ({signal_524, signal_272}), .b ({signal_529, signal_277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .a ({signal_504, signal_252}), .b ({signal_515, signal_263}), .c ({signal_532, signal_280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .a ({signal_495, signal_243}), .b ({signal_515, signal_263}), .c ({signal_533, signal_281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .a ({signal_523, signal_271}), .b ({signal_524, signal_272}), .c ({signal_534, signal_282}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_267 ( .a ({signal_532, signal_280}), .b ({signal_535, signal_283}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_268 ( .a ({signal_533, signal_281}), .b ({signal_536, signal_284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .a ({signal_520, signal_268}), .b ({signal_533, signal_281}), .c ({signal_541, signal_289}) ) ;
    buf_clk cell_672 ( .C ( clk ), .D ( signal_1035 ), .Q ( signal_1036 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_453 ( .C ( clk ), .D ( signal_262 ), .Q ( signal_817 ) ) ;
    buf_clk cell_459 ( .C ( clk ), .D ( signal_514 ), .Q ( signal_823 ) ) ;
    buf_clk cell_465 ( .C ( clk ), .D ( signal_243 ), .Q ( signal_829 ) ) ;
    buf_clk cell_471 ( .C ( clk ), .D ( signal_495 ), .Q ( signal_835 ) ) ;
    buf_clk cell_477 ( .C ( clk ), .D ( signal_252 ), .Q ( signal_841 ) ) ;
    buf_clk cell_483 ( .C ( clk ), .D ( signal_504 ), .Q ( signal_847 ) ) ;
    buf_clk cell_489 ( .C ( clk ), .D ( signal_263 ), .Q ( signal_853 ) ) ;
    buf_clk cell_495 ( .C ( clk ), .D ( signal_515 ), .Q ( signal_859 ) ) ;
    buf_clk cell_501 ( .C ( clk ), .D ( signal_259 ), .Q ( signal_865 ) ) ;
    buf_clk cell_507 ( .C ( clk ), .D ( signal_511 ), .Q ( signal_871 ) ) ;
    buf_clk cell_513 ( .C ( clk ), .D ( signal_260 ), .Q ( signal_877 ) ) ;
    buf_clk cell_519 ( .C ( clk ), .D ( signal_512 ), .Q ( signal_883 ) ) ;
    buf_clk cell_525 ( .C ( clk ), .D ( signal_261 ), .Q ( signal_889 ) ) ;
    buf_clk cell_531 ( .C ( clk ), .D ( signal_513 ), .Q ( signal_895 ) ) ;
    buf_clk cell_537 ( .C ( clk ), .D ( signal_253 ), .Q ( signal_901 ) ) ;
    buf_clk cell_543 ( .C ( clk ), .D ( signal_505 ), .Q ( signal_907 ) ) ;
    buf_clk cell_549 ( .C ( clk ), .D ( signal_267 ), .Q ( signal_913 ) ) ;
    buf_clk cell_555 ( .C ( clk ), .D ( signal_519 ), .Q ( signal_919 ) ) ;
    buf_clk cell_561 ( .C ( clk ), .D ( signal_280 ), .Q ( signal_925 ) ) ;
    buf_clk cell_567 ( .C ( clk ), .D ( signal_532 ), .Q ( signal_931 ) ) ;
    buf_clk cell_573 ( .C ( clk ), .D ( signal_268 ), .Q ( signal_937 ) ) ;
    buf_clk cell_579 ( .C ( clk ), .D ( signal_520 ), .Q ( signal_943 ) ) ;
    buf_clk cell_585 ( .C ( clk ), .D ( signal_281 ), .Q ( signal_949 ) ) ;
    buf_clk cell_591 ( .C ( clk ), .D ( signal_533 ), .Q ( signal_955 ) ) ;
    buf_clk cell_597 ( .C ( clk ), .D ( signal_270 ), .Q ( signal_961 ) ) ;
    buf_clk cell_603 ( .C ( clk ), .D ( signal_522 ), .Q ( signal_967 ) ) ;
    buf_clk cell_609 ( .C ( clk ), .D ( signal_269 ), .Q ( signal_973 ) ) ;
    buf_clk cell_615 ( .C ( clk ), .D ( signal_521 ), .Q ( signal_979 ) ) ;
    buf_clk cell_621 ( .C ( clk ), .D ( signal_272 ), .Q ( signal_985 ) ) ;
    buf_clk cell_627 ( .C ( clk ), .D ( signal_524 ), .Q ( signal_991 ) ) ;
    buf_clk cell_633 ( .C ( clk ), .D ( signal_271 ), .Q ( signal_997 ) ) ;
    buf_clk cell_639 ( .C ( clk ), .D ( signal_523 ), .Q ( signal_1003 ) ) ;
    buf_clk cell_645 ( .C ( clk ), .D ( signal_289 ), .Q ( signal_1009 ) ) ;
    buf_clk cell_651 ( .C ( clk ), .D ( signal_541 ), .Q ( signal_1015 ) ) ;
    buf_clk cell_657 ( .C ( clk ), .D ( signal_282 ), .Q ( signal_1021 ) ) ;
    buf_clk cell_663 ( .C ( clk ), .D ( signal_534 ), .Q ( signal_1027 ) ) ;
    buf_clk cell_673 ( .C ( clk ), .D ( signal_1036 ), .Q ( signal_1037 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .a ({signal_511, signal_259}), .b ({signal_514, signal_262}), .clk ( clk ), .r ( Fresh[24] ), .c ({signal_516, signal_264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .a ({signal_495, signal_243}), .b ({signal_512, signal_260}), .clk ( clk ), .r ( Fresh[25] ), .c ({signal_517, signal_265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .a ({signal_504, signal_252}), .b ({signal_513, signal_261}), .clk ( clk ), .r ( Fresh[26] ), .c ({signal_518, signal_266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .a ({signal_519, signal_267}), .b ({signal_522, signal_270}), .clk ( clk ), .r ( Fresh[27] ), .c ({signal_530, signal_278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .a ({signal_520, signal_268}), .b ({signal_524, signal_272}), .clk ( clk ), .r ( Fresh[28] ), .c ({signal_531, signal_279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .a ({signal_526, signal_274}), .b ({signal_529, signal_277}), .clk ( clk ), .r ( Fresh[29] ), .c ({signal_537, signal_285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .a ({signal_508, signal_256}), .b ({signal_525, signal_273}), .clk ( clk ), .r ( Fresh[30] ), .c ({signal_538, signal_286}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .a ({signal_521, signal_269}), .b ({signal_532, signal_280}), .clk ( clk ), .r ( Fresh[31] ), .c ({signal_539, signal_287}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .a ({signal_523, signal_271}), .b ({signal_533, signal_281}), .clk ( clk ), .r ( Fresh[32] ), .c ({signal_540, signal_288}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .a ({signal_528, signal_276}), .b ({signal_536, signal_284}), .clk ( clk ), .r ( Fresh[33] ), .c ({signal_542, signal_290}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .a ({signal_527, signal_275}), .b ({signal_535, signal_283}), .clk ( clk ), .r ( Fresh[34] ), .c ({signal_543, signal_291}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .a ({signal_534, signal_282}), .b ({signal_541, signal_289}), .clk ( clk ), .r ( Fresh[35] ), .c ({signal_544, signal_292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .a ({signal_517, signal_265}), .b ({signal_537, signal_285}), .c ({signal_545, signal_293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .a ({signal_530, signal_278}), .b ({signal_540, signal_288}), .c ({signal_546, signal_294}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .a ({signal_538, signal_286}), .b ({signal_539, signal_287}), .c ({signal_547, signal_295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_280 ( .a ({signal_516, signal_264}), .b ({signal_542, signal_290}), .c ({signal_548, signal_296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_281 ( .a ({signal_518, signal_266}), .b ({signal_543, signal_291}), .c ({signal_549, signal_297}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_282 ( .a ({signal_530, signal_278}), .b ({signal_544, signal_292}), .c ({signal_550, signal_298}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_283 ( .a ({signal_545, signal_293}), .b ({signal_546, signal_294}), .c ({signal_551, signal_299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_284 ( .a ({signal_540, signal_288}), .b ({signal_544, signal_292}), .c ({signal_552, signal_300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_285 ( .a ({signal_531, signal_279}), .b ({signal_547, signal_295}), .c ({signal_553, signal_301}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_286 ( .a ({signal_551, signal_299}), .b ({signal_554, signal_302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_287 ( .a ({signal_548, signal_296}), .b ({signal_550, signal_298}), .c ({signal_555, signal_303}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_288 ( .a ({signal_549, signal_297}), .b ({signal_552, signal_300}), .c ({signal_556, signal_304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_289 ( .a ({signal_540, signal_288}), .b ({signal_553, signal_301}), .c ({signal_557, signal_305}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_290 ( .a ({signal_555, signal_303}), .b ({signal_558, signal_306}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_291 ( .a ({signal_556, signal_304}), .b ({signal_559, signal_307}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_292 ( .a ({signal_557, signal_305}), .b ({signal_560, signal_308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_294 ( .a ({signal_551, signal_299}), .b ({signal_555, signal_303}), .c ({signal_562, signal_310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_295 ( .a ({signal_556, signal_304}), .b ({signal_557, signal_305}), .c ({signal_563, signal_311}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_296 ( .a ({signal_562, signal_310}), .b ({signal_564, signal_312}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_297 ( .a ({signal_563, signal_311}), .b ({signal_565, signal_313}) ) ;
    buf_clk cell_454 ( .C ( clk ), .D ( signal_817 ), .Q ( signal_818 ) ) ;
    buf_clk cell_460 ( .C ( clk ), .D ( signal_823 ), .Q ( signal_824 ) ) ;
    buf_clk cell_466 ( .C ( clk ), .D ( signal_829 ), .Q ( signal_830 ) ) ;
    buf_clk cell_472 ( .C ( clk ), .D ( signal_835 ), .Q ( signal_836 ) ) ;
    buf_clk cell_478 ( .C ( clk ), .D ( signal_841 ), .Q ( signal_842 ) ) ;
    buf_clk cell_484 ( .C ( clk ), .D ( signal_847 ), .Q ( signal_848 ) ) ;
    buf_clk cell_490 ( .C ( clk ), .D ( signal_853 ), .Q ( signal_854 ) ) ;
    buf_clk cell_496 ( .C ( clk ), .D ( signal_859 ), .Q ( signal_860 ) ) ;
    buf_clk cell_502 ( .C ( clk ), .D ( signal_865 ), .Q ( signal_866 ) ) ;
    buf_clk cell_508 ( .C ( clk ), .D ( signal_871 ), .Q ( signal_872 ) ) ;
    buf_clk cell_514 ( .C ( clk ), .D ( signal_877 ), .Q ( signal_878 ) ) ;
    buf_clk cell_520 ( .C ( clk ), .D ( signal_883 ), .Q ( signal_884 ) ) ;
    buf_clk cell_526 ( .C ( clk ), .D ( signal_889 ), .Q ( signal_890 ) ) ;
    buf_clk cell_532 ( .C ( clk ), .D ( signal_895 ), .Q ( signal_896 ) ) ;
    buf_clk cell_538 ( .C ( clk ), .D ( signal_901 ), .Q ( signal_902 ) ) ;
    buf_clk cell_544 ( .C ( clk ), .D ( signal_907 ), .Q ( signal_908 ) ) ;
    buf_clk cell_550 ( .C ( clk ), .D ( signal_913 ), .Q ( signal_914 ) ) ;
    buf_clk cell_556 ( .C ( clk ), .D ( signal_919 ), .Q ( signal_920 ) ) ;
    buf_clk cell_562 ( .C ( clk ), .D ( signal_925 ), .Q ( signal_926 ) ) ;
    buf_clk cell_568 ( .C ( clk ), .D ( signal_931 ), .Q ( signal_932 ) ) ;
    buf_clk cell_574 ( .C ( clk ), .D ( signal_937 ), .Q ( signal_938 ) ) ;
    buf_clk cell_580 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_944 ) ) ;
    buf_clk cell_586 ( .C ( clk ), .D ( signal_949 ), .Q ( signal_950 ) ) ;
    buf_clk cell_592 ( .C ( clk ), .D ( signal_955 ), .Q ( signal_956 ) ) ;
    buf_clk cell_598 ( .C ( clk ), .D ( signal_961 ), .Q ( signal_962 ) ) ;
    buf_clk cell_604 ( .C ( clk ), .D ( signal_967 ), .Q ( signal_968 ) ) ;
    buf_clk cell_610 ( .C ( clk ), .D ( signal_973 ), .Q ( signal_974 ) ) ;
    buf_clk cell_616 ( .C ( clk ), .D ( signal_979 ), .Q ( signal_980 ) ) ;
    buf_clk cell_622 ( .C ( clk ), .D ( signal_985 ), .Q ( signal_986 ) ) ;
    buf_clk cell_628 ( .C ( clk ), .D ( signal_991 ), .Q ( signal_992 ) ) ;
    buf_clk cell_634 ( .C ( clk ), .D ( signal_997 ), .Q ( signal_998 ) ) ;
    buf_clk cell_640 ( .C ( clk ), .D ( signal_1003 ), .Q ( signal_1004 ) ) ;
    buf_clk cell_646 ( .C ( clk ), .D ( signal_1009 ), .Q ( signal_1010 ) ) ;
    buf_clk cell_652 ( .C ( clk ), .D ( signal_1015 ), .Q ( signal_1016 ) ) ;
    buf_clk cell_658 ( .C ( clk ), .D ( signal_1021 ), .Q ( signal_1022 ) ) ;
    buf_clk cell_664 ( .C ( clk ), .D ( signal_1027 ), .Q ( signal_1028 ) ) ;
    buf_clk cell_674 ( .C ( clk ), .D ( signal_1037 ), .Q ( signal_1038 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_429 ( .C ( clk ), .D ( signal_308 ), .Q ( signal_793 ) ) ;
    buf_clk cell_431 ( .C ( clk ), .D ( signal_560 ), .Q ( signal_795 ) ) ;
    buf_clk cell_433 ( .C ( clk ), .D ( signal_302 ), .Q ( signal_797 ) ) ;
    buf_clk cell_435 ( .C ( clk ), .D ( signal_554 ), .Q ( signal_799 ) ) ;
    buf_clk cell_437 ( .C ( clk ), .D ( signal_307 ), .Q ( signal_801 ) ) ;
    buf_clk cell_439 ( .C ( clk ), .D ( signal_559 ), .Q ( signal_803 ) ) ;
    buf_clk cell_441 ( .C ( clk ), .D ( signal_306 ), .Q ( signal_805 ) ) ;
    buf_clk cell_443 ( .C ( clk ), .D ( signal_558 ), .Q ( signal_807 ) ) ;
    buf_clk cell_445 ( .C ( clk ), .D ( signal_311 ), .Q ( signal_809 ) ) ;
    buf_clk cell_447 ( .C ( clk ), .D ( signal_563 ), .Q ( signal_811 ) ) ;
    buf_clk cell_449 ( .C ( clk ), .D ( signal_310 ), .Q ( signal_813 ) ) ;
    buf_clk cell_451 ( .C ( clk ), .D ( signal_562 ), .Q ( signal_815 ) ) ;
    buf_clk cell_455 ( .C ( clk ), .D ( signal_818 ), .Q ( signal_819 ) ) ;
    buf_clk cell_461 ( .C ( clk ), .D ( signal_824 ), .Q ( signal_825 ) ) ;
    buf_clk cell_467 ( .C ( clk ), .D ( signal_830 ), .Q ( signal_831 ) ) ;
    buf_clk cell_473 ( .C ( clk ), .D ( signal_836 ), .Q ( signal_837 ) ) ;
    buf_clk cell_479 ( .C ( clk ), .D ( signal_842 ), .Q ( signal_843 ) ) ;
    buf_clk cell_485 ( .C ( clk ), .D ( signal_848 ), .Q ( signal_849 ) ) ;
    buf_clk cell_491 ( .C ( clk ), .D ( signal_854 ), .Q ( signal_855 ) ) ;
    buf_clk cell_497 ( .C ( clk ), .D ( signal_860 ), .Q ( signal_861 ) ) ;
    buf_clk cell_503 ( .C ( clk ), .D ( signal_866 ), .Q ( signal_867 ) ) ;
    buf_clk cell_509 ( .C ( clk ), .D ( signal_872 ), .Q ( signal_873 ) ) ;
    buf_clk cell_515 ( .C ( clk ), .D ( signal_878 ), .Q ( signal_879 ) ) ;
    buf_clk cell_521 ( .C ( clk ), .D ( signal_884 ), .Q ( signal_885 ) ) ;
    buf_clk cell_527 ( .C ( clk ), .D ( signal_890 ), .Q ( signal_891 ) ) ;
    buf_clk cell_533 ( .C ( clk ), .D ( signal_896 ), .Q ( signal_897 ) ) ;
    buf_clk cell_539 ( .C ( clk ), .D ( signal_902 ), .Q ( signal_903 ) ) ;
    buf_clk cell_545 ( .C ( clk ), .D ( signal_908 ), .Q ( signal_909 ) ) ;
    buf_clk cell_551 ( .C ( clk ), .D ( signal_914 ), .Q ( signal_915 ) ) ;
    buf_clk cell_557 ( .C ( clk ), .D ( signal_920 ), .Q ( signal_921 ) ) ;
    buf_clk cell_563 ( .C ( clk ), .D ( signal_926 ), .Q ( signal_927 ) ) ;
    buf_clk cell_569 ( .C ( clk ), .D ( signal_932 ), .Q ( signal_933 ) ) ;
    buf_clk cell_575 ( .C ( clk ), .D ( signal_938 ), .Q ( signal_939 ) ) ;
    buf_clk cell_581 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_945 ) ) ;
    buf_clk cell_587 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_951 ) ) ;
    buf_clk cell_593 ( .C ( clk ), .D ( signal_956 ), .Q ( signal_957 ) ) ;
    buf_clk cell_599 ( .C ( clk ), .D ( signal_962 ), .Q ( signal_963 ) ) ;
    buf_clk cell_605 ( .C ( clk ), .D ( signal_968 ), .Q ( signal_969 ) ) ;
    buf_clk cell_611 ( .C ( clk ), .D ( signal_974 ), .Q ( signal_975 ) ) ;
    buf_clk cell_617 ( .C ( clk ), .D ( signal_980 ), .Q ( signal_981 ) ) ;
    buf_clk cell_623 ( .C ( clk ), .D ( signal_986 ), .Q ( signal_987 ) ) ;
    buf_clk cell_629 ( .C ( clk ), .D ( signal_992 ), .Q ( signal_993 ) ) ;
    buf_clk cell_635 ( .C ( clk ), .D ( signal_998 ), .Q ( signal_999 ) ) ;
    buf_clk cell_641 ( .C ( clk ), .D ( signal_1004 ), .Q ( signal_1005 ) ) ;
    buf_clk cell_647 ( .C ( clk ), .D ( signal_1010 ), .Q ( signal_1011 ) ) ;
    buf_clk cell_653 ( .C ( clk ), .D ( signal_1016 ), .Q ( signal_1017 ) ) ;
    buf_clk cell_659 ( .C ( clk ), .D ( signal_1022 ), .Q ( signal_1023 ) ) ;
    buf_clk cell_665 ( .C ( clk ), .D ( signal_1028 ), .Q ( signal_1029 ) ) ;
    buf_clk cell_675 ( .C ( clk ), .D ( signal_1038 ), .Q ( signal_1039 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_293 ( .a ({signal_555, signal_303}), .b ({signal_556, signal_304}), .clk ( clk ), .r ( Fresh[36] ), .c ({signal_561, signal_309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_298 ( .a ({signal_554, signal_302}), .b ({signal_560, signal_308}), .clk ( clk ), .r ( Fresh[37] ), .c ({signal_566, signal_314}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_299 ( .a ({signal_562, signal_310}), .b ({signal_563, signal_311}), .clk ( clk ), .r ( Fresh[38] ), .c ({signal_567, signal_315}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_300 ( .a ({signal_564, signal_312}), .b ({signal_565, signal_313}), .clk ( clk ), .r ( Fresh[39] ), .c ({signal_568, signal_316}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_301 ( .a ({signal_561, signal_309}), .b ({signal_567, signal_315}), .c ({signal_569, signal_317}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_302 ( .a ({signal_569, signal_317}), .b ({signal_570, signal_318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_303 ( .a ({signal_566, signal_314}), .b ({signal_568, signal_316}), .c ({signal_571, signal_319}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_304 ( .a ({signal_571, signal_319}), .b ({signal_572, signal_320}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_307 ( .a ({signal_569, signal_317}), .b ({signal_571, signal_319}), .c ({signal_575, signal_323}) ) ;
    buf_clk cell_430 ( .C ( clk ), .D ( signal_793 ), .Q ( signal_794 ) ) ;
    buf_clk cell_432 ( .C ( clk ), .D ( signal_795 ), .Q ( signal_796 ) ) ;
    buf_clk cell_434 ( .C ( clk ), .D ( signal_797 ), .Q ( signal_798 ) ) ;
    buf_clk cell_436 ( .C ( clk ), .D ( signal_799 ), .Q ( signal_800 ) ) ;
    buf_clk cell_438 ( .C ( clk ), .D ( signal_801 ), .Q ( signal_802 ) ) ;
    buf_clk cell_440 ( .C ( clk ), .D ( signal_803 ), .Q ( signal_804 ) ) ;
    buf_clk cell_442 ( .C ( clk ), .D ( signal_805 ), .Q ( signal_806 ) ) ;
    buf_clk cell_444 ( .C ( clk ), .D ( signal_807 ), .Q ( signal_808 ) ) ;
    buf_clk cell_446 ( .C ( clk ), .D ( signal_809 ), .Q ( signal_810 ) ) ;
    buf_clk cell_448 ( .C ( clk ), .D ( signal_811 ), .Q ( signal_812 ) ) ;
    buf_clk cell_450 ( .C ( clk ), .D ( signal_813 ), .Q ( signal_814 ) ) ;
    buf_clk cell_452 ( .C ( clk ), .D ( signal_815 ), .Q ( signal_816 ) ) ;
    buf_clk cell_456 ( .C ( clk ), .D ( signal_819 ), .Q ( signal_820 ) ) ;
    buf_clk cell_462 ( .C ( clk ), .D ( signal_825 ), .Q ( signal_826 ) ) ;
    buf_clk cell_468 ( .C ( clk ), .D ( signal_831 ), .Q ( signal_832 ) ) ;
    buf_clk cell_474 ( .C ( clk ), .D ( signal_837 ), .Q ( signal_838 ) ) ;
    buf_clk cell_480 ( .C ( clk ), .D ( signal_843 ), .Q ( signal_844 ) ) ;
    buf_clk cell_486 ( .C ( clk ), .D ( signal_849 ), .Q ( signal_850 ) ) ;
    buf_clk cell_492 ( .C ( clk ), .D ( signal_855 ), .Q ( signal_856 ) ) ;
    buf_clk cell_498 ( .C ( clk ), .D ( signal_861 ), .Q ( signal_862 ) ) ;
    buf_clk cell_504 ( .C ( clk ), .D ( signal_867 ), .Q ( signal_868 ) ) ;
    buf_clk cell_510 ( .C ( clk ), .D ( signal_873 ), .Q ( signal_874 ) ) ;
    buf_clk cell_516 ( .C ( clk ), .D ( signal_879 ), .Q ( signal_880 ) ) ;
    buf_clk cell_522 ( .C ( clk ), .D ( signal_885 ), .Q ( signal_886 ) ) ;
    buf_clk cell_528 ( .C ( clk ), .D ( signal_891 ), .Q ( signal_892 ) ) ;
    buf_clk cell_534 ( .C ( clk ), .D ( signal_897 ), .Q ( signal_898 ) ) ;
    buf_clk cell_540 ( .C ( clk ), .D ( signal_903 ), .Q ( signal_904 ) ) ;
    buf_clk cell_546 ( .C ( clk ), .D ( signal_909 ), .Q ( signal_910 ) ) ;
    buf_clk cell_552 ( .C ( clk ), .D ( signal_915 ), .Q ( signal_916 ) ) ;
    buf_clk cell_558 ( .C ( clk ), .D ( signal_921 ), .Q ( signal_922 ) ) ;
    buf_clk cell_564 ( .C ( clk ), .D ( signal_927 ), .Q ( signal_928 ) ) ;
    buf_clk cell_570 ( .C ( clk ), .D ( signal_933 ), .Q ( signal_934 ) ) ;
    buf_clk cell_576 ( .C ( clk ), .D ( signal_939 ), .Q ( signal_940 ) ) ;
    buf_clk cell_582 ( .C ( clk ), .D ( signal_945 ), .Q ( signal_946 ) ) ;
    buf_clk cell_588 ( .C ( clk ), .D ( signal_951 ), .Q ( signal_952 ) ) ;
    buf_clk cell_594 ( .C ( clk ), .D ( signal_957 ), .Q ( signal_958 ) ) ;
    buf_clk cell_600 ( .C ( clk ), .D ( signal_963 ), .Q ( signal_964 ) ) ;
    buf_clk cell_606 ( .C ( clk ), .D ( signal_969 ), .Q ( signal_970 ) ) ;
    buf_clk cell_612 ( .C ( clk ), .D ( signal_975 ), .Q ( signal_976 ) ) ;
    buf_clk cell_618 ( .C ( clk ), .D ( signal_981 ), .Q ( signal_982 ) ) ;
    buf_clk cell_624 ( .C ( clk ), .D ( signal_987 ), .Q ( signal_988 ) ) ;
    buf_clk cell_630 ( .C ( clk ), .D ( signal_993 ), .Q ( signal_994 ) ) ;
    buf_clk cell_636 ( .C ( clk ), .D ( signal_999 ), .Q ( signal_1000 ) ) ;
    buf_clk cell_642 ( .C ( clk ), .D ( signal_1005 ), .Q ( signal_1006 ) ) ;
    buf_clk cell_648 ( .C ( clk ), .D ( signal_1011 ), .Q ( signal_1012 ) ) ;
    buf_clk cell_654 ( .C ( clk ), .D ( signal_1017 ), .Q ( signal_1018 ) ) ;
    buf_clk cell_660 ( .C ( clk ), .D ( signal_1023 ), .Q ( signal_1024 ) ) ;
    buf_clk cell_666 ( .C ( clk ), .D ( signal_1029 ), .Q ( signal_1030 ) ) ;
    buf_clk cell_676 ( .C ( clk ), .D ( signal_1039 ), .Q ( signal_1040 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_457 ( .C ( clk ), .D ( signal_820 ), .Q ( signal_821 ) ) ;
    buf_clk cell_463 ( .C ( clk ), .D ( signal_826 ), .Q ( signal_827 ) ) ;
    buf_clk cell_469 ( .C ( clk ), .D ( signal_832 ), .Q ( signal_833 ) ) ;
    buf_clk cell_475 ( .C ( clk ), .D ( signal_838 ), .Q ( signal_839 ) ) ;
    buf_clk cell_481 ( .C ( clk ), .D ( signal_844 ), .Q ( signal_845 ) ) ;
    buf_clk cell_487 ( .C ( clk ), .D ( signal_850 ), .Q ( signal_851 ) ) ;
    buf_clk cell_493 ( .C ( clk ), .D ( signal_856 ), .Q ( signal_857 ) ) ;
    buf_clk cell_499 ( .C ( clk ), .D ( signal_862 ), .Q ( signal_863 ) ) ;
    buf_clk cell_505 ( .C ( clk ), .D ( signal_868 ), .Q ( signal_869 ) ) ;
    buf_clk cell_511 ( .C ( clk ), .D ( signal_874 ), .Q ( signal_875 ) ) ;
    buf_clk cell_517 ( .C ( clk ), .D ( signal_880 ), .Q ( signal_881 ) ) ;
    buf_clk cell_523 ( .C ( clk ), .D ( signal_886 ), .Q ( signal_887 ) ) ;
    buf_clk cell_529 ( .C ( clk ), .D ( signal_892 ), .Q ( signal_893 ) ) ;
    buf_clk cell_535 ( .C ( clk ), .D ( signal_898 ), .Q ( signal_899 ) ) ;
    buf_clk cell_541 ( .C ( clk ), .D ( signal_904 ), .Q ( signal_905 ) ) ;
    buf_clk cell_547 ( .C ( clk ), .D ( signal_910 ), .Q ( signal_911 ) ) ;
    buf_clk cell_553 ( .C ( clk ), .D ( signal_916 ), .Q ( signal_917 ) ) ;
    buf_clk cell_559 ( .C ( clk ), .D ( signal_922 ), .Q ( signal_923 ) ) ;
    buf_clk cell_565 ( .C ( clk ), .D ( signal_928 ), .Q ( signal_929 ) ) ;
    buf_clk cell_571 ( .C ( clk ), .D ( signal_934 ), .Q ( signal_935 ) ) ;
    buf_clk cell_577 ( .C ( clk ), .D ( signal_940 ), .Q ( signal_941 ) ) ;
    buf_clk cell_583 ( .C ( clk ), .D ( signal_946 ), .Q ( signal_947 ) ) ;
    buf_clk cell_589 ( .C ( clk ), .D ( signal_952 ), .Q ( signal_953 ) ) ;
    buf_clk cell_595 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_959 ) ) ;
    buf_clk cell_601 ( .C ( clk ), .D ( signal_964 ), .Q ( signal_965 ) ) ;
    buf_clk cell_607 ( .C ( clk ), .D ( signal_970 ), .Q ( signal_971 ) ) ;
    buf_clk cell_613 ( .C ( clk ), .D ( signal_976 ), .Q ( signal_977 ) ) ;
    buf_clk cell_619 ( .C ( clk ), .D ( signal_982 ), .Q ( signal_983 ) ) ;
    buf_clk cell_625 ( .C ( clk ), .D ( signal_988 ), .Q ( signal_989 ) ) ;
    buf_clk cell_631 ( .C ( clk ), .D ( signal_994 ), .Q ( signal_995 ) ) ;
    buf_clk cell_637 ( .C ( clk ), .D ( signal_1000 ), .Q ( signal_1001 ) ) ;
    buf_clk cell_643 ( .C ( clk ), .D ( signal_1006 ), .Q ( signal_1007 ) ) ;
    buf_clk cell_649 ( .C ( clk ), .D ( signal_1012 ), .Q ( signal_1013 ) ) ;
    buf_clk cell_655 ( .C ( clk ), .D ( signal_1018 ), .Q ( signal_1019 ) ) ;
    buf_clk cell_661 ( .C ( clk ), .D ( signal_1024 ), .Q ( signal_1025 ) ) ;
    buf_clk cell_667 ( .C ( clk ), .D ( signal_1030 ), .Q ( signal_1031 ) ) ;
    buf_clk cell_677 ( .C ( clk ), .D ( signal_1040 ), .Q ( signal_1041 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_305 ( .a ({signal_796, signal_794}), .b ({signal_570, signal_318}), .clk ( clk ), .r ( Fresh[40] ), .c ({signal_573, signal_321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_306 ( .a ({signal_800, signal_798}), .b ({signal_570, signal_318}), .clk ( clk ), .r ( Fresh[41] ), .c ({signal_574, signal_322}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_308 ( .a ({signal_804, signal_802}), .b ({signal_572, signal_320}), .clk ( clk ), .r ( Fresh[42] ), .c ({signal_576, signal_324}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_309 ( .a ({signal_808, signal_806}), .b ({signal_572, signal_320}), .clk ( clk ), .r ( Fresh[43] ), .c ({signal_577, signal_325}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_310 ( .a ({signal_812, signal_810}), .b ({signal_575, signal_323}), .clk ( clk ), .r ( Fresh[44] ), .c ({signal_578, signal_326}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_311 ( .a ({signal_816, signal_814}), .b ({signal_575, signal_323}), .clk ( clk ), .r ( Fresh[45] ), .c ({signal_579, signal_327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_312 ( .a ({signal_576, signal_324}), .b ({signal_578, signal_326}), .c ({signal_580, signal_328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_313 ( .a ({signal_573, signal_321}), .b ({signal_578, signal_326}), .c ({signal_581, signal_329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_314 ( .a ({signal_577, signal_325}), .b ({signal_579, signal_327}), .c ({signal_582, signal_330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_315 ( .a ({signal_574, signal_322}), .b ({signal_579, signal_327}), .c ({signal_583, signal_331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_324 ( .a ({signal_582, signal_330}), .b ({signal_583, signal_331}), .c ({signal_592, signal_340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_325 ( .a ({signal_580, signal_328}), .b ({signal_581, signal_329}), .c ({signal_593, signal_341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_326 ( .a ({signal_581, signal_329}), .b ({signal_583, signal_331}), .c ({signal_594, signal_342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_327 ( .a ({signal_580, signal_328}), .b ({signal_582, signal_330}), .c ({signal_595, signal_343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_336 ( .a ({signal_594, signal_342}), .b ({signal_595, signal_343}), .c ({signal_604, signal_352}) ) ;
    buf_clk cell_458 ( .C ( clk ), .D ( signal_821 ), .Q ( signal_822 ) ) ;
    buf_clk cell_464 ( .C ( clk ), .D ( signal_827 ), .Q ( signal_828 ) ) ;
    buf_clk cell_470 ( .C ( clk ), .D ( signal_833 ), .Q ( signal_834 ) ) ;
    buf_clk cell_476 ( .C ( clk ), .D ( signal_839 ), .Q ( signal_840 ) ) ;
    buf_clk cell_482 ( .C ( clk ), .D ( signal_845 ), .Q ( signal_846 ) ) ;
    buf_clk cell_488 ( .C ( clk ), .D ( signal_851 ), .Q ( signal_852 ) ) ;
    buf_clk cell_494 ( .C ( clk ), .D ( signal_857 ), .Q ( signal_858 ) ) ;
    buf_clk cell_500 ( .C ( clk ), .D ( signal_863 ), .Q ( signal_864 ) ) ;
    buf_clk cell_506 ( .C ( clk ), .D ( signal_869 ), .Q ( signal_870 ) ) ;
    buf_clk cell_512 ( .C ( clk ), .D ( signal_875 ), .Q ( signal_876 ) ) ;
    buf_clk cell_518 ( .C ( clk ), .D ( signal_881 ), .Q ( signal_882 ) ) ;
    buf_clk cell_524 ( .C ( clk ), .D ( signal_887 ), .Q ( signal_888 ) ) ;
    buf_clk cell_530 ( .C ( clk ), .D ( signal_893 ), .Q ( signal_894 ) ) ;
    buf_clk cell_536 ( .C ( clk ), .D ( signal_899 ), .Q ( signal_900 ) ) ;
    buf_clk cell_542 ( .C ( clk ), .D ( signal_905 ), .Q ( signal_906 ) ) ;
    buf_clk cell_548 ( .C ( clk ), .D ( signal_911 ), .Q ( signal_912 ) ) ;
    buf_clk cell_554 ( .C ( clk ), .D ( signal_917 ), .Q ( signal_918 ) ) ;
    buf_clk cell_560 ( .C ( clk ), .D ( signal_923 ), .Q ( signal_924 ) ) ;
    buf_clk cell_566 ( .C ( clk ), .D ( signal_929 ), .Q ( signal_930 ) ) ;
    buf_clk cell_572 ( .C ( clk ), .D ( signal_935 ), .Q ( signal_936 ) ) ;
    buf_clk cell_578 ( .C ( clk ), .D ( signal_941 ), .Q ( signal_942 ) ) ;
    buf_clk cell_584 ( .C ( clk ), .D ( signal_947 ), .Q ( signal_948 ) ) ;
    buf_clk cell_590 ( .C ( clk ), .D ( signal_953 ), .Q ( signal_954 ) ) ;
    buf_clk cell_596 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_960 ) ) ;
    buf_clk cell_602 ( .C ( clk ), .D ( signal_965 ), .Q ( signal_966 ) ) ;
    buf_clk cell_608 ( .C ( clk ), .D ( signal_971 ), .Q ( signal_972 ) ) ;
    buf_clk cell_614 ( .C ( clk ), .D ( signal_977 ), .Q ( signal_978 ) ) ;
    buf_clk cell_620 ( .C ( clk ), .D ( signal_983 ), .Q ( signal_984 ) ) ;
    buf_clk cell_626 ( .C ( clk ), .D ( signal_989 ), .Q ( signal_990 ) ) ;
    buf_clk cell_632 ( .C ( clk ), .D ( signal_995 ), .Q ( signal_996 ) ) ;
    buf_clk cell_638 ( .C ( clk ), .D ( signal_1001 ), .Q ( signal_1002 ) ) ;
    buf_clk cell_644 ( .C ( clk ), .D ( signal_1007 ), .Q ( signal_1008 ) ) ;
    buf_clk cell_650 ( .C ( clk ), .D ( signal_1013 ), .Q ( signal_1014 ) ) ;
    buf_clk cell_656 ( .C ( clk ), .D ( signal_1019 ), .Q ( signal_1020 ) ) ;
    buf_clk cell_662 ( .C ( clk ), .D ( signal_1025 ), .Q ( signal_1026 ) ) ;
    buf_clk cell_668 ( .C ( clk ), .D ( signal_1031 ), .Q ( signal_1032 ) ) ;
    buf_clk cell_678 ( .C ( clk ), .D ( signal_1041 ), .Q ( signal_1042 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_679 ( .C ( clk ), .D ( signal_1042 ), .Q ( signal_1043 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_316 ( .a ({signal_828, signal_822}), .b ({signal_580, signal_328}), .clk ( clk ), .r ( Fresh[46] ), .c ({signal_584, signal_332}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_317 ( .a ({signal_840, signal_834}), .b ({signal_581, signal_329}), .clk ( clk ), .r ( Fresh[47] ), .c ({signal_585, signal_333}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_318 ( .a ({signal_852, signal_846}), .b ({signal_582, signal_330}), .clk ( clk ), .r ( Fresh[48] ), .c ({signal_586, signal_334}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_319 ( .a ({signal_864, signal_858}), .b ({signal_583, signal_331}), .clk ( clk ), .r ( Fresh[49] ), .c ({signal_587, signal_335}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_320 ( .a ({signal_876, signal_870}), .b ({signal_580, signal_328}), .clk ( clk ), .r ( Fresh[50] ), .c ({signal_588, signal_336}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_321 ( .a ({signal_888, signal_882}), .b ({signal_581, signal_329}), .clk ( clk ), .r ( Fresh[51] ), .c ({signal_589, signal_337}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_322 ( .a ({signal_900, signal_894}), .b ({signal_582, signal_330}), .clk ( clk ), .r ( Fresh[52] ), .c ({signal_590, signal_338}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_323 ( .a ({signal_912, signal_906}), .b ({signal_583, signal_331}), .clk ( clk ), .r ( Fresh[53] ), .c ({signal_591, signal_339}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_328 ( .a ({signal_924, signal_918}), .b ({signal_593, signal_341}), .clk ( clk ), .r ( Fresh[54] ), .c ({signal_596, signal_344}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_329 ( .a ({signal_936, signal_930}), .b ({signal_592, signal_340}), .clk ( clk ), .r ( Fresh[55] ), .c ({signal_597, signal_345}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_330 ( .a ({signal_948, signal_942}), .b ({signal_595, signal_343}), .clk ( clk ), .r ( Fresh[56] ), .c ({signal_598, signal_346}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_331 ( .a ({signal_960, signal_954}), .b ({signal_594, signal_342}), .clk ( clk ), .r ( Fresh[57] ), .c ({signal_599, signal_347}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_332 ( .a ({signal_972, signal_966}), .b ({signal_593, signal_341}), .clk ( clk ), .r ( Fresh[58] ), .c ({signal_600, signal_348}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_333 ( .a ({signal_984, signal_978}), .b ({signal_592, signal_340}), .clk ( clk ), .r ( Fresh[59] ), .c ({signal_601, signal_349}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_334 ( .a ({signal_996, signal_990}), .b ({signal_595, signal_343}), .clk ( clk ), .r ( Fresh[60] ), .c ({signal_602, signal_350}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_335 ( .a ({signal_1008, signal_1002}), .b ({signal_594, signal_342}), .clk ( clk ), .r ( Fresh[61] ), .c ({signal_603, signal_351}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_337 ( .a ({signal_1020, signal_1014}), .b ({signal_604, signal_352}), .clk ( clk ), .r ( Fresh[62] ), .c ({signal_605, signal_353}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_338 ( .a ({signal_1032, signal_1026}), .b ({signal_604, signal_352}), .clk ( clk ), .r ( Fresh[63] ), .c ({signal_606, signal_354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_339 ( .a ({signal_584, signal_332}), .b ({signal_596, signal_344}), .c ({signal_607, signal_355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_340 ( .a ({signal_585, signal_333}), .b ({signal_596, signal_344}), .c ({signal_608, signal_356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_341 ( .a ({signal_586, signal_334}), .b ({signal_597, signal_345}), .c ({signal_609, signal_357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_342 ( .a ({signal_587, signal_335}), .b ({signal_597, signal_345}), .c ({signal_610, signal_358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_343 ( .a ({signal_598, signal_346}), .b ({signal_599, signal_347}), .c ({signal_611, signal_359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_344 ( .a ({signal_588, signal_336}), .b ({signal_600, signal_348}), .c ({signal_612, signal_360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_345 ( .a ({signal_589, signal_337}), .b ({signal_600, signal_348}), .c ({signal_613, signal_361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_346 ( .a ({signal_590, signal_338}), .b ({signal_601, signal_349}), .c ({signal_614, signal_362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_347 ( .a ({signal_591, signal_339}), .b ({signal_601, signal_349}), .c ({signal_615, signal_363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_348 ( .a ({signal_602, signal_350}), .b ({signal_603, signal_351}), .c ({signal_616, signal_364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_349 ( .a ({signal_608, signal_356}), .b ({signal_611, signal_359}), .c ({signal_617, signal_365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_350 ( .a ({signal_610, signal_358}), .b ({signal_611, signal_359}), .c ({signal_618, signal_366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_351 ( .a ({signal_599, signal_347}), .b ({signal_605, signal_353}), .c ({signal_619, signal_367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_352 ( .a ({signal_613, signal_361}), .b ({signal_616, signal_364}), .c ({signal_620, signal_368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_353 ( .a ({signal_615, signal_363}), .b ({signal_616, signal_364}), .c ({signal_621, signal_369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_354 ( .a ({signal_603, signal_351}), .b ({signal_606, signal_354}), .c ({signal_622, signal_370}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_355 ( .a ({signal_620, signal_368}), .b ({signal_623, signal_371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_356 ( .a ({signal_617, signal_365}), .b ({signal_621, signal_369}), .c ({signal_624, signal_372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_357 ( .a ({signal_617, signal_365}), .b ({signal_618, signal_366}), .c ({signal_625, signal_373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_358 ( .a ({signal_607, signal_355}), .b ({signal_619, signal_367}), .c ({signal_626, signal_374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_359 ( .a ({signal_609, signal_357}), .b ({signal_619, signal_367}), .c ({signal_627, signal_375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_360 ( .a ({signal_612, signal_360}), .b ({signal_622, signal_370}), .c ({signal_628, signal_376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_361 ( .a ({signal_614, signal_362}), .b ({signal_622, signal_370}), .c ({signal_629, signal_377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_364 ( .a ({signal_627, signal_375}), .b ({signal_629, signal_377}), .c ({signal_632, signal_380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_365 ( .a ({signal_618, signal_366}), .b ({signal_629, signal_377}), .c ({signal_633, signal_381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_366 ( .a ({signal_617, signal_365}), .b ({signal_629, signal_377}), .c ({signal_634, signal_382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_367 ( .a ({signal_626, signal_374}), .b ({signal_628, signal_376}), .c ({signal_635, signal_383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_368 ( .a ({signal_627, signal_375}), .b ({signal_628, signal_376}), .c ({signal_636, signal_384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_369 ( .a ({signal_625, signal_373}), .b ({signal_629, signal_377}), .c ({signal_637, signal_385}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_370 ( .a ({signal_632, signal_380}), .b ({signal_638, signal_386}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_371 ( .a ({signal_633, signal_381}), .b ({signal_639, signal_387}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_372 ( .a ({signal_634, signal_382}), .b ({signal_640, signal_388}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_373 ( .a ({signal_636, signal_384}), .b ({signal_641, signal_389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_378 ( .a ({signal_618, signal_366}), .b ({signal_632, signal_380}), .c ({signal_646, signal_394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_379 ( .a ({signal_627, signal_375}), .b ({signal_635, signal_383}), .c ({signal_647, signal_395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_380 ( .a ({signal_620, signal_368}), .b ({signal_636, signal_384}), .c ({signal_648, signal_396}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_381 ( .a ({signal_647, signal_395}), .b ({signal_649, signal_397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_389 ( .a ({signal_626, signal_374}), .b ({signal_646, signal_394}), .c ({signal_657, signal_405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_390 ( .a ({signal_624, signal_372}), .b ({signal_647, signal_395}), .c ({signal_658, signal_406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_391 ( .a ({signal_637, signal_385}), .b ({signal_648, signal_396}), .c ({signal_659, signal_407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_392 ( .a ({signal_625, signal_373}), .b ({signal_647, signal_395}), .c ({signal_660, signal_408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_393 ( .a ({signal_624, signal_372}), .b ({signal_648, signal_396}), .c ({signal_661, signal_409}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_396 ( .a ({signal_657, signal_405}), .b ({signal_664, signal_412}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_397 ( .a ({signal_659, signal_407}), .b ({signal_665, signal_413}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_398 ( .a ({signal_660, signal_408}), .b ({signal_666, signal_414}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_399 ( .a ({signal_661, signal_409}), .b ({signal_667, signal_415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_405 ( .a ({signal_629, signal_377}), .b ({signal_658, signal_406}), .c ({signal_673, signal_420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_406 ( .a ({signal_620, signal_368}), .b ({signal_658, signal_406}), .c ({signal_674, signal_421}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_408 ( .a ({signal_673, signal_420}), .b ({signal_676, signal_423}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_409 ( .a ({signal_674, signal_421}), .b ({signal_677, signal_424}) ) ;
    buf_clk cell_680 ( .C ( clk ), .D ( signal_1043 ), .Q ( signal_1044 ) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_362 ( .a ({1'b0, signal_1044}), .b ({signal_623, signal_371}), .clk ( clk ), .r ( Fresh[64] ), .c ({signal_630, signal_378}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_363 ( .a ({1'b0, 1'b1}), .b ({signal_624, signal_372}), .clk ( clk ), .r ( Fresh[65] ), .c ({signal_631, signal_379}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_374 ( .a ({signal_630, signal_378}), .b ({signal_642, signal_390}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_375 ( .a ({signal_631, signal_379}), .b ({signal_643, signal_391}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_637, signal_385}), .clk ( clk ), .r ( Fresh[66] ), .c ({signal_644, signal_392}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_377 ( .a ({1'b0, 1'b1}), .b ({signal_635, signal_383}), .clk ( clk ), .r ( Fresh[67] ), .c ({signal_645, signal_393}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_382 ( .a ({signal_644, signal_392}), .b ({signal_650, signal_398}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_383 ( .a ({signal_645, signal_393}), .b ({signal_651, signal_399}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_384 ( .a ({1'b0, signal_1044}), .b ({signal_639, signal_387}), .clk ( clk ), .r ( Fresh[68] ), .c ({signal_652, signal_400}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_385 ( .a ({1'b0, 1'b1}), .b ({signal_641, signal_389}), .clk ( clk ), .r ( Fresh[69] ), .c ({signal_653, signal_401}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_386 ( .a ({1'b0, signal_1044}), .b ({signal_640, signal_388}), .clk ( clk ), .r ( Fresh[70] ), .c ({signal_654, signal_402}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_387 ( .a ({1'b0, signal_1044}), .b ({signal_638, signal_386}), .clk ( clk ), .r ( Fresh[71] ), .c ({signal_655, signal_403}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_388 ( .a ({1'b0, 1'b1}), .b ({signal_646, signal_394}), .clk ( clk ), .r ( Fresh[72] ), .c ({signal_656, signal_404}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_394 ( .a ({signal_652, signal_400}), .b ({signal_662, signal_410}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_395 ( .a ({signal_653, signal_401}), .b ({signal_663, signal_411}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_400 ( .a ({signal_654, signal_402}), .b ({signal_668, signal_416}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_401 ( .a ({signal_655, signal_403}), .b ({signal_669, signal_417}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_402 ( .a ({signal_656, signal_404}), .b ({signal_670, signal_418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_404 ( .a ({1'b0, 1'b1}), .b ({signal_649, signal_397}), .clk ( clk ), .r ( Fresh[73] ), .c ({signal_672, signal_419}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_407 ( .a ({signal_672, signal_419}), .b ({signal_675, signal_422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_412 ( .a ({1'b0, signal_1044}), .b ({signal_665, signal_413}), .clk ( clk ), .r ( Fresh[74] ), .c ({signal_680, signal_425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_413 ( .a ({1'b0, 1'b1}), .b ({signal_666, signal_414}), .clk ( clk ), .r ( Fresh[75] ), .c ({signal_681, signal_426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_414 ( .a ({1'b0, signal_1044}), .b ({signal_664, signal_412}), .clk ( clk ), .r ( Fresh[76] ), .c ({signal_682, signal_427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_415 ( .a ({1'b0, 1'b1}), .b ({signal_667, signal_415}), .clk ( clk ), .r ( Fresh[77] ), .c ({signal_683, signal_428}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_416 ( .a ({signal_680, signal_425}), .b ({signal_684, signal_429}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_417 ( .a ({signal_681, signal_426}), .b ({signal_685, signal_430}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_418 ( .a ({signal_682, signal_427}), .b ({signal_686, signal_431}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_419 ( .a ({signal_683, signal_428}), .b ({signal_687, signal_432}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_421 ( .a ({1'b0, signal_1044}), .b ({signal_676, signal_423}), .clk ( clk ), .r ( Fresh[78] ), .c ({signal_689, signal_433}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_422 ( .a ({1'b0, signal_1044}), .b ({signal_677, signal_424}), .clk ( clk ), .r ( Fresh[79] ), .c ({signal_690, signal_434}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_423 ( .a ({signal_689, signal_433}), .b ({signal_691, signal_435}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_424 ( .a ({signal_690, signal_434}), .b ({signal_692, signal_436}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_403 ( .a ({signal_642, signal_390}), .b ({signal_650, signal_398}), .clk ( clk ), .r ( Fresh[80] ), .c ({signal_671, signal_167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_410 ( .a ({signal_662, signal_410}), .b ({signal_663, signal_411}), .clk ( clk ), .r ( Fresh[81] ), .c ({signal_678, signal_160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_411 ( .a ({signal_669, signal_417}), .b ({signal_670, signal_418}), .clk ( clk ), .r ( Fresh[82] ), .c ({signal_679, signal_166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_420 ( .a ({signal_668, signal_416}), .b ({signal_675, signal_422}), .clk ( clk ), .r ( Fresh[83] ), .c ({signal_688, signal_163}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_425 ( .a ({signal_684, signal_429}), .b ({signal_685, signal_430}), .clk ( clk ), .r ( Fresh[84] ), .c ({signal_693, signal_164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_426 ( .a ({signal_686, signal_431}), .b ({signal_687, signal_432}), .clk ( clk ), .r ( Fresh[85] ), .c ({signal_694, signal_165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_427 ( .a ({signal_691, signal_435}), .b ({signal_651, signal_399}), .clk ( clk ), .r ( Fresh[86] ), .c ({signal_695, signal_161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_428 ( .a ({signal_692, signal_436}), .b ({signal_643, signal_391}), .clk ( clk ), .r ( Fresh[87] ), .c ({signal_696, signal_162}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_678, signal_160}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_695, signal_161}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_696, signal_162}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_688, signal_163}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_693, signal_164}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_694, signal_165}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_679, signal_166}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_671, signal_167}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
