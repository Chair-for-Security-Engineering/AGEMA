/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* 17 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 18 register stage(s) in total */

module sbox_GHPCLL_Pipeline_d1 (SI_s0, clk, SI_s1, Fresh, SO_s0, SO_s1);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [3471:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;

    /* cells in depth 0 */
    not_masked #(.low_latency(1), .pipeline(1)) U1938 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_943, n2796}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1939 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_945, n2810}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1940 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_947, n2462}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1941 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_949, n2760}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1942 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_951, n2791}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1944 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_953, n2813}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1945 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_955, n2630}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1946 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_957, n2765}) ) ;

    /* cells in depth 1 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1937 ( .a ({new_AGEMA_signal_943, n2796}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_970, n2719}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1943 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1023, n2672}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1947 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[7], Fresh[6], Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_958, n2635}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1948 ( .a ({new_AGEMA_signal_947, n2462}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_971, n2641}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1949 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_959, n2790}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1950 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_960, n2519}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1951 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_972, n2750}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1952 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_973, n2615}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1953 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1024, n2640}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1955 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ({Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_974, n2699}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1956 ( .a ({new_AGEMA_signal_974, n2699}), .b ({new_AGEMA_signal_1025, n2737}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1957 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_975, n2816}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1958 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1026, n2767}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1961 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_976, n2780}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1962 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1027, n2789}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1963 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_977, n2317}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1965 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ({Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_978, n2694}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1966 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1028, n2769}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1969 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_979, n2073}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1970 ( .a ({new_AGEMA_signal_979, n2073}), .b ({new_AGEMA_signal_1029, n2707}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1971 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_961, n2315}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1972 ( .a ({SI_s1[0], SI_s0[0]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[55], Fresh[54], Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_962, n2682}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1973 ( .a ({new_AGEMA_signal_962, n2682}), .b ({new_AGEMA_signal_980, n2713}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1975 ( .a ({new_AGEMA_signal_953, n2813}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_981, n2723}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1976 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1031, n2688}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1978 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_982, n2725}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1979 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1032, n2541}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1984 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_983, n2815}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1985 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1033, n2086}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1987 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68]}), .c ({new_AGEMA_signal_984, n2600}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1990 ( .a ({new_AGEMA_signal_947, n2462}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_985, n2538}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1991 ( .a ({new_AGEMA_signal_985, n2538}), .b ({new_AGEMA_signal_1035, n2786}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1995 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76]}), .c ({new_AGEMA_signal_963, n2595}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1996 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_986, n2742}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1999 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_987, n2753}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2000 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1037, n2577}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2004 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_988, n2400}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2008 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[91], Fresh[90], Fresh[89], Fresh[88]}), .c ({new_AGEMA_signal_989, n2785}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2009 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1039, n2792}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2013 ( .a ({new_AGEMA_signal_953, n2813}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92]}), .c ({new_AGEMA_signal_990, n2609}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2014 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_1040, n2724}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2017 ( .a ({new_AGEMA_signal_949, n2760}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_991, n2661}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2018 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1041, n2174}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2020 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_964, n2708}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2021 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_992, n2493}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2025 ( .a ({new_AGEMA_signal_943, n2796}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104]}), .c ({new_AGEMA_signal_993, n2587}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2028 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1044, n2570}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2029 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_965, n2559}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2035 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .c ({new_AGEMA_signal_994, n2643}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2036 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1045, n2442}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2038 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_995, n2739}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2044 ( .a ({new_AGEMA_signal_947, n2462}), .b ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116]}), .c ({new_AGEMA_signal_996, n2437}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2045 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_966, n2261}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2046 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_997, n2778}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2052 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124]}), .c ({new_AGEMA_signal_998, n2452}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2055 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1050, n2766}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2068 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .c ({new_AGEMA_signal_1000, n2772}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2070 ( .a ({new_AGEMA_signal_951, n2791}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1001, n2824}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2071 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1053, n2612}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2074 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_1054, n2313}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2089 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136]}), .c ({new_AGEMA_signal_1002, n2395}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2090 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1058, n2818}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2094 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_967, n2779}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2096 ( .a ({new_AGEMA_signal_955, n2630}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ({Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1003, n2624}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2097 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[151], Fresh[150], Fresh[149], Fresh[148]}), .c ({new_AGEMA_signal_968, n2242}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2100 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152]}), .c ({new_AGEMA_signal_1004, n2356}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2119 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_1063, n2823}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2122 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1005, n2611}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2131 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1065, n2828}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2133 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({new_AGEMA_signal_1006, n2616}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2134 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1066, n2679}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2138 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164]}), .c ({new_AGEMA_signal_1007, n2563}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2139 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1067, n2809}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2150 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_1068, n2709}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2163 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .r ({Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1008, n2401}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2211 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[175], Fresh[174], Fresh[173], Fresh[172]}), .c ({new_AGEMA_signal_1010, n2061}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2232 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176]}), .c ({new_AGEMA_signal_1011, n2721}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2276 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .r ({Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1012, n2298}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2278 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_1080, n2118}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2307 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ({Fresh[187], Fresh[186], Fresh[185], Fresh[184]}), .c ({new_AGEMA_signal_1013, n2346}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2341 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188]}), .c ({new_AGEMA_signal_1015, n2430}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2383 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_969, n2712}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2402 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ({Fresh[199], Fresh[198], Fresh[197], Fresh[196]}), .c ({new_AGEMA_signal_1017, n2777}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2615 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_947, n2462}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .c ({new_AGEMA_signal_1019, n2463}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2627 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1020, n2474}) ) ;
    buf_clk new_AGEMA_reg_buffer_927 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( new_AGEMA_signal_5349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( new_AGEMA_signal_5350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( new_AGEMA_signal_5351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( new_AGEMA_signal_5352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( new_AGEMA_signal_5353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( new_AGEMA_signal_5354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( new_AGEMA_signal_5355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( new_AGEMA_signal_5356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_5357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_5358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C ( clk ), .D ( n2630 ), .Q ( new_AGEMA_signal_5359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C ( clk ), .D ( new_AGEMA_signal_955 ), .Q ( new_AGEMA_signal_5360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( new_AGEMA_signal_5361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( new_AGEMA_signal_5362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C ( clk ), .D ( n2462 ), .Q ( new_AGEMA_signal_5363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C ( clk ), .D ( new_AGEMA_signal_947 ), .Q ( new_AGEMA_signal_5364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C ( clk ), .D ( n2760 ), .Q ( new_AGEMA_signal_5365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C ( clk ), .D ( new_AGEMA_signal_949 ), .Q ( new_AGEMA_signal_5366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C ( clk ), .D ( n2796 ), .Q ( new_AGEMA_signal_5367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C ( clk ), .D ( new_AGEMA_signal_943 ), .Q ( new_AGEMA_signal_5368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C ( clk ), .D ( n2765 ), .Q ( new_AGEMA_signal_5369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C ( clk ), .D ( new_AGEMA_signal_957 ), .Q ( new_AGEMA_signal_5370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C ( clk ), .D ( n2791 ), .Q ( new_AGEMA_signal_5371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C ( clk ), .D ( new_AGEMA_signal_951 ), .Q ( new_AGEMA_signal_5372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_5373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_5374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C ( clk ), .D ( n2813 ), .Q ( new_AGEMA_signal_5375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C ( clk ), .D ( new_AGEMA_signal_953 ), .Q ( new_AGEMA_signal_5376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C ( clk ), .D ( n2810 ), .Q ( new_AGEMA_signal_5377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C ( clk ), .D ( new_AGEMA_signal_945 ), .Q ( new_AGEMA_signal_5378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_5635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_5638 ) ) ;

    /* cells in depth 2 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1954 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ({Fresh[211], Fresh[210], Fresh[209], Fresh[208]}), .c ({new_AGEMA_signal_1127, n2575}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1959 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212]}), .c ({new_AGEMA_signal_1128, n1962}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1964 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ({Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1129, n1922}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1974 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ({Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .c ({new_AGEMA_signal_1030, n2755}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1977 ( .a ({new_AGEMA_signal_977, n2317}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224]}), .c ({new_AGEMA_signal_1130, n1926}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1980 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1032, n2541}), .clk ( clk ), .r ({Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1131, n1925}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1986 ( .a ({new_AGEMA_signal_1033, n2086}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ({Fresh[235], Fresh[234], Fresh[233], Fresh[232]}), .c ({new_AGEMA_signal_1132, n2151}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1988 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236]}), .c ({new_AGEMA_signal_1034, n2631}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U1989 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_1133, n2734}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1992 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ({Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1134, n2763}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1997 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ({Fresh[247], Fresh[246], Fresh[245], Fresh[244]}), .c ({new_AGEMA_signal_1036, n1930}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2005 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248]}), .c ({new_AGEMA_signal_1038, n2492}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2006 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1135, n2732}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2010 ( .a ({new_AGEMA_signal_5350, new_AGEMA_signal_5349}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ({Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1136, n1937}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2022 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5351}), .b ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .r ({Fresh[259], Fresh[258], Fresh[257], Fresh[256]}), .c ({new_AGEMA_signal_1042, n1942}) ) ;
    or_GHPC #(.low_latency(1), .pipeline(1)) U2026 ( .a ({new_AGEMA_signal_993, n2587}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .c ({new_AGEMA_signal_1043, n2676}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2030 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ({Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1139, n1944}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2037 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ({Fresh[271], Fresh[270], Fresh[269], Fresh[268]}), .c ({new_AGEMA_signal_1140, n1950}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2039 ( .a ({new_AGEMA_signal_5354, new_AGEMA_signal_5353}), .b ({new_AGEMA_signal_995, n2739}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272]}), .c ({new_AGEMA_signal_1046, n1949}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2042 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ({Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1047, n2677}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2043 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1141, n2662}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2047 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ({Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .c ({new_AGEMA_signal_1048, n2627}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2053 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_998, n2452}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284]}), .c ({new_AGEMA_signal_1049, n1957}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2056 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ({Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1142, n2088}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2062 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ({Fresh[295], Fresh[294], Fresh[293], Fresh[292]}), .c ({new_AGEMA_signal_999, n1964}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2063 ( .a ({new_AGEMA_signal_5356, new_AGEMA_signal_5355}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296]}), .c ({new_AGEMA_signal_1051, n2736}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2069 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_5358, new_AGEMA_signal_5357}), .clk ( clk ), .r ({Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1052, n2673}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2072 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ({Fresh[307], Fresh[306], Fresh[305], Fresh[304]}), .c ({new_AGEMA_signal_1144, n2761}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2073 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1323, n2720}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2075 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308]}), .c ({new_AGEMA_signal_1145, n2412}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2076 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_1324, n2417}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2079 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_966, n2261}), .clk ( clk ), .r ({Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1055, n2571}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2080 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1146, n2505}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2081 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316]}), .c ({new_AGEMA_signal_1056, n2651}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2083 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_5358, new_AGEMA_signal_5357}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .c ({new_AGEMA_signal_1147, n2359}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2086 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ({Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1057, n2101}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2087 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1148, n2625}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2091 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ({Fresh[331], Fresh[330], Fresh[329], Fresh[328]}), .c ({new_AGEMA_signal_1059, n2190}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2095 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332]}), .c ({new_AGEMA_signal_1060, n1976}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2098 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ({Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1150, n2535}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2101 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .r ({Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .c ({new_AGEMA_signal_1151, n1973}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2105 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344]}), .c ({new_AGEMA_signal_1061, n2690}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2111 ( .a ({new_AGEMA_signal_992, n2493}), .b ({new_AGEMA_signal_5360, new_AGEMA_signal_5359}), .clk ( clk ), .r ({Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1062, n2817}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2113 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ({Fresh[355], Fresh[354], Fresh[353], Fresh[352]}), .c ({new_AGEMA_signal_1153, n2741}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2118 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356]}), .c ({new_AGEMA_signal_1154, n1992}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2120 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ({Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1155, n1991}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2123 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ({Fresh[367], Fresh[366], Fresh[365], Fresh[364]}), .c ({new_AGEMA_signal_1064, n1993}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2125 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368]}), .c ({new_AGEMA_signal_1156, n1995}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2132 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ({Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1157, n2241}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2135 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361}), .b ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .r ({Fresh[379], Fresh[378], Fresh[377], Fresh[376]}), .c ({new_AGEMA_signal_1158, n2003}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2140 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .c ({new_AGEMA_signal_1159, n2008}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2141 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ({Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1160, n2572}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2143 ( .a ({new_AGEMA_signal_1067, n2809}), .b ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .r ({Fresh[391], Fresh[390], Fresh[389], Fresh[388]}), .c ({new_AGEMA_signal_1161, n2004}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2147 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392]}), .c ({new_AGEMA_signal_1162, n2009}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2151 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_5360, new_AGEMA_signal_5359}), .clk ( clk ), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1163, n2533}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2157 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ({Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .c ({new_AGEMA_signal_1069, n2026}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2158 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404]}), .c ({new_AGEMA_signal_1164, n2022}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2159 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ({Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1070, n2227}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2167 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_5360, new_AGEMA_signal_5359}), .clk ( clk ), .r ({Fresh[415], Fresh[414], Fresh[413], Fresh[412]}), .c ({new_AGEMA_signal_1009, n2027}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2171 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416]}), .c ({new_AGEMA_signal_1167, n2214}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2173 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1168, n2290}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2174 ( .a ({new_AGEMA_signal_5356, new_AGEMA_signal_5355}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ({Fresh[427], Fresh[426], Fresh[425], Fresh[424]}), .c ({new_AGEMA_signal_1169, n2376}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2178 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428]}), .c ({new_AGEMA_signal_1072, n2034}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2182 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ({Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1073, n2171}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2183 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ({Fresh[439], Fresh[438], Fresh[437], Fresh[436]}), .c ({new_AGEMA_signal_1170, n2039}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2188 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440]}), .c ({new_AGEMA_signal_1172, n2042}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2191 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ({Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1173, n2754}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2192 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_959, n2790}), .clk ( clk ), .r ({Fresh[451], Fresh[450], Fresh[449], Fresh[448]}), .c ({new_AGEMA_signal_1174, n2044}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2198 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452]}), .c ({new_AGEMA_signal_1175, n2654}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2202 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1037, n2577}), .clk ( clk ), .r ({Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1176, n2055}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2205 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ({Fresh[463], Fresh[462], Fresh[461], Fresh[460]}), .c ({new_AGEMA_signal_1177, n2057}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2208 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464]}), .c ({new_AGEMA_signal_1178, n2407}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2212 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1010, n2061}), .clk ( clk ), .r ({Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1179, n2062}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2216 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ({Fresh[475], Fresh[474], Fresh[473], Fresh[472]}), .c ({new_AGEMA_signal_1180, n2731}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2220 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1181, n2068}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2224 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476]}), .c ({new_AGEMA_signal_1074, n2642}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2225 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ({Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1182, n2252}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2228 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ({Fresh[487], Fresh[486], Fresh[485], Fresh[484]}), .c ({new_AGEMA_signal_1075, n2075}) ) ;
    or_GHPC #(.low_latency(1), .pipeline(1)) U2233 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488]}), .c ({new_AGEMA_signal_1076, n2081}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2234 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ({Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1183, n2080}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2237 ( .a ({new_AGEMA_signal_984, n2600}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ({Fresh[499], Fresh[498], Fresh[497], Fresh[496]}), .c ({new_AGEMA_signal_1077, n2498}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2238 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_1184, n2773}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2239 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500]}), .c ({new_AGEMA_signal_1185, n2083}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2244 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361}), .b ({new_AGEMA_signal_1033, n2086}), .clk ( clk ), .r ({Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1186, n2562}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2247 ( .a ({new_AGEMA_signal_5356, new_AGEMA_signal_5355}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ({Fresh[511], Fresh[510], Fresh[509], Fresh[508]}), .c ({new_AGEMA_signal_1078, n2087}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2251 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1041, n2174}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512]}), .c ({new_AGEMA_signal_1187, n2156}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2260 ( .a ({new_AGEMA_signal_1028, n2769}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ({Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1188, n2100}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2277 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_1012, n2298}), .clk ( clk ), .r ({Fresh[523], Fresh[522], Fresh[521], Fresh[520]}), .c ({new_AGEMA_signal_1079, n2544}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2279 ( .a ({new_AGEMA_signal_1004, n2356}), .b ({new_AGEMA_signal_1080, n2118}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524]}), .c ({new_AGEMA_signal_1191, n2121}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2284 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ({Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1193, n2122}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2286 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ({Fresh[535], Fresh[534], Fresh[533], Fresh[532]}), .c ({new_AGEMA_signal_1194, n2811}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2294 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536]}), .c ({new_AGEMA_signal_1081, n2647}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2297 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ({Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1082, n2132}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2304 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[547], Fresh[546], Fresh[545], Fresh[544]}), .c ({new_AGEMA_signal_1199, n2220}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2305 ( .a ({new_AGEMA_signal_5350, new_AGEMA_signal_5349}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548]}), .c ({new_AGEMA_signal_1200, n2138}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2312 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_5366, new_AGEMA_signal_5365}), .clk ( clk ), .r ({Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1201, n2555}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2322 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367}), .clk ( clk ), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556]}), .c ({new_AGEMA_signal_1202, n2429}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2328 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_5360, new_AGEMA_signal_5359}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .c ({new_AGEMA_signal_1083, n2162}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2337 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ({Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1014, n2545}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2340 ( .a ({new_AGEMA_signal_965, n2559}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ({Fresh[571], Fresh[570], Fresh[569], Fresh[568]}), .c ({new_AGEMA_signal_1085, n2178}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2342 ( .a ({new_AGEMA_signal_1015, n2430}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572]}), .c ({new_AGEMA_signal_1204, n2176}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2343 ( .a ({new_AGEMA_signal_1041, n2174}), .b ({new_AGEMA_signal_5362, new_AGEMA_signal_5361}), .clk ( clk ), .r ({Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1205, n2175}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2348 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367}), .clk ( clk ), .r ({Fresh[583], Fresh[582], Fresh[581], Fresh[580]}), .c ({new_AGEMA_signal_1016, n2182}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2353 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584]}), .c ({new_AGEMA_signal_1206, n2188}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2355 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ({Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1207, n2189}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2357 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ({Fresh[595], Fresh[594], Fresh[593], Fresh[592]}), .c ({new_AGEMA_signal_1208, n2446}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2362 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596]}), .c ({new_AGEMA_signal_1087, n2576}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2363 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_5370, new_AGEMA_signal_5369}), .clk ( clk ), .r ({Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1088, n2748}) ) ;
    not_masked #(.low_latency(1), .pipeline(1)) U2368 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_1375, n2674}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2378 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ({Fresh[607], Fresh[606], Fresh[605], Fresh[604]}), .c ({new_AGEMA_signal_1089, n2213}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2380 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_5356, new_AGEMA_signal_5355}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608]}), .c ({new_AGEMA_signal_1090, n2215}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2384 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ({Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1211, n2218}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2386 ( .a ({new_AGEMA_signal_1012, n2298}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ({Fresh[619], Fresh[618], Fresh[617], Fresh[616]}), .c ({new_AGEMA_signal_1212, n2219}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2405 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620]}), .c ({new_AGEMA_signal_1217, n2240}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2407 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ({Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1218, n2561}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2408 ( .a ({new_AGEMA_signal_5362, new_AGEMA_signal_5361}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ({Fresh[631], Fresh[630], Fresh[629], Fresh[628]}), .c ({new_AGEMA_signal_1219, n2243}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2411 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632]}), .c ({new_AGEMA_signal_1220, n2245}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2422 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1221, n2540}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2423 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ({Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .c ({new_AGEMA_signal_1222, n2259}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2426 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644]}), .c ({new_AGEMA_signal_1091, n2262}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2431 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ({Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1092, n2266}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2432 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_5368, new_AGEMA_signal_5367}), .clk ( clk ), .r ({Fresh[655], Fresh[654], Fresh[653], Fresh[652]}), .c ({new_AGEMA_signal_1093, n2645}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2436 ( .a ({new_AGEMA_signal_5350, new_AGEMA_signal_5349}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656]}), .c ({new_AGEMA_signal_1094, n2268}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2443 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ({Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1225, n2278}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2448 ( .a ({new_AGEMA_signal_5372, new_AGEMA_signal_5371}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ({Fresh[667], Fresh[666], Fresh[665], Fresh[664]}), .c ({new_AGEMA_signal_1095, n2383}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2455 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668]}), .c ({new_AGEMA_signal_1228, n2774}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2458 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ({Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1229, n2287}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2470 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[679], Fresh[678], Fresh[677], Fresh[676]}), .c ({new_AGEMA_signal_1231, n2438}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2471 ( .a ({new_AGEMA_signal_1012, n2298}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680]}), .c ({new_AGEMA_signal_1096, n2299}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2481 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1054, n2313}), .clk ( clk ), .r ({Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1232, n2371}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2484 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ({Fresh[691], Fresh[690], Fresh[689], Fresh[688]}), .c ({new_AGEMA_signal_1018, n2316}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2486 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692]}), .c ({new_AGEMA_signal_1098, n2318}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2492 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ({Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1235, n2325}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2494 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[703], Fresh[702], Fresh[701], Fresh[700]}), .c ({new_AGEMA_signal_1236, n2328}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2495 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704]}), .c ({new_AGEMA_signal_1099, n2327}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2505 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .r ({Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1237, n2343}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2510 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ({Fresh[715], Fresh[714], Fresh[713], Fresh[712]}), .c ({new_AGEMA_signal_1239, n2344}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) U2512 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1013, n2346}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716]}), .c ({new_AGEMA_signal_1100, n2348}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2513 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ({Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1101, n2347}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2520 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ({Fresh[727], Fresh[726], Fresh[725], Fresh[724]}), .c ({new_AGEMA_signal_1102, n2363}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2521 ( .a ({new_AGEMA_signal_1067, n2809}), .b ({new_AGEMA_signal_5358, new_AGEMA_signal_5357}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728]}), .c ({new_AGEMA_signal_1243, n2353}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2524 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ({Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1244, n2355}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2530 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ({Fresh[739], Fresh[738], Fresh[737], Fresh[736]}), .c ({new_AGEMA_signal_1245, n2364}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2543 ( .a ({new_AGEMA_signal_5350, new_AGEMA_signal_5349}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740]}), .c ({new_AGEMA_signal_1103, n2415}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2558 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ({Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1104, n2700}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2563 ( .a ({new_AGEMA_signal_5374, new_AGEMA_signal_5373}), .b ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .r ({Fresh[751], Fresh[750], Fresh[749], Fresh[748]}), .c ({new_AGEMA_signal_1105, n2594}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2564 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_5360, new_AGEMA_signal_5359}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752]}), .c ({new_AGEMA_signal_1106, n2402}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2585 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ({Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1255, n2428}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2588 ( .a ({new_AGEMA_signal_1015, n2430}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ({Fresh[763], Fresh[762], Fresh[761], Fresh[760]}), .c ({new_AGEMA_signal_1256, n2431}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2594 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764]}), .c ({new_AGEMA_signal_1107, n2483}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2599 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ({Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1258, n2443}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2606 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ({Fresh[775], Fresh[774], Fresh[773], Fresh[772]}), .c ({new_AGEMA_signal_1259, n2693}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2608 ( .a ({new_AGEMA_signal_998, n2452}), .b ({new_AGEMA_signal_5376, new_AGEMA_signal_5375}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776]}), .c ({new_AGEMA_signal_1108, n2453}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2616 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1019, n2463}), .clk ( clk ), .r ({Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1109, n2464}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2620 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ({Fresh[787], Fresh[786], Fresh[785], Fresh[784]}), .c ({new_AGEMA_signal_1110, n2468}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2624 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_5358, new_AGEMA_signal_5357}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788]}), .c ({new_AGEMA_signal_1111, n2473}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2625 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ({Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1112, n2472}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2628 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1020, n2474}), .clk ( clk ), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796]}), .c ({new_AGEMA_signal_1113, n2475}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2632 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377}), .b ({new_AGEMA_signal_1065, n2828}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .c ({new_AGEMA_signal_1263, n2480}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2638 ( .a ({new_AGEMA_signal_1037, n2577}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ({Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1264, n2487}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2641 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ({Fresh[811], Fresh[810], Fresh[809], Fresh[808]}), .c ({new_AGEMA_signal_1114, n2488}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2665 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812]}), .c ({new_AGEMA_signal_1270, n2520}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2667 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_993, n2587}), .clk ( clk ), .r ({Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1115, n2521}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2674 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_963, n2595}), .clk ( clk ), .r ({Fresh[823], Fresh[822], Fresh[821], Fresh[820]}), .c ({new_AGEMA_signal_1271, n2531}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2689 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824]}), .c ({new_AGEMA_signal_1273, n2553}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2691 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ({Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1274, n2554}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) U2695 ( .a ({new_AGEMA_signal_965, n2559}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ({Fresh[835], Fresh[834], Fresh[833], Fresh[832]}), .c ({new_AGEMA_signal_1116, n2560}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2698 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836]}), .c ({new_AGEMA_signal_1275, n2564}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2714 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .r ({Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_1278, n2586}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2720 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ({Fresh[847], Fresh[846], Fresh[845], Fresh[844]}), .c ({new_AGEMA_signal_1117, n2597}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2721 ( .a ({new_AGEMA_signal_1024, n2640}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848]}), .c ({new_AGEMA_signal_1280, n2596}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2723 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ({Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_1281, n2598}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2725 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_5356, new_AGEMA_signal_5355}), .clk ( clk ), .r ({Fresh[859], Fresh[858], Fresh[857], Fresh[856]}), .c ({new_AGEMA_signal_1021, n2599}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2732 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860]}), .c ({new_AGEMA_signal_1283, n2610}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2734 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ({Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_1284, n2614}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2735 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ({Fresh[871], Fresh[870], Fresh[869], Fresh[868]}), .c ({new_AGEMA_signal_1285, n2613}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2737 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872]}), .c ({new_AGEMA_signal_1119, n2617}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2742 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_1120, n2629}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2751 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ({Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .c ({new_AGEMA_signal_1287, n2784}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2757 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884]}), .c ({new_AGEMA_signal_1121, n2650}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2775 ( .a ({new_AGEMA_signal_5366, new_AGEMA_signal_5365}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ({Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_1022, n2683}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2789 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ({Fresh[895], Fresh[894], Fresh[893], Fresh[892]}), .c ({new_AGEMA_signal_1294, n2711}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2790 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896]}), .c ({new_AGEMA_signal_1295, n2710}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2792 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_969, n2712}), .clk ( clk ), .r ({Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_1122, n2714}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2797 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1011, n2721}), .clk ( clk ), .r ({Fresh[907], Fresh[906], Fresh[905], Fresh[904]}), .c ({new_AGEMA_signal_1123, n2722}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2799 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908]}), .c ({new_AGEMA_signal_1297, n2726}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2806 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ({Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_1298, n2738}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2822 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .r ({Fresh[919], Fresh[918], Fresh[917], Fresh[916]}), .c ({new_AGEMA_signal_1301, n2768}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2828 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920]}), .c ({new_AGEMA_signal_1124, n2782}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2829 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ({Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_1125, n2781}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2832 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_989, n2785}), .clk ( clk ), .r ({Fresh[931], Fresh[930], Fresh[929], Fresh[928]}), .c ({new_AGEMA_signal_1303, n2787}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2834 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932]}), .c ({new_AGEMA_signal_1304, n2794}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2835 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_5372, new_AGEMA_signal_5371}), .clk ( clk ), .r ({Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_1305, n2793}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2844 ( .a ({new_AGEMA_signal_5378, new_AGEMA_signal_5377}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ({Fresh[943], Fresh[942], Fresh[941], Fresh[940]}), .c ({new_AGEMA_signal_1306, n2812}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2847 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944]}), .c ({new_AGEMA_signal_1126, n2820}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2851 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ({Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_1308, n2825}) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C ( clk ), .D ( n2769 ), .Q ( new_AGEMA_signal_5379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_5380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C ( clk ), .D ( new_AGEMA_signal_5373 ), .Q ( new_AGEMA_signal_5381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C ( clk ), .D ( new_AGEMA_signal_5374 ), .Q ( new_AGEMA_signal_5382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C ( clk ), .D ( new_AGEMA_signal_5351 ), .Q ( new_AGEMA_signal_5383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C ( clk ), .D ( new_AGEMA_signal_5352 ), .Q ( new_AGEMA_signal_5384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C ( clk ), .D ( n2174 ), .Q ( new_AGEMA_signal_5385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C ( clk ), .D ( new_AGEMA_signal_1041 ), .Q ( new_AGEMA_signal_5386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C ( clk ), .D ( new_AGEMA_signal_5349 ), .Q ( new_AGEMA_signal_5387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C ( clk ), .D ( new_AGEMA_signal_5350 ), .Q ( new_AGEMA_signal_5388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C ( clk ), .D ( new_AGEMA_signal_5355 ), .Q ( new_AGEMA_signal_5389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C ( clk ), .D ( new_AGEMA_signal_5356 ), .Q ( new_AGEMA_signal_5390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C ( clk ), .D ( n2570 ), .Q ( new_AGEMA_signal_5391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_5392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C ( clk ), .D ( n2792 ), .Q ( new_AGEMA_signal_5393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C ( clk ), .D ( new_AGEMA_signal_1039 ), .Q ( new_AGEMA_signal_5394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C ( clk ), .D ( n2635 ), .Q ( new_AGEMA_signal_5395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C ( clk ), .D ( new_AGEMA_signal_958 ), .Q ( new_AGEMA_signal_5396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C ( clk ), .D ( n2587 ), .Q ( new_AGEMA_signal_5397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C ( clk ), .D ( new_AGEMA_signal_993 ), .Q ( new_AGEMA_signal_5398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C ( clk ), .D ( n2725 ), .Q ( new_AGEMA_signal_5399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C ( clk ), .D ( new_AGEMA_signal_982 ), .Q ( new_AGEMA_signal_5400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C ( clk ), .D ( n2708 ), .Q ( new_AGEMA_signal_5401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_5402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C ( clk ), .D ( n2818 ), .Q ( new_AGEMA_signal_5403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_5404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C ( clk ), .D ( n2790 ), .Q ( new_AGEMA_signal_5405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C ( clk ), .D ( new_AGEMA_signal_959 ), .Q ( new_AGEMA_signal_5406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C ( clk ), .D ( n2786 ), .Q ( new_AGEMA_signal_5407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C ( clk ), .D ( new_AGEMA_signal_1035 ), .Q ( new_AGEMA_signal_5408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C ( clk ), .D ( n2400 ), .Q ( new_AGEMA_signal_5409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C ( clk ), .D ( new_AGEMA_signal_988 ), .Q ( new_AGEMA_signal_5410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C ( clk ), .D ( new_AGEMA_signal_5357 ), .Q ( new_AGEMA_signal_5411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C ( clk ), .D ( new_AGEMA_signal_5358 ), .Q ( new_AGEMA_signal_5412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C ( clk ), .D ( n2815 ), .Q ( new_AGEMA_signal_5413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C ( clk ), .D ( new_AGEMA_signal_983 ), .Q ( new_AGEMA_signal_5414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C ( clk ), .D ( n2723 ), .Q ( new_AGEMA_signal_5415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C ( clk ), .D ( new_AGEMA_signal_981 ), .Q ( new_AGEMA_signal_5416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C ( clk ), .D ( n2709 ), .Q ( new_AGEMA_signal_5417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_5418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C ( clk ), .D ( n2753 ), .Q ( new_AGEMA_signal_5419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C ( clk ), .D ( new_AGEMA_signal_987 ), .Q ( new_AGEMA_signal_5420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C ( clk ), .D ( n2401 ), .Q ( new_AGEMA_signal_5421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_5422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C ( clk ), .D ( new_AGEMA_signal_5369 ), .Q ( new_AGEMA_signal_5423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C ( clk ), .D ( new_AGEMA_signal_5370 ), .Q ( new_AGEMA_signal_5424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C ( clk ), .D ( new_AGEMA_signal_5359 ), .Q ( new_AGEMA_signal_5425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C ( clk ), .D ( new_AGEMA_signal_5360 ), .Q ( new_AGEMA_signal_5426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C ( clk ), .D ( n2615 ), .Q ( new_AGEMA_signal_5427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C ( clk ), .D ( new_AGEMA_signal_973 ), .Q ( new_AGEMA_signal_5428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C ( clk ), .D ( n2643 ), .Q ( new_AGEMA_signal_5429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C ( clk ), .D ( new_AGEMA_signal_994 ), .Q ( new_AGEMA_signal_5430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C ( clk ), .D ( n2563 ), .Q ( new_AGEMA_signal_5431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_5432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C ( clk ), .D ( n2612 ), .Q ( new_AGEMA_signal_5433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C ( clk ), .D ( new_AGEMA_signal_1053 ), .Q ( new_AGEMA_signal_5434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C ( clk ), .D ( n2824 ), .Q ( new_AGEMA_signal_5435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C ( clk ), .D ( new_AGEMA_signal_1001 ), .Q ( new_AGEMA_signal_5436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C ( clk ), .D ( n2816 ), .Q ( new_AGEMA_signal_5437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C ( clk ), .D ( new_AGEMA_signal_975 ), .Q ( new_AGEMA_signal_5438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C ( clk ), .D ( n2073 ), .Q ( new_AGEMA_signal_5439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C ( clk ), .D ( new_AGEMA_signal_979 ), .Q ( new_AGEMA_signal_5440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C ( clk ), .D ( n2519 ), .Q ( new_AGEMA_signal_5441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C ( clk ), .D ( new_AGEMA_signal_960 ), .Q ( new_AGEMA_signal_5442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C ( clk ), .D ( n2616 ), .Q ( new_AGEMA_signal_5443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_5444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C ( clk ), .D ( new_AGEMA_signal_5371 ), .Q ( new_AGEMA_signal_5445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C ( clk ), .D ( new_AGEMA_signal_5372 ), .Q ( new_AGEMA_signal_5446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C ( clk ), .D ( n2780 ), .Q ( new_AGEMA_signal_5447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C ( clk ), .D ( new_AGEMA_signal_976 ), .Q ( new_AGEMA_signal_5448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C ( clk ), .D ( new_AGEMA_signal_5375 ), .Q ( new_AGEMA_signal_5449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C ( clk ), .D ( new_AGEMA_signal_5376 ), .Q ( new_AGEMA_signal_5450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C ( clk ), .D ( n2742 ), .Q ( new_AGEMA_signal_5451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C ( clk ), .D ( new_AGEMA_signal_986 ), .Q ( new_AGEMA_signal_5452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C ( clk ), .D ( n2724 ), .Q ( new_AGEMA_signal_5453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C ( clk ), .D ( new_AGEMA_signal_1040 ), .Q ( new_AGEMA_signal_5454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C ( clk ), .D ( n2317 ), .Q ( new_AGEMA_signal_5455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C ( clk ), .D ( new_AGEMA_signal_977 ), .Q ( new_AGEMA_signal_5456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C ( clk ), .D ( n2688 ), .Q ( new_AGEMA_signal_5457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_5458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C ( clk ), .D ( n2609 ), .Q ( new_AGEMA_signal_5459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C ( clk ), .D ( new_AGEMA_signal_990 ), .Q ( new_AGEMA_signal_5460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C ( clk ), .D ( n2672 ), .Q ( new_AGEMA_signal_5461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C ( clk ), .D ( new_AGEMA_signal_1023 ), .Q ( new_AGEMA_signal_5462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C ( clk ), .D ( n2640 ), .Q ( new_AGEMA_signal_5463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C ( clk ), .D ( new_AGEMA_signal_1024 ), .Q ( new_AGEMA_signal_5464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C ( clk ), .D ( n2713 ), .Q ( new_AGEMA_signal_5465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C ( clk ), .D ( new_AGEMA_signal_980 ), .Q ( new_AGEMA_signal_5466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C ( clk ), .D ( n2777 ), .Q ( new_AGEMA_signal_5467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C ( clk ), .D ( new_AGEMA_signal_1017 ), .Q ( new_AGEMA_signal_5468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C ( clk ), .D ( n2789 ), .Q ( new_AGEMA_signal_5469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_5470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C ( clk ), .D ( n2661 ), .Q ( new_AGEMA_signal_5471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C ( clk ), .D ( new_AGEMA_signal_991 ), .Q ( new_AGEMA_signal_5472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C ( clk ), .D ( new_AGEMA_signal_5363 ), .Q ( new_AGEMA_signal_5473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C ( clk ), .D ( new_AGEMA_signal_5364 ), .Q ( new_AGEMA_signal_5474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C ( clk ), .D ( n2694 ), .Q ( new_AGEMA_signal_5475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C ( clk ), .D ( new_AGEMA_signal_978 ), .Q ( new_AGEMA_signal_5476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C ( clk ), .D ( new_AGEMA_signal_5365 ), .Q ( new_AGEMA_signal_5477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C ( clk ), .D ( new_AGEMA_signal_5366 ), .Q ( new_AGEMA_signal_5478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C ( clk ), .D ( n2682 ), .Q ( new_AGEMA_signal_5479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C ( clk ), .D ( new_AGEMA_signal_962 ), .Q ( new_AGEMA_signal_5480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C ( clk ), .D ( new_AGEMA_signal_5377 ), .Q ( new_AGEMA_signal_5481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C ( clk ), .D ( new_AGEMA_signal_5378 ), .Q ( new_AGEMA_signal_5482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C ( clk ), .D ( n2624 ), .Q ( new_AGEMA_signal_5483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_5484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C ( clk ), .D ( n2356 ), .Q ( new_AGEMA_signal_5485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_5486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C ( clk ), .D ( n2778 ), .Q ( new_AGEMA_signal_5487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C ( clk ), .D ( new_AGEMA_signal_997 ), .Q ( new_AGEMA_signal_5488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C ( clk ), .D ( n2766 ), .Q ( new_AGEMA_signal_5489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C ( clk ), .D ( new_AGEMA_signal_1050 ), .Q ( new_AGEMA_signal_5490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C ( clk ), .D ( n2767 ), .Q ( new_AGEMA_signal_5491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_5492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C ( clk ), .D ( n2641 ), .Q ( new_AGEMA_signal_5493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C ( clk ), .D ( new_AGEMA_signal_971 ), .Q ( new_AGEMA_signal_5494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C ( clk ), .D ( n2719 ), .Q ( new_AGEMA_signal_5495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C ( clk ), .D ( new_AGEMA_signal_970 ), .Q ( new_AGEMA_signal_5496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C ( clk ), .D ( n2707 ), .Q ( new_AGEMA_signal_5497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C ( clk ), .D ( new_AGEMA_signal_1029 ), .Q ( new_AGEMA_signal_5498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C ( clk ), .D ( n2493 ), .Q ( new_AGEMA_signal_5499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C ( clk ), .D ( new_AGEMA_signal_992 ), .Q ( new_AGEMA_signal_5500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C ( clk ), .D ( n2577 ), .Q ( new_AGEMA_signal_5501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C ( clk ), .D ( new_AGEMA_signal_1037 ), .Q ( new_AGEMA_signal_5502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C ( clk ), .D ( n2541 ), .Q ( new_AGEMA_signal_5503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_5504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C ( clk ), .D ( n2679 ), .Q ( new_AGEMA_signal_5505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_5506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C ( clk ), .D ( n2699 ), .Q ( new_AGEMA_signal_5507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C ( clk ), .D ( new_AGEMA_signal_974 ), .Q ( new_AGEMA_signal_5508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C ( clk ), .D ( n2611 ), .Q ( new_AGEMA_signal_5509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C ( clk ), .D ( new_AGEMA_signal_1005 ), .Q ( new_AGEMA_signal_5510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C ( clk ), .D ( n2739 ), .Q ( new_AGEMA_signal_5511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C ( clk ), .D ( new_AGEMA_signal_995 ), .Q ( new_AGEMA_signal_5512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C ( clk ), .D ( n2772 ), .Q ( new_AGEMA_signal_5513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C ( clk ), .D ( new_AGEMA_signal_1000 ), .Q ( new_AGEMA_signal_5514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C ( clk ), .D ( n2442 ), .Q ( new_AGEMA_signal_5519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_5521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C ( clk ), .D ( n2779 ), .Q ( new_AGEMA_signal_5545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C ( clk ), .D ( new_AGEMA_signal_967 ), .Q ( new_AGEMA_signal_5547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C ( clk ), .D ( n2721 ), .Q ( new_AGEMA_signal_5563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C ( clk ), .D ( new_AGEMA_signal_1011 ), .Q ( new_AGEMA_signal_5565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C ( clk ), .D ( n2823 ), .Q ( new_AGEMA_signal_5577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C ( clk ), .D ( new_AGEMA_signal_1063 ), .Q ( new_AGEMA_signal_5579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C ( clk ), .D ( n2346 ), .Q ( new_AGEMA_signal_5587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C ( clk ), .D ( new_AGEMA_signal_1013 ), .Q ( new_AGEMA_signal_5589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C ( clk ), .D ( n2315 ), .Q ( new_AGEMA_signal_5597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C ( clk ), .D ( new_AGEMA_signal_961 ), .Q ( new_AGEMA_signal_5599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C ( clk ), .D ( new_AGEMA_signal_5635 ), .Q ( new_AGEMA_signal_5636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C ( clk ), .D ( new_AGEMA_signal_5638 ), .Q ( new_AGEMA_signal_5639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C ( clk ), .D ( new_AGEMA_signal_5353 ), .Q ( new_AGEMA_signal_5647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C ( clk ), .D ( new_AGEMA_signal_5354 ), .Q ( new_AGEMA_signal_5649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C ( clk ), .D ( n2600 ), .Q ( new_AGEMA_signal_5657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C ( clk ), .D ( new_AGEMA_signal_984 ), .Q ( new_AGEMA_signal_5659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C ( clk ), .D ( n2750 ), .Q ( new_AGEMA_signal_5675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C ( clk ), .D ( new_AGEMA_signal_972 ), .Q ( new_AGEMA_signal_5677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C ( clk ), .D ( new_AGEMA_signal_5367 ), .Q ( new_AGEMA_signal_5683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C ( clk ), .D ( new_AGEMA_signal_5368 ), .Q ( new_AGEMA_signal_5685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C ( clk ), .D ( n2737 ), .Q ( new_AGEMA_signal_5757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C ( clk ), .D ( new_AGEMA_signal_1025 ), .Q ( new_AGEMA_signal_5760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C ( clk ), .D ( n2785 ), .Q ( new_AGEMA_signal_5783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C ( clk ), .D ( new_AGEMA_signal_989 ), .Q ( new_AGEMA_signal_5786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C ( clk ), .D ( n2595 ), .Q ( new_AGEMA_signal_5899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C ( clk ), .D ( new_AGEMA_signal_963 ), .Q ( new_AGEMA_signal_5903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C ( clk ), .D ( n2437 ), .Q ( new_AGEMA_signal_5909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C ( clk ), .D ( new_AGEMA_signal_996 ), .Q ( new_AGEMA_signal_5913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C ( clk ), .D ( n2828 ), .Q ( new_AGEMA_signal_5985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C ( clk ), .D ( new_AGEMA_signal_1065 ), .Q ( new_AGEMA_signal_5989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C ( clk ), .D ( n2538 ), .Q ( new_AGEMA_signal_6071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C ( clk ), .D ( new_AGEMA_signal_985 ), .Q ( new_AGEMA_signal_6075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C ( clk ), .D ( n2809 ), .Q ( new_AGEMA_signal_6101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_6105 ) ) ;

    /* cells in depth 3 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1960 ( .a ({new_AGEMA_signal_1127, n2575}), .b ({new_AGEMA_signal_1128, n1962}), .clk ( clk ), .r ({Fresh[955], Fresh[954], Fresh[953], Fresh[952]}), .c ({new_AGEMA_signal_1309, n1924}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1967 ( .a ({new_AGEMA_signal_1129, n1922}), .b ({new_AGEMA_signal_5380, new_AGEMA_signal_5379}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956]}), .c ({new_AGEMA_signal_1310, n1923}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1981 ( .a ({new_AGEMA_signal_1130, n1926}), .b ({new_AGEMA_signal_1131, n1925}), .clk ( clk ), .r ({Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_1311, n1927}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1993 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_1134, n2763}), .clk ( clk ), .r ({Fresh[967], Fresh[966], Fresh[965], Fresh[964]}), .c ({new_AGEMA_signal_1312, n1929}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2007 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968]}), .c ({new_AGEMA_signal_1313, n2665}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2011 ( .a ({new_AGEMA_signal_5384, new_AGEMA_signal_5383}), .b ({new_AGEMA_signal_1136, n1937}), .clk ( clk ), .r ({Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_1314, n1938}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2019 ( .a ({new_AGEMA_signal_5386, new_AGEMA_signal_5385}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ({Fresh[979], Fresh[978], Fresh[977], Fresh[976]}), .c ({new_AGEMA_signal_1315, n2235}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2023 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387}), .b ({new_AGEMA_signal_1042, n1942}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980]}), .c ({new_AGEMA_signal_1137, n1943}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2027 ( .a ({new_AGEMA_signal_1043, n2676}), .b ({new_AGEMA_signal_5390, new_AGEMA_signal_5389}), .clk ( clk ), .r ({Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_1138, n1946}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2031 ( .a ({new_AGEMA_signal_5392, new_AGEMA_signal_5391}), .b ({new_AGEMA_signal_1139, n1944}), .clk ( clk ), .r ({Fresh[991], Fresh[990], Fresh[989], Fresh[988]}), .c ({new_AGEMA_signal_1316, n1945}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2034 ( .a ({new_AGEMA_signal_5394, new_AGEMA_signal_5393}), .b ({new_AGEMA_signal_1133, n2734}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992]}), .c ({new_AGEMA_signal_1317, n1956}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2040 ( .a ({new_AGEMA_signal_1140, n1950}), .b ({new_AGEMA_signal_1046, n1949}), .clk ( clk ), .r ({Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_1318, n1951}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2048 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ({Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000]}), .c ({new_AGEMA_signal_1319, n1952}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2057 ( .a ({new_AGEMA_signal_5396, new_AGEMA_signal_5395}), .b ({new_AGEMA_signal_1142, n2088}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004]}), .c ({new_AGEMA_signal_1320, n2687}) ) ;
    or_GHPC #(.low_latency(1), .pipeline(1)) U2061 ( .a ({new_AGEMA_signal_1128, n1962}), .b ({new_AGEMA_signal_5398, new_AGEMA_signal_5397}), .clk ( clk ), .r ({Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_1321, n1966}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2064 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_5400, new_AGEMA_signal_5399}), .clk ( clk ), .r ({Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012]}), .c ({new_AGEMA_signal_1143, n1963}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2077 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016]}), .c ({new_AGEMA_signal_1480, n1968}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2082 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_1325, n2684}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2088 ( .a ({new_AGEMA_signal_5402, new_AGEMA_signal_5401}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ({Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024]}), .c ({new_AGEMA_signal_1326, n1972}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2092 ( .a ({new_AGEMA_signal_5404, new_AGEMA_signal_5403}), .b ({new_AGEMA_signal_1059, n2190}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028]}), .c ({new_AGEMA_signal_1149, n1971}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2099 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405}), .b ({new_AGEMA_signal_1150, n2535}), .clk ( clk ), .r ({Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_1327, n1974}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2106 ( .a ({new_AGEMA_signal_1135, n2732}), .b ({new_AGEMA_signal_5396, new_AGEMA_signal_5395}), .clk ( clk ), .r ({Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036]}), .c ({new_AGEMA_signal_1328, n1979}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2112 ( .a ({new_AGEMA_signal_5408, new_AGEMA_signal_5407}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040]}), .c ({new_AGEMA_signal_1152, n1985}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2121 ( .a ({new_AGEMA_signal_1154, n1992}), .b ({new_AGEMA_signal_1155, n1991}), .clk ( clk ), .r ({Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_1330, n1994}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2126 ( .a ({new_AGEMA_signal_5410, new_AGEMA_signal_5409}), .b ({new_AGEMA_signal_1156, n1995}), .clk ( clk ), .r ({Fresh[1051], Fresh[1050], Fresh[1049], Fresh[1048]}), .c ({new_AGEMA_signal_1331, n1996}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2136 ( .a ({new_AGEMA_signal_5412, new_AGEMA_signal_5411}), .b ({new_AGEMA_signal_1158, n2003}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052]}), .c ({new_AGEMA_signal_1332, n2137}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2142 ( .a ({new_AGEMA_signal_5414, new_AGEMA_signal_5413}), .b ({new_AGEMA_signal_1160, n2572}), .clk ( clk ), .r ({Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_1333, n2006}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2144 ( .a ({new_AGEMA_signal_5416, new_AGEMA_signal_5415}), .b ({new_AGEMA_signal_1161, n2004}), .clk ( clk ), .r ({Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060]}), .c ({new_AGEMA_signal_1334, n2005}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2152 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064]}), .c ({new_AGEMA_signal_1335, n2013}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2160 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419}), .b ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .r ({Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_1165, n2020}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2164 ( .a ({new_AGEMA_signal_1062, n2817}), .b ({new_AGEMA_signal_5422, new_AGEMA_signal_5421}), .clk ( clk ), .r ({Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072]}), .c ({new_AGEMA_signal_1166, n2023}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2168 ( .a ({new_AGEMA_signal_1009, n2027}), .b ({new_AGEMA_signal_5424, new_AGEMA_signal_5423}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076]}), .c ({new_AGEMA_signal_1071, n2028}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2172 ( .a ({new_AGEMA_signal_1167, n2214}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_1337, n2033}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2175 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_5428, new_AGEMA_signal_5427}), .clk ( clk ), .r ({Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084]}), .c ({new_AGEMA_signal_1338, n2031}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2184 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1170, n2039}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088]}), .c ({new_AGEMA_signal_1339, n2040}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2187 ( .a ({new_AGEMA_signal_5430, new_AGEMA_signal_5429}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ({Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_1171, n2050}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2193 ( .a ({new_AGEMA_signal_5432, new_AGEMA_signal_5431}), .b ({new_AGEMA_signal_1174, n2044}), .clk ( clk ), .r ({Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096]}), .c ({new_AGEMA_signal_1340, n2045}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2199 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_5396, new_AGEMA_signal_5395}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100]}), .c ({new_AGEMA_signal_1341, n2051}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2203 ( .a ({new_AGEMA_signal_5434, new_AGEMA_signal_5433}), .b ({new_AGEMA_signal_1176, n2055}), .clk ( clk ), .r ({Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_1342, n2056}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2209 ( .a ({new_AGEMA_signal_1178, n2407}), .b ({new_AGEMA_signal_5436, new_AGEMA_signal_5435}), .clk ( clk ), .r ({Fresh[1111], Fresh[1110], Fresh[1109], Fresh[1108]}), .c ({new_AGEMA_signal_1343, n2060}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2215 ( .a ({new_AGEMA_signal_5438, new_AGEMA_signal_5437}), .b ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112]}), .c ({new_AGEMA_signal_1344, n2066}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2217 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5423}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ({Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_1345, n2065}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2221 ( .a ({new_AGEMA_signal_1181, n2068}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ({Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120]}), .c ({new_AGEMA_signal_1346, n2069}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2226 ( .a ({new_AGEMA_signal_5440, new_AGEMA_signal_5439}), .b ({new_AGEMA_signal_1182, n2252}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124]}), .c ({new_AGEMA_signal_1347, n2074}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2235 ( .a ({new_AGEMA_signal_1076, n2081}), .b ({new_AGEMA_signal_1183, n2080}), .clk ( clk ), .r ({Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_1348, n2082}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2240 ( .a ({new_AGEMA_signal_5416, new_AGEMA_signal_5415}), .b ({new_AGEMA_signal_1185, n2083}), .clk ( clk ), .r ({Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132]}), .c ({new_AGEMA_signal_1349, n2084}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2242 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136]}), .c ({new_AGEMA_signal_1350, n2085}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2245 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441}), .b ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .r ({Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_1351, n2131}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2248 ( .a ({new_AGEMA_signal_1142, n2088}), .b ({new_AGEMA_signal_1078, n2087}), .clk ( clk ), .r ({Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144]}), .c ({new_AGEMA_signal_1352, n2089}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2252 ( .a ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .b ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148]}), .c ({new_AGEMA_signal_1353, n2330}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2254 ( .a ({new_AGEMA_signal_5444, new_AGEMA_signal_5443}), .b ({new_AGEMA_signal_1132, n2151}), .clk ( clk ), .r ({Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_1354, n2092}) ) ;
    or_GHPC #(.low_latency(1), .pipeline(1)) U2256 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1147, n2359}), .clk ( clk ), .r ({Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156]}), .c ({new_AGEMA_signal_1355, n2094}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2261 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1188, n2100}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160]}), .c ({new_AGEMA_signal_1356, n2160}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2265 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_1189, n2504}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2271 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ({Fresh[1171], Fresh[1170], Fresh[1169], Fresh[1168]}), .c ({new_AGEMA_signal_1504, n2114}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2273 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_5416, new_AGEMA_signal_5415}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172]}), .c ({new_AGEMA_signal_1190, n2115}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2280 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ({Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_1358, n2291}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2281 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ({Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180]}), .c ({new_AGEMA_signal_1192, n2119}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2291 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184]}), .c ({new_AGEMA_signal_1195, n2130}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2292 ( .a ({new_AGEMA_signal_1062, n2817}), .b ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .r ({Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_1196, n2129}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2295 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .clk ( clk ), .r ({Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192]}), .c ({new_AGEMA_signal_1197, n2150}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2298 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1082, n2132}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196]}), .c ({new_AGEMA_signal_1198, n2133}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2302 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_5452, new_AGEMA_signal_5451}), .clk ( clk ), .r ({Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_1361, n2136}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2306 ( .a ({new_AGEMA_signal_1160, n2572}), .b ({new_AGEMA_signal_1200, n2138}), .clk ( clk ), .r ({Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204]}), .c ({new_AGEMA_signal_1362, n2139}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2313 ( .a ({new_AGEMA_signal_5454, new_AGEMA_signal_5453}), .b ({new_AGEMA_signal_1201, n2555}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208]}), .c ({new_AGEMA_signal_1363, n2144}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2318 ( .a ({new_AGEMA_signal_1132, n2151}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ({Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_1364, n2152}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2321 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .r ({Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216]}), .c ({new_AGEMA_signal_1365, n2170}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2323 ( .a ({new_AGEMA_signal_1202, n2429}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220]}), .c ({new_AGEMA_signal_1366, n2157}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2329 ( .a ({new_AGEMA_signal_5456, new_AGEMA_signal_5455}), .b ({new_AGEMA_signal_1083, n2162}), .clk ( clk ), .r ({Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_1203, n2163}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2335 ( .a ({new_AGEMA_signal_1073, n2171}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ({Fresh[1231], Fresh[1230], Fresh[1229], Fresh[1228]}), .c ({new_AGEMA_signal_1368, n2172}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2338 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_1014, n2545}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232]}), .c ({new_AGEMA_signal_1084, n2186}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2339 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405}), .b ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .r ({Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_1369, n2181}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2344 ( .a ({new_AGEMA_signal_1204, n2176}), .b ({new_AGEMA_signal_1205, n2175}), .clk ( clk ), .r ({Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240]}), .c ({new_AGEMA_signal_1370, n2177}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2349 ( .a ({new_AGEMA_signal_5396, new_AGEMA_signal_5395}), .b ({new_AGEMA_signal_1016, n2182}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244]}), .c ({new_AGEMA_signal_1086, n2183}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2354 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457}), .b ({new_AGEMA_signal_1206, n2188}), .clk ( clk ), .r ({Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_1371, n2195}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2356 ( .a ({new_AGEMA_signal_1059, n2190}), .b ({new_AGEMA_signal_1207, n2189}), .clk ( clk ), .r ({Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252]}), .c ({new_AGEMA_signal_1372, n2193}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2358 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .b ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256]}), .c ({new_AGEMA_signal_1373, n2191}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2364 ( .a ({new_AGEMA_signal_1087, n2576}), .b ({new_AGEMA_signal_1088, n2748}), .clk ( clk ), .r ({Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_1209, n2196}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2367 ( .a ({new_AGEMA_signal_5390, new_AGEMA_signal_5389}), .b ({new_AGEMA_signal_1146, n2505}), .clk ( clk ), .r ({Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264]}), .c ({new_AGEMA_signal_1374, n2201}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2369 ( .a ({new_AGEMA_signal_1375, n2674}), .b ({new_AGEMA_signal_5462, new_AGEMA_signal_5461}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268]}), .c ({new_AGEMA_signal_1515, n2200}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2371 ( .s ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .b ({new_AGEMA_signal_1133, n2734}), .a ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ({Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_1516, n2202}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2379 ( .a ({new_AGEMA_signal_1167, n2214}), .b ({new_AGEMA_signal_1089, n2213}), .clk ( clk ), .r ({Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276]}), .c ({new_AGEMA_signal_1376, n2217}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2381 ( .a ({new_AGEMA_signal_5464, new_AGEMA_signal_5463}), .b ({new_AGEMA_signal_1090, n2215}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280]}), .c ({new_AGEMA_signal_1210, n2216}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2385 ( .a ({new_AGEMA_signal_1211, n2218}), .b ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .clk ( clk ), .r ({Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_1377, n2222}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2387 ( .a ({new_AGEMA_signal_1199, n2220}), .b ({new_AGEMA_signal_1212, n2219}), .clk ( clk ), .r ({Fresh[1291], Fresh[1290], Fresh[1289], Fresh[1288]}), .c ({new_AGEMA_signal_1378, n2221}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2391 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_5466, new_AGEMA_signal_5465}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292]}), .c ({new_AGEMA_signal_1213, n2226}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2393 ( .s ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .b ({new_AGEMA_signal_1056, n2651}), .a ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .r ({Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_1214, n2228}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2397 ( .a ({new_AGEMA_signal_5420, new_AGEMA_signal_5419}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ({Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300]}), .c ({new_AGEMA_signal_1215, n2237}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2398 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304]}), .c ({new_AGEMA_signal_1520, n2233}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2403 ( .a ({new_AGEMA_signal_5468, new_AGEMA_signal_5467}), .b ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .r ({Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_1216, n2238}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2406 ( .a ({new_AGEMA_signal_1157, n2241}), .b ({new_AGEMA_signal_1217, n2240}), .clk ( clk ), .r ({Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312]}), .c ({new_AGEMA_signal_1380, n2248}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2409 ( .a ({new_AGEMA_signal_1218, n2561}), .b ({new_AGEMA_signal_1219, n2243}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316]}), .c ({new_AGEMA_signal_1381, n2244}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2414 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_5380, new_AGEMA_signal_5379}), .clk ( clk ), .r ({Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_1382, n2249}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2417 ( .s ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .b ({new_AGEMA_signal_1182, n2252}), .a ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ({Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324]}), .c ({new_AGEMA_signal_1383, n2253}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2424 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_1222, n2259}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328]}), .c ({new_AGEMA_signal_1384, n2260}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2429 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_5470, new_AGEMA_signal_5469}), .clk ( clk ), .r ({Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_1524, n2273}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2430 ( .a ({new_AGEMA_signal_5472, new_AGEMA_signal_5471}), .b ({new_AGEMA_signal_1323, n2720}), .clk ( clk ), .r ({Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336]}), .c ({new_AGEMA_signal_1525, n2752}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2433 ( .a ({new_AGEMA_signal_1093, n2645}), .b ({new_AGEMA_signal_5446, new_AGEMA_signal_5445}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340]}), .c ({new_AGEMA_signal_1223, n2265}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2437 ( .a ({new_AGEMA_signal_5474, new_AGEMA_signal_5473}), .b ({new_AGEMA_signal_1094, n2268}), .clk ( clk ), .r ({Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_1224, n2269}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2444 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ({Fresh[1351], Fresh[1350], Fresh[1349], Fresh[1348]}), .c ({new_AGEMA_signal_1226, n2277}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2449 ( .a ({new_AGEMA_signal_5476, new_AGEMA_signal_5475}), .b ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352]}), .c ({new_AGEMA_signal_1227, n2282}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2452 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ({Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_1389, n2284}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2456 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_5478, new_AGEMA_signal_5477}), .clk ( clk ), .r ({Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360]}), .c ({new_AGEMA_signal_1390, n2459}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2459 ( .a ({new_AGEMA_signal_5384, new_AGEMA_signal_5383}), .b ({new_AGEMA_signal_1229, n2287}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364]}), .c ({new_AGEMA_signal_1391, n2288}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2462 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_1144, n2761}), .clk ( clk ), .r ({Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_1392, n2458}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2464 ( .a ({new_AGEMA_signal_5456, new_AGEMA_signal_5455}), .b ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .r ({Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372]}), .c ({new_AGEMA_signal_1393, n2293}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2467 ( .a ({new_AGEMA_signal_5444, new_AGEMA_signal_5443}), .b ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376]}), .c ({new_AGEMA_signal_1230, n2294}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2472 ( .a ({new_AGEMA_signal_1231, n2438}), .b ({new_AGEMA_signal_1096, n2299}), .clk ( clk ), .r ({Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_1394, n2300}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2480 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .clk ( clk ), .r ({Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384]}), .c ({new_AGEMA_signal_1395, n2323}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) U2482 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1232, n2371}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388]}), .c ({new_AGEMA_signal_1396, n2314}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2485 ( .a ({new_AGEMA_signal_1018, n2316}), .b ({new_AGEMA_signal_5480, new_AGEMA_signal_5479}), .clk ( clk ), .r ({Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_1097, n2319}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2491 ( .a ({new_AGEMA_signal_1074, n2642}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ({Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396]}), .c ({new_AGEMA_signal_1234, n2326}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2496 ( .a ({new_AGEMA_signal_1236, n2328}), .b ({new_AGEMA_signal_1099, n2327}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400]}), .c ({new_AGEMA_signal_1398, n2329}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2501 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ({Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_1537, n2335}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2506 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ({Fresh[1411], Fresh[1410], Fresh[1409], Fresh[1408]}), .c ({new_AGEMA_signal_1399, n2341}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2507 ( .a ({new_AGEMA_signal_5482, new_AGEMA_signal_5481}), .b ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412]}), .c ({new_AGEMA_signal_1238, n2340}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2514 ( .a ({new_AGEMA_signal_1100, n2348}), .b ({new_AGEMA_signal_1101, n2347}), .clk ( clk ), .r ({Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_1240, n2349}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2517 ( .a ({new_AGEMA_signal_5484, new_AGEMA_signal_5483}), .b ({new_AGEMA_signal_1061, n2690}), .clk ( clk ), .r ({Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420]}), .c ({new_AGEMA_signal_1241, n2375}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2518 ( .a ({new_AGEMA_signal_5454, new_AGEMA_signal_5453}), .b ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424]}), .c ({new_AGEMA_signal_1242, n2352}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2522 ( .a ({new_AGEMA_signal_1243, n2353}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ({Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_1401, n2354}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2525 ( .a ({new_AGEMA_signal_5486, new_AGEMA_signal_5485}), .b ({new_AGEMA_signal_1244, n2355}), .clk ( clk ), .r ({Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432]}), .c ({new_AGEMA_signal_1402, n2357}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2527 ( .a ({new_AGEMA_signal_1147, n2359}), .b ({new_AGEMA_signal_5488, new_AGEMA_signal_5487}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436]}), .c ({new_AGEMA_signal_1403, n2360}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2534 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ({Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_1540, n2369}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2536 ( .a ({new_AGEMA_signal_1232, n2371}), .b ({new_AGEMA_signal_5466, new_AGEMA_signal_5465}), .clk ( clk ), .r ({Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444]}), .c ({new_AGEMA_signal_1404, n2372}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2539 ( .a ({new_AGEMA_signal_1087, n2576}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448]}), .c ({new_AGEMA_signal_1405, n2377}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2544 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .b ({new_AGEMA_signal_1103, n2415}), .clk ( clk ), .r ({Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_1246, n2467}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2545 ( .a ({new_AGEMA_signal_5490, new_AGEMA_signal_5489}), .b ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .r ({Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456]}), .c ({new_AGEMA_signal_1247, n2385}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2546 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460]}), .c ({new_AGEMA_signal_1248, n2384}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2548 ( .a ({new_AGEMA_signal_5416, new_AGEMA_signal_5415}), .b ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .r ({Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_1407, n2386}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2552 ( .a ({new_AGEMA_signal_5458, new_AGEMA_signal_5457}), .b ({new_AGEMA_signal_1081, n2647}), .clk ( clk ), .r ({Fresh[1471], Fresh[1470], Fresh[1469], Fresh[1468]}), .c ({new_AGEMA_signal_1249, n2394}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2553 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472]}), .c ({new_AGEMA_signal_1250, n2391}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2554 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_1408, n2390}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2559 ( .a ({new_AGEMA_signal_5444, new_AGEMA_signal_5443}), .b ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .r ({Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480]}), .c ({new_AGEMA_signal_1251, n2396}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2562 ( .a ({new_AGEMA_signal_5492, new_AGEMA_signal_5491}), .b ({new_AGEMA_signal_1231, n2438}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484]}), .c ({new_AGEMA_signal_1409, n2406}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2565 ( .a ({new_AGEMA_signal_1105, n2594}), .b ({new_AGEMA_signal_1106, n2402}), .clk ( clk ), .r ({Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_1252, n2403}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2569 ( .a ({new_AGEMA_signal_1178, n2407}), .b ({new_AGEMA_signal_5452, new_AGEMA_signal_5451}), .clk ( clk ), .r ({Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492]}), .c ({new_AGEMA_signal_1411, n2408}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2573 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5467}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496]}), .c ({new_AGEMA_signal_1412, n2574}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2574 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_5432, new_AGEMA_signal_5431}), .clk ( clk ), .r ({Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_1253, n2413}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2577 ( .a ({new_AGEMA_signal_1103, n2415}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504]}), .c ({new_AGEMA_signal_1254, n2416}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2586 ( .a ({new_AGEMA_signal_1255, n2428}), .b ({new_AGEMA_signal_5494, new_AGEMA_signal_5493}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508]}), .c ({new_AGEMA_signal_1414, n2433}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2587 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .b ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .r ({Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_1415, n2689}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2591 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .r ({Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516]}), .c ({new_AGEMA_signal_1257, n2434}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2595 ( .a ({new_AGEMA_signal_1231, n2438}), .b ({new_AGEMA_signal_1107, n2483}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520]}), .c ({new_AGEMA_signal_1417, n2439}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2598 ( .a ({new_AGEMA_signal_5490, new_AGEMA_signal_5489}), .b ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .r ({Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_1418, n2445}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2600 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1258, n2443}), .clk ( clk ), .r ({Fresh[1531], Fresh[1530], Fresh[1529], Fresh[1528]}), .c ({new_AGEMA_signal_1419, n2444}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2602 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405}), .b ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532]}), .c ({new_AGEMA_signal_1420, n2447}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2607 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .r ({Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_1421, n2454}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2617 ( .a ({new_AGEMA_signal_5446, new_AGEMA_signal_5445}), .b ({new_AGEMA_signal_1109, n2464}), .clk ( clk ), .r ({Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540]}), .c ({new_AGEMA_signal_1260, n2465}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2622 ( .a ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .b ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544]}), .c ({new_AGEMA_signal_1261, n2470}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2626 ( .a ({new_AGEMA_signal_1111, n2473}), .b ({new_AGEMA_signal_1112, n2472}), .clk ( clk ), .r ({Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_1262, n2476}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2633 ( .a ({new_AGEMA_signal_5496, new_AGEMA_signal_5495}), .b ({new_AGEMA_signal_1263, n2480}), .clk ( clk ), .r ({Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552]}), .c ({new_AGEMA_signal_1424, n2481}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2639 ( .a ({new_AGEMA_signal_5498, new_AGEMA_signal_5497}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556]}), .c ({new_AGEMA_signal_1265, n2486}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2642 ( .a ({new_AGEMA_signal_5472, new_AGEMA_signal_5471}), .b ({new_AGEMA_signal_1114, n2488}), .clk ( clk ), .r ({Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_1266, n2489}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2645 ( .a ({new_AGEMA_signal_5500, new_AGEMA_signal_5499}), .b ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .r ({Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564]}), .c ({new_AGEMA_signal_1267, n2497}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2646 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501}), .b ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568]}), .c ({new_AGEMA_signal_1268, n2495}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2647 ( .a ({new_AGEMA_signal_5448, new_AGEMA_signal_5447}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ({Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_1426, n2494}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2650 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_5390, new_AGEMA_signal_5389}), .clk ( clk ), .r ({Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576]}), .c ({new_AGEMA_signal_1269, n2499}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2653 ( .a ({new_AGEMA_signal_5390, new_AGEMA_signal_5389}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580]}), .c ({new_AGEMA_signal_1557, n2503}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2655 ( .s ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .b ({new_AGEMA_signal_1146, n2505}), .a ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ({Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_1427, n2506}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2662 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_5412, new_AGEMA_signal_5411}), .clk ( clk ), .r ({Fresh[1591], Fresh[1590], Fresh[1589], Fresh[1588]}), .c ({new_AGEMA_signal_1428, n2518}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2663 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592]}), .c ({new_AGEMA_signal_1558, n2517}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2666 ( .a ({new_AGEMA_signal_1270, n2520}), .b ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .clk ( clk ), .r ({Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_1429, n2523}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2668 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_1115, n2521}), .clk ( clk ), .r ({Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600]}), .c ({new_AGEMA_signal_1430, n2522}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2675 ( .a ({new_AGEMA_signal_5412, new_AGEMA_signal_5411}), .b ({new_AGEMA_signal_1271, n2531}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604]}), .c ({new_AGEMA_signal_1431, n2532}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2677 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ({Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_1432, n2534}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2681 ( .a ({new_AGEMA_signal_5504, new_AGEMA_signal_5503}), .b ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .r ({Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612]}), .c ({new_AGEMA_signal_1433, n2542}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2683 ( .a ({new_AGEMA_signal_1014, n2545}), .b ({new_AGEMA_signal_1079, n2544}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616]}), .c ({new_AGEMA_signal_1272, n2546}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2687 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ({Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_1435, n2551}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2690 ( .a ({new_AGEMA_signal_1273, n2553}), .b ({new_AGEMA_signal_5506, new_AGEMA_signal_5505}), .clk ( clk ), .r ({Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624]}), .c ({new_AGEMA_signal_1436, n2558}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2692 ( .a ({new_AGEMA_signal_1201, n2555}), .b ({new_AGEMA_signal_1274, n2554}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628]}), .c ({new_AGEMA_signal_1437, n2556}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2696 ( .a ({new_AGEMA_signal_1218, n2561}), .b ({new_AGEMA_signal_1116, n2560}), .clk ( clk ), .r ({Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_1438, n2566}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2697 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507}), .b ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .r ({Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636]}), .c ({new_AGEMA_signal_1439, n2715}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2703 ( .a ({new_AGEMA_signal_1160, n2572}), .b ({new_AGEMA_signal_1055, n2571}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640]}), .c ({new_AGEMA_signal_1440, n2573}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2705 ( .a ({new_AGEMA_signal_5492, new_AGEMA_signal_5491}), .b ({new_AGEMA_signal_1173, n2754}), .clk ( clk ), .r ({Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_1441, n2585}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2706 ( .a ({new_AGEMA_signal_5470, new_AGEMA_signal_5469}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ({Fresh[1651], Fresh[1650], Fresh[1649], Fresh[1648]}), .c ({new_AGEMA_signal_1276, n2581}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2707 ( .a ({new_AGEMA_signal_1127, n2575}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652]}), .c ({new_AGEMA_signal_1442, n2579}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2708 ( .a ({new_AGEMA_signal_5502, new_AGEMA_signal_5501}), .b ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .r ({Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_1277, n2578}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2711 ( .a ({new_AGEMA_signal_1148, n2625}), .b ({new_AGEMA_signal_5462, new_AGEMA_signal_5461}), .clk ( clk ), .r ({Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660]}), .c ({new_AGEMA_signal_1443, n2582}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2715 ( .a ({new_AGEMA_signal_5398, new_AGEMA_signal_5397}), .b ({new_AGEMA_signal_1278, n2586}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664]}), .c ({new_AGEMA_signal_1444, n2588}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2719 ( .a ({new_AGEMA_signal_1105, n2594}), .b ({new_AGEMA_signal_5492, new_AGEMA_signal_5491}), .clk ( clk ), .r ({Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_1279, n2607}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2722 ( .a ({new_AGEMA_signal_1117, n2597}), .b ({new_AGEMA_signal_1280, n2596}), .clk ( clk ), .r ({Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672]}), .c ({new_AGEMA_signal_1445, n2605}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2724 ( .a ({new_AGEMA_signal_1281, n2598}), .b ({new_AGEMA_signal_5510, new_AGEMA_signal_5509}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676]}), .c ({new_AGEMA_signal_1446, n2603}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2726 ( .a ({new_AGEMA_signal_1021, n2599}), .b ({new_AGEMA_signal_5468, new_AGEMA_signal_5467}), .clk ( clk ), .r ({Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_1118, n2601}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2733 ( .a ({new_AGEMA_signal_1283, n2610}), .b ({new_AGEMA_signal_5460, new_AGEMA_signal_5459}), .clk ( clk ), .r ({Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684]}), .c ({new_AGEMA_signal_1447, n2620}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2736 ( .a ({new_AGEMA_signal_1284, n2614}), .b ({new_AGEMA_signal_1285, n2613}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688]}), .c ({new_AGEMA_signal_1448, n2618}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2743 ( .a ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ({Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_1449, n2626}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2746 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_5426, new_AGEMA_signal_5425}), .clk ( clk ), .r ({Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696]}), .c ({new_AGEMA_signal_1286, n2632}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2752 ( .a ({new_AGEMA_signal_1287, n2784}), .b ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700]}), .c ({new_AGEMA_signal_1450, n2644}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2754 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387}), .b ({new_AGEMA_signal_1093, n2645}), .clk ( clk ), .r ({Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_1288, n2646}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2758 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_1121, n2650}), .clk ( clk ), .r ({Fresh[1711], Fresh[1710], Fresh[1709], Fresh[1708]}), .c ({new_AGEMA_signal_1289, n2653}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2760 ( .a ({new_AGEMA_signal_5468, new_AGEMA_signal_5467}), .b ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712]}), .c ({new_AGEMA_signal_1452, n2655}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2764 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471}), .clk ( clk ), .r ({Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_1453, n2663}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2770 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_5462, new_AGEMA_signal_5461}), .clk ( clk ), .r ({Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720]}), .c ({new_AGEMA_signal_1290, n2675}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2772 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1043, n2676}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724]}), .c ({new_AGEMA_signal_1291, n2678}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2780 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_5470, new_AGEMA_signal_5469}), .clk ( clk ), .r ({Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_1292, n2691}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2782 ( .a ({new_AGEMA_signal_5476, new_AGEMA_signal_5475}), .b ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .r ({Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732]}), .c ({new_AGEMA_signal_1455, n2695}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2785 ( .a ({new_AGEMA_signal_1104, n2700}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736]}), .c ({new_AGEMA_signal_1293, n2701}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2791 ( .a ({new_AGEMA_signal_1294, n2711}), .b ({new_AGEMA_signal_1295, n2710}), .clk ( clk ), .r ({Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_1456, n2717}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2796 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_5450, new_AGEMA_signal_5449}), .clk ( clk ), .r ({Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744]}), .c ({new_AGEMA_signal_1576, n2729}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2798 ( .a ({new_AGEMA_signal_5416, new_AGEMA_signal_5415}), .b ({new_AGEMA_signal_1123, n2722}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748]}), .c ({new_AGEMA_signal_1296, n2727}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2803 ( .a ({new_AGEMA_signal_1135, n2732}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ({Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_1458, n2733}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2807 ( .a ({new_AGEMA_signal_5512, new_AGEMA_signal_5511}), .b ({new_AGEMA_signal_1298, n2738}), .clk ( clk ), .r ({Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756]}), .c ({new_AGEMA_signal_1459, n2740}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2812 ( .a ({new_AGEMA_signal_1088, n2748}), .b ({new_AGEMA_signal_5380, new_AGEMA_signal_5379}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760]}), .c ({new_AGEMA_signal_1299, n2749}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2815 ( .a ({new_AGEMA_signal_1173, n2754}), .b ({new_AGEMA_signal_5420, new_AGEMA_signal_5419}), .clk ( clk ), .r ({Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_1461, n2757}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2816 ( .a ({new_AGEMA_signal_1030, n2755}), .b ({new_AGEMA_signal_5514, new_AGEMA_signal_5513}), .clk ( clk ), .r ({Fresh[1771], Fresh[1770], Fresh[1769], Fresh[1768]}), .c ({new_AGEMA_signal_1300, n2756}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2819 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_5478, new_AGEMA_signal_5477}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772]}), .c ({new_AGEMA_signal_1462, n2762}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2823 ( .a ({new_AGEMA_signal_5380, new_AGEMA_signal_5379}), .b ({new_AGEMA_signal_1301, n2768}), .clk ( clk ), .r ({Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_1463, n2770}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2825 ( .a ({new_AGEMA_signal_1184, n2773}), .b ({new_AGEMA_signal_5514, new_AGEMA_signal_5513}), .clk ( clk ), .r ({Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780]}), .c ({new_AGEMA_signal_1464, n2776}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2826 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_5382, new_AGEMA_signal_5381}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784]}), .c ({new_AGEMA_signal_1465, n2775}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2830 ( .a ({new_AGEMA_signal_1124, n2782}), .b ({new_AGEMA_signal_1125, n2781}), .clk ( clk ), .r ({Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_1302, n2783}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2836 ( .a ({new_AGEMA_signal_1304, n2794}), .b ({new_AGEMA_signal_1305, n2793}), .clk ( clk ), .r ({Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792]}), .c ({new_AGEMA_signal_1467, n2795}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2845 ( .a ({new_AGEMA_signal_1306, n2812}), .b ({new_AGEMA_signal_1194, n2811}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796]}), .c ({new_AGEMA_signal_1468, n2814}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2848 ( .a ({new_AGEMA_signal_5404, new_AGEMA_signal_5403}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ({Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_1307, n2819}) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C ( clk ), .D ( n2755 ), .Q ( new_AGEMA_signal_5515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_5516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C ( clk ), .D ( n2151 ), .Q ( new_AGEMA_signal_5517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C ( clk ), .D ( new_AGEMA_signal_1132 ), .Q ( new_AGEMA_signal_5518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C ( clk ), .D ( new_AGEMA_signal_5519 ), .Q ( new_AGEMA_signal_5520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C ( clk ), .D ( new_AGEMA_signal_5521 ), .Q ( new_AGEMA_signal_5522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C ( clk ), .D ( new_AGEMA_signal_5395 ), .Q ( new_AGEMA_signal_5523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C ( clk ), .D ( new_AGEMA_signal_5396 ), .Q ( new_AGEMA_signal_5524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C ( clk ), .D ( new_AGEMA_signal_5389 ), .Q ( new_AGEMA_signal_5525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C ( clk ), .D ( new_AGEMA_signal_5390 ), .Q ( new_AGEMA_signal_5526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C ( clk ), .D ( n1964 ), .Q ( new_AGEMA_signal_5527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C ( clk ), .D ( new_AGEMA_signal_999 ), .Q ( new_AGEMA_signal_5528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C ( clk ), .D ( n2673 ), .Q ( new_AGEMA_signal_5529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C ( clk ), .D ( new_AGEMA_signal_1052 ), .Q ( new_AGEMA_signal_5530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C ( clk ), .D ( n2359 ), .Q ( new_AGEMA_signal_5531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C ( clk ), .D ( new_AGEMA_signal_1147 ), .Q ( new_AGEMA_signal_5532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C ( clk ), .D ( n1973 ), .Q ( new_AGEMA_signal_5533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C ( clk ), .D ( new_AGEMA_signal_1151 ), .Q ( new_AGEMA_signal_5534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C ( clk ), .D ( n2690 ), .Q ( new_AGEMA_signal_5535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_5536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C ( clk ), .D ( n2741 ), .Q ( new_AGEMA_signal_5537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C ( clk ), .D ( new_AGEMA_signal_1153 ), .Q ( new_AGEMA_signal_5538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C ( clk ), .D ( n1993 ), .Q ( new_AGEMA_signal_5539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_5540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C ( clk ), .D ( n2241 ), .Q ( new_AGEMA_signal_5541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C ( clk ), .D ( new_AGEMA_signal_1157 ), .Q ( new_AGEMA_signal_5542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C ( clk ), .D ( new_AGEMA_signal_5449 ), .Q ( new_AGEMA_signal_5543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C ( clk ), .D ( new_AGEMA_signal_5450 ), .Q ( new_AGEMA_signal_5544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C ( clk ), .D ( new_AGEMA_signal_5545 ), .Q ( new_AGEMA_signal_5546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C ( clk ), .D ( new_AGEMA_signal_5547 ), .Q ( new_AGEMA_signal_5548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C ( clk ), .D ( n2290 ), .Q ( new_AGEMA_signal_5549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C ( clk ), .D ( new_AGEMA_signal_1168 ), .Q ( new_AGEMA_signal_5550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C ( clk ), .D ( n2171 ), .Q ( new_AGEMA_signal_5551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_5552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C ( clk ), .D ( n2042 ), .Q ( new_AGEMA_signal_5553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C ( clk ), .D ( new_AGEMA_signal_1172 ), .Q ( new_AGEMA_signal_5554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C ( clk ), .D ( n2754 ), .Q ( new_AGEMA_signal_5555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C ( clk ), .D ( new_AGEMA_signal_1173 ), .Q ( new_AGEMA_signal_5556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C ( clk ), .D ( new_AGEMA_signal_5379 ), .Q ( new_AGEMA_signal_5557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C ( clk ), .D ( new_AGEMA_signal_5380 ), .Q ( new_AGEMA_signal_5558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C ( clk ), .D ( n2535 ), .Q ( new_AGEMA_signal_5559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C ( clk ), .D ( new_AGEMA_signal_1150 ), .Q ( new_AGEMA_signal_5560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C ( clk ), .D ( n2642 ), .Q ( new_AGEMA_signal_5561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_5562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C ( clk ), .D ( new_AGEMA_signal_5563 ), .Q ( new_AGEMA_signal_5564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C ( clk ), .D ( new_AGEMA_signal_5565 ), .Q ( new_AGEMA_signal_5566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C ( clk ), .D ( n2773 ), .Q ( new_AGEMA_signal_5567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C ( clk ), .D ( new_AGEMA_signal_1184 ), .Q ( new_AGEMA_signal_5568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C ( clk ), .D ( n2627 ), .Q ( new_AGEMA_signal_5569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C ( clk ), .D ( new_AGEMA_signal_1048 ), .Q ( new_AGEMA_signal_5570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C ( clk ), .D ( new_AGEMA_signal_5419 ), .Q ( new_AGEMA_signal_5571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C ( clk ), .D ( new_AGEMA_signal_5420 ), .Q ( new_AGEMA_signal_5572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C ( clk ), .D ( n2631 ), .Q ( new_AGEMA_signal_5573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C ( clk ), .D ( new_AGEMA_signal_1034 ), .Q ( new_AGEMA_signal_5574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C ( clk ), .D ( n2376 ), .Q ( new_AGEMA_signal_5575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C ( clk ), .D ( new_AGEMA_signal_1169 ), .Q ( new_AGEMA_signal_5576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C ( clk ), .D ( new_AGEMA_signal_5577 ), .Q ( new_AGEMA_signal_5578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C ( clk ), .D ( new_AGEMA_signal_5579 ), .Q ( new_AGEMA_signal_5580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C ( clk ), .D ( new_AGEMA_signal_5465 ), .Q ( new_AGEMA_signal_5581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C ( clk ), .D ( new_AGEMA_signal_5466 ), .Q ( new_AGEMA_signal_5582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C ( clk ), .D ( new_AGEMA_signal_5429 ), .Q ( new_AGEMA_signal_5583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C ( clk ), .D ( new_AGEMA_signal_5430 ), .Q ( new_AGEMA_signal_5584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C ( clk ), .D ( new_AGEMA_signal_5437 ), .Q ( new_AGEMA_signal_5585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C ( clk ), .D ( new_AGEMA_signal_5438 ), .Q ( new_AGEMA_signal_5586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C ( clk ), .D ( new_AGEMA_signal_5587 ), .Q ( new_AGEMA_signal_5588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C ( clk ), .D ( new_AGEMA_signal_5589 ), .Q ( new_AGEMA_signal_5590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C ( clk ), .D ( new_AGEMA_signal_5505 ), .Q ( new_AGEMA_signal_5591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C ( clk ), .D ( new_AGEMA_signal_5506 ), .Q ( new_AGEMA_signal_5592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C ( clk ), .D ( n2498 ), .Q ( new_AGEMA_signal_5593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C ( clk ), .D ( new_AGEMA_signal_1077 ), .Q ( new_AGEMA_signal_5594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C ( clk ), .D ( n2178 ), .Q ( new_AGEMA_signal_5595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_5596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C ( clk ), .D ( new_AGEMA_signal_5597 ), .Q ( new_AGEMA_signal_5598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C ( clk ), .D ( new_AGEMA_signal_5599 ), .Q ( new_AGEMA_signal_5600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C ( clk ), .D ( n2505 ), .Q ( new_AGEMA_signal_5601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C ( clk ), .D ( new_AGEMA_signal_1146 ), .Q ( new_AGEMA_signal_5602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C ( clk ), .D ( n2540 ), .Q ( new_AGEMA_signal_5603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C ( clk ), .D ( new_AGEMA_signal_1221 ), .Q ( new_AGEMA_signal_5604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C ( clk ), .D ( n2266 ), .Q ( new_AGEMA_signal_5605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_5606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C ( clk ), .D ( n2278 ), .Q ( new_AGEMA_signal_5607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C ( clk ), .D ( new_AGEMA_signal_1225 ), .Q ( new_AGEMA_signal_5608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C ( clk ), .D ( new_AGEMA_signal_5461 ), .Q ( new_AGEMA_signal_5609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C ( clk ), .D ( new_AGEMA_signal_5462 ), .Q ( new_AGEMA_signal_5610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C ( clk ), .D ( new_AGEMA_signal_5483 ), .Q ( new_AGEMA_signal_5611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C ( clk ), .D ( new_AGEMA_signal_5484 ), .Q ( new_AGEMA_signal_5612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C ( clk ), .D ( new_AGEMA_signal_5415 ), .Q ( new_AGEMA_signal_5613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C ( clk ), .D ( new_AGEMA_signal_5416 ), .Q ( new_AGEMA_signal_5614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C ( clk ), .D ( new_AGEMA_signal_5411 ), .Q ( new_AGEMA_signal_5615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C ( clk ), .D ( new_AGEMA_signal_5412 ), .Q ( new_AGEMA_signal_5616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C ( clk ), .D ( n2318 ), .Q ( new_AGEMA_signal_5617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C ( clk ), .D ( new_AGEMA_signal_1098 ), .Q ( new_AGEMA_signal_5618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C ( clk ), .D ( n2325 ), .Q ( new_AGEMA_signal_5619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C ( clk ), .D ( new_AGEMA_signal_1235 ), .Q ( new_AGEMA_signal_5620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C ( clk ), .D ( n2677 ), .Q ( new_AGEMA_signal_5621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C ( clk ), .D ( new_AGEMA_signal_1047 ), .Q ( new_AGEMA_signal_5622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C ( clk ), .D ( new_AGEMA_signal_5501 ), .Q ( new_AGEMA_signal_5623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C ( clk ), .D ( new_AGEMA_signal_5502 ), .Q ( new_AGEMA_signal_5624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C ( clk ), .D ( new_AGEMA_signal_5509 ), .Q ( new_AGEMA_signal_5625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C ( clk ), .D ( new_AGEMA_signal_5510 ), .Q ( new_AGEMA_signal_5626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C ( clk ), .D ( new_AGEMA_signal_5433 ), .Q ( new_AGEMA_signal_5627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C ( clk ), .D ( new_AGEMA_signal_5434 ), .Q ( new_AGEMA_signal_5628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C ( clk ), .D ( new_AGEMA_signal_5383 ), .Q ( new_AGEMA_signal_5629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C ( clk ), .D ( new_AGEMA_signal_5384 ), .Q ( new_AGEMA_signal_5630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C ( clk ), .D ( n2625 ), .Q ( new_AGEMA_signal_5631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C ( clk ), .D ( new_AGEMA_signal_1148 ), .Q ( new_AGEMA_signal_5632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C ( clk ), .D ( n2431 ), .Q ( new_AGEMA_signal_5633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C ( clk ), .D ( new_AGEMA_signal_1256 ), .Q ( new_AGEMA_signal_5634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C ( clk ), .D ( new_AGEMA_signal_5636 ), .Q ( new_AGEMA_signal_5637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C ( clk ), .D ( new_AGEMA_signal_5639 ), .Q ( new_AGEMA_signal_5640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C ( clk ), .D ( n2453 ), .Q ( new_AGEMA_signal_5641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_5642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C ( clk ), .D ( n2475 ), .Q ( new_AGEMA_signal_5643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C ( clk ), .D ( new_AGEMA_signal_1113 ), .Q ( new_AGEMA_signal_5644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C ( clk ), .D ( n2487 ), .Q ( new_AGEMA_signal_5645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C ( clk ), .D ( new_AGEMA_signal_1264 ), .Q ( new_AGEMA_signal_5646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C ( clk ), .D ( new_AGEMA_signal_5647 ), .Q ( new_AGEMA_signal_5648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C ( clk ), .D ( new_AGEMA_signal_5649 ), .Q ( new_AGEMA_signal_5650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C ( clk ), .D ( new_AGEMA_signal_5453 ), .Q ( new_AGEMA_signal_5651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C ( clk ), .D ( new_AGEMA_signal_5454 ), .Q ( new_AGEMA_signal_5652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C ( clk ), .D ( new_AGEMA_signal_5457 ), .Q ( new_AGEMA_signal_5653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C ( clk ), .D ( new_AGEMA_signal_5458 ), .Q ( new_AGEMA_signal_5654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C ( clk ), .D ( n2564 ), .Q ( new_AGEMA_signal_5655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C ( clk ), .D ( new_AGEMA_signal_1275 ), .Q ( new_AGEMA_signal_5656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C ( clk ), .D ( new_AGEMA_signal_5657 ), .Q ( new_AGEMA_signal_5658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C ( clk ), .D ( new_AGEMA_signal_5659 ), .Q ( new_AGEMA_signal_5660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C ( clk ), .D ( n2617 ), .Q ( new_AGEMA_signal_5661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C ( clk ), .D ( new_AGEMA_signal_1119 ), .Q ( new_AGEMA_signal_5662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C ( clk ), .D ( n2647 ), .Q ( new_AGEMA_signal_5663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_5664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C ( clk ), .D ( n2674 ), .Q ( new_AGEMA_signal_5665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C ( clk ), .D ( new_AGEMA_signal_1375 ), .Q ( new_AGEMA_signal_5666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C ( clk ), .D ( n2683 ), .Q ( new_AGEMA_signal_5667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C ( clk ), .D ( new_AGEMA_signal_1022 ), .Q ( new_AGEMA_signal_5668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C ( clk ), .D ( n2714 ), .Q ( new_AGEMA_signal_5669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C ( clk ), .D ( new_AGEMA_signal_1122 ), .Q ( new_AGEMA_signal_5670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C ( clk ), .D ( n2726 ), .Q ( new_AGEMA_signal_5671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C ( clk ), .D ( new_AGEMA_signal_1297 ), .Q ( new_AGEMA_signal_5672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C ( clk ), .D ( n2734 ), .Q ( new_AGEMA_signal_5673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C ( clk ), .D ( new_AGEMA_signal_1133 ), .Q ( new_AGEMA_signal_5674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C ( clk ), .D ( new_AGEMA_signal_5675 ), .Q ( new_AGEMA_signal_5676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C ( clk ), .D ( new_AGEMA_signal_5677 ), .Q ( new_AGEMA_signal_5678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C ( clk ), .D ( n2763 ), .Q ( new_AGEMA_signal_5679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C ( clk ), .D ( new_AGEMA_signal_1134 ), .Q ( new_AGEMA_signal_5680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C ( clk ), .D ( n2784 ), .Q ( new_AGEMA_signal_5681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C ( clk ), .D ( new_AGEMA_signal_1287 ), .Q ( new_AGEMA_signal_5682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C ( clk ), .D ( new_AGEMA_signal_5683 ), .Q ( new_AGEMA_signal_5684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C ( clk ), .D ( new_AGEMA_signal_5685 ), .Q ( new_AGEMA_signal_5686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C ( clk ), .D ( n2820 ), .Q ( new_AGEMA_signal_5687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C ( clk ), .D ( new_AGEMA_signal_1126 ), .Q ( new_AGEMA_signal_5688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C ( clk ), .D ( new_AGEMA_signal_5497 ), .Q ( new_AGEMA_signal_5689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C ( clk ), .D ( new_AGEMA_signal_5498 ), .Q ( new_AGEMA_signal_5691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C ( clk ), .D ( n1930 ), .Q ( new_AGEMA_signal_5693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C ( clk ), .D ( new_AGEMA_signal_1036 ), .Q ( new_AGEMA_signal_5695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C ( clk ), .D ( n1976 ), .Q ( new_AGEMA_signal_5701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_5703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C ( clk ), .D ( new_AGEMA_signal_5413 ), .Q ( new_AGEMA_signal_5707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C ( clk ), .D ( new_AGEMA_signal_5414 ), .Q ( new_AGEMA_signal_5709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C ( clk ), .D ( n2008 ), .Q ( new_AGEMA_signal_5713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C ( clk ), .D ( new_AGEMA_signal_1159 ), .Q ( new_AGEMA_signal_5715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C ( clk ), .D ( n2022 ), .Q ( new_AGEMA_signal_5717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C ( clk ), .D ( new_AGEMA_signal_1164 ), .Q ( new_AGEMA_signal_5719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C ( clk ), .D ( n2057 ), .Q ( new_AGEMA_signal_5729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C ( clk ), .D ( new_AGEMA_signal_1177 ), .Q ( new_AGEMA_signal_5731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C ( clk ), .D ( n2062 ), .Q ( new_AGEMA_signal_5733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C ( clk ), .D ( new_AGEMA_signal_1179 ), .Q ( new_AGEMA_signal_5735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C ( clk ), .D ( n2075 ), .Q ( new_AGEMA_signal_5737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_5739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C ( clk ), .D ( n2121 ), .Q ( new_AGEMA_signal_5747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C ( clk ), .D ( new_AGEMA_signal_1191 ), .Q ( new_AGEMA_signal_5749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C ( clk ), .D ( new_AGEMA_signal_5403 ), .Q ( new_AGEMA_signal_5753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C ( clk ), .D ( new_AGEMA_signal_5404 ), .Q ( new_AGEMA_signal_5755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C ( clk ), .D ( new_AGEMA_signal_5757 ), .Q ( new_AGEMA_signal_5758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C ( clk ), .D ( new_AGEMA_signal_5760 ), .Q ( new_AGEMA_signal_5761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C ( clk ), .D ( new_AGEMA_signal_5475 ), .Q ( new_AGEMA_signal_5763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C ( clk ), .D ( new_AGEMA_signal_5476 ), .Q ( new_AGEMA_signal_5765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C ( clk ), .D ( new_AGEMA_signal_5489 ), .Q ( new_AGEMA_signal_5767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C ( clk ), .D ( new_AGEMA_signal_5490 ), .Q ( new_AGEMA_signal_5769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C ( clk ), .D ( n2245 ), .Q ( new_AGEMA_signal_5779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C ( clk ), .D ( new_AGEMA_signal_1220 ), .Q ( new_AGEMA_signal_5781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C ( clk ), .D ( new_AGEMA_signal_5783 ), .Q ( new_AGEMA_signal_5784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C ( clk ), .D ( new_AGEMA_signal_5786 ), .Q ( new_AGEMA_signal_5787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C ( clk ), .D ( n2262 ), .Q ( new_AGEMA_signal_5789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C ( clk ), .D ( new_AGEMA_signal_1091 ), .Q ( new_AGEMA_signal_5791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C ( clk ), .D ( n2343 ), .Q ( new_AGEMA_signal_5799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C ( clk ), .D ( new_AGEMA_signal_1237 ), .Q ( new_AGEMA_signal_5801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C ( clk ), .D ( new_AGEMA_signal_5477 ), .Q ( new_AGEMA_signal_5807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C ( clk ), .D ( new_AGEMA_signal_5478 ), .Q ( new_AGEMA_signal_5809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C ( clk ), .D ( new_AGEMA_signal_5469 ), .Q ( new_AGEMA_signal_5811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C ( clk ), .D ( new_AGEMA_signal_5470 ), .Q ( new_AGEMA_signal_5813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C ( clk ), .D ( new_AGEMA_signal_5399 ), .Q ( new_AGEMA_signal_5815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C ( clk ), .D ( new_AGEMA_signal_5400 ), .Q ( new_AGEMA_signal_5817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C ( clk ), .D ( new_AGEMA_signal_5425 ), .Q ( new_AGEMA_signal_5819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C ( clk ), .D ( new_AGEMA_signal_5426 ), .Q ( new_AGEMA_signal_5821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C ( clk ), .D ( n2417 ), .Q ( new_AGEMA_signal_5823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C ( clk ), .D ( new_AGEMA_signal_1324 ), .Q ( new_AGEMA_signal_5825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C ( clk ), .D ( new_AGEMA_signal_5495 ), .Q ( new_AGEMA_signal_5835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C ( clk ), .D ( new_AGEMA_signal_5496 ), .Q ( new_AGEMA_signal_5837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C ( clk ), .D ( n2483 ), .Q ( new_AGEMA_signal_5839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C ( clk ), .D ( new_AGEMA_signal_1107 ), .Q ( new_AGEMA_signal_5841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C ( clk ), .D ( n2629 ), .Q ( new_AGEMA_signal_5861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C ( clk ), .D ( new_AGEMA_signal_1120 ), .Q ( new_AGEMA_signal_5863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C ( clk ), .D ( n2736 ), .Q ( new_AGEMA_signal_5875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C ( clk ), .D ( new_AGEMA_signal_1051 ), .Q ( new_AGEMA_signal_5877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C ( clk ), .D ( new_AGEMA_signal_5451 ), .Q ( new_AGEMA_signal_5879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C ( clk ), .D ( new_AGEMA_signal_5452 ), .Q ( new_AGEMA_signal_5881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C ( clk ), .D ( new_AGEMA_signal_5423 ), .Q ( new_AGEMA_signal_5883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C ( clk ), .D ( new_AGEMA_signal_5424 ), .Q ( new_AGEMA_signal_5885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C ( clk ), .D ( n2787 ), .Q ( new_AGEMA_signal_5887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C ( clk ), .D ( new_AGEMA_signal_1303 ), .Q ( new_AGEMA_signal_5889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C ( clk ), .D ( new_AGEMA_signal_5899 ), .Q ( new_AGEMA_signal_5900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C ( clk ), .D ( new_AGEMA_signal_5903 ), .Q ( new_AGEMA_signal_5904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C ( clk ), .D ( new_AGEMA_signal_5909 ), .Q ( new_AGEMA_signal_5910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C ( clk ), .D ( new_AGEMA_signal_5913 ), .Q ( new_AGEMA_signal_5914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C ( clk ), .D ( n2009 ), .Q ( new_AGEMA_signal_5917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C ( clk ), .D ( new_AGEMA_signal_1162 ), .Q ( new_AGEMA_signal_5920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C ( clk ), .D ( n2034 ), .Q ( new_AGEMA_signal_5927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_5930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C ( clk ), .D ( new_AGEMA_signal_5493 ), .Q ( new_AGEMA_signal_5935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C ( clk ), .D ( new_AGEMA_signal_5494 ), .Q ( new_AGEMA_signal_5938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C ( clk ), .D ( new_AGEMA_signal_5507 ), .Q ( new_AGEMA_signal_5941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C ( clk ), .D ( new_AGEMA_signal_5508 ), .Q ( new_AGEMA_signal_5944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C ( clk ), .D ( new_AGEMA_signal_5381 ), .Q ( new_AGEMA_signal_5953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C ( clk ), .D ( new_AGEMA_signal_5382 ), .Q ( new_AGEMA_signal_5956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C ( clk ), .D ( n2122 ), .Q ( new_AGEMA_signal_5959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C ( clk ), .D ( new_AGEMA_signal_1193 ), .Q ( new_AGEMA_signal_5962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C ( clk ), .D ( n2220 ), .Q ( new_AGEMA_signal_5967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C ( clk ), .D ( new_AGEMA_signal_1199 ), .Q ( new_AGEMA_signal_5970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C ( clk ), .D ( new_AGEMA_signal_5985 ), .Q ( new_AGEMA_signal_5986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C ( clk ), .D ( new_AGEMA_signal_5989 ), .Q ( new_AGEMA_signal_5990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C ( clk ), .D ( new_AGEMA_signal_5431 ), .Q ( new_AGEMA_signal_5993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C ( clk ), .D ( new_AGEMA_signal_5432 ), .Q ( new_AGEMA_signal_5996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C ( clk ), .D ( n2344 ), .Q ( new_AGEMA_signal_6021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C ( clk ), .D ( new_AGEMA_signal_1239 ), .Q ( new_AGEMA_signal_6024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C ( clk ), .D ( n2468 ), .Q ( new_AGEMA_signal_6053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C ( clk ), .D ( new_AGEMA_signal_1110 ), .Q ( new_AGEMA_signal_6056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C ( clk ), .D ( n2761 ), .Q ( new_AGEMA_signal_6059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C ( clk ), .D ( new_AGEMA_signal_1144 ), .Q ( new_AGEMA_signal_6062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C ( clk ), .D ( new_AGEMA_signal_6071 ), .Q ( new_AGEMA_signal_6072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C ( clk ), .D ( new_AGEMA_signal_6075 ), .Q ( new_AGEMA_signal_6076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C ( clk ), .D ( new_AGEMA_signal_6101 ), .Q ( new_AGEMA_signal_6102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C ( clk ), .D ( new_AGEMA_signal_6105 ), .Q ( new_AGEMA_signal_6106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C ( clk ), .D ( n2825 ), .Q ( new_AGEMA_signal_6117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C ( clk ), .D ( new_AGEMA_signal_1308 ), .Q ( new_AGEMA_signal_6120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C ( clk ), .D ( n1957 ), .Q ( new_AGEMA_signal_6125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C ( clk ), .D ( new_AGEMA_signal_1049 ), .Q ( new_AGEMA_signal_6129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C ( clk ), .D ( n2026 ), .Q ( new_AGEMA_signal_6139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_6143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C ( clk ), .D ( n2811 ), .Q ( new_AGEMA_signal_6159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C ( clk ), .D ( new_AGEMA_signal_1194 ), .Q ( new_AGEMA_signal_6163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C ( clk ), .D ( new_AGEMA_signal_5513 ), .Q ( new_AGEMA_signal_6205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C ( clk ), .D ( new_AGEMA_signal_5514 ), .Q ( new_AGEMA_signal_6209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C ( clk ), .D ( n2363 ), .Q ( new_AGEMA_signal_6223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_6227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C ( clk ), .D ( new_AGEMA_signal_5491 ), .Q ( new_AGEMA_signal_6255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C ( clk ), .D ( new_AGEMA_signal_5492 ), .Q ( new_AGEMA_signal_6259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C ( clk ), .D ( new_AGEMA_signal_5391 ), .Q ( new_AGEMA_signal_6263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C ( clk ), .D ( new_AGEMA_signal_5392 ), .Q ( new_AGEMA_signal_6267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C ( clk ), .D ( n2544 ), .Q ( new_AGEMA_signal_6349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C ( clk ), .D ( new_AGEMA_signal_1079 ), .Q ( new_AGEMA_signal_6354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C ( clk ), .D ( n2364 ), .Q ( new_AGEMA_signal_6399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C ( clk ), .D ( new_AGEMA_signal_1245 ), .Q ( new_AGEMA_signal_6404 ) ) ;

    /* cells in depth 4 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1968 ( .a ({new_AGEMA_signal_1309, n1924}), .b ({new_AGEMA_signal_1310, n1923}), .clk ( clk ), .r ({Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804]}), .c ({new_AGEMA_signal_1470, n1936}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1982 ( .a ({new_AGEMA_signal_5516, new_AGEMA_signal_5515}), .b ({new_AGEMA_signal_1311, n1927}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808]}), .c ({new_AGEMA_signal_1471, n1928}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U1994 ( .a ({new_AGEMA_signal_5518, new_AGEMA_signal_5517}), .b ({new_AGEMA_signal_1312, n1929}), .clk ( clk ), .r ({Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_1472, n1931}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2012 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_1314, n1938}), .clk ( clk ), .r ({Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816]}), .c ({new_AGEMA_signal_1473, n1939}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2024 ( .a ({new_AGEMA_signal_1315, n2235}), .b ({new_AGEMA_signal_1137, n1943}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820]}), .c ({new_AGEMA_signal_1474, n1948}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2032 ( .a ({new_AGEMA_signal_1138, n1946}), .b ({new_AGEMA_signal_1316, n1945}), .clk ( clk ), .r ({Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_1475, n1947}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2041 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5520}), .b ({new_AGEMA_signal_1318, n1951}), .clk ( clk ), .r ({Fresh[1831], Fresh[1830], Fresh[1829], Fresh[1828]}), .c ({new_AGEMA_signal_1476, n1954}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2049 ( .a ({new_AGEMA_signal_5524, new_AGEMA_signal_5523}), .b ({new_AGEMA_signal_1319, n1952}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832]}), .c ({new_AGEMA_signal_1477, n1953}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2058 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525}), .b ({new_AGEMA_signal_1320, n2687}), .clk ( clk ), .r ({Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_1478, n2658}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2065 ( .a ({new_AGEMA_signal_5528, new_AGEMA_signal_5527}), .b ({new_AGEMA_signal_1143, n1963}), .clk ( clk ), .r ({Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840]}), .c ({new_AGEMA_signal_1322, n1965}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2078 ( .a ({new_AGEMA_signal_5530, new_AGEMA_signal_5529}), .b ({new_AGEMA_signal_1480, n1968}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844]}), .c ({new_AGEMA_signal_1591, n1970}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2084 ( .a ({new_AGEMA_signal_1325, n2684}), .b ({new_AGEMA_signal_5532, new_AGEMA_signal_5531}), .clk ( clk ), .r ({Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_1481, n1969}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2093 ( .a ({new_AGEMA_signal_1326, n1972}), .b ({new_AGEMA_signal_1149, n1971}), .clk ( clk ), .r ({Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852]}), .c ({new_AGEMA_signal_1482, n1978}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2102 ( .a ({new_AGEMA_signal_1327, n1974}), .b ({new_AGEMA_signal_5534, new_AGEMA_signal_5533}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856]}), .c ({new_AGEMA_signal_1483, n1975}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2107 ( .a ({new_AGEMA_signal_5536, new_AGEMA_signal_5535}), .b ({new_AGEMA_signal_1328, n1979}), .clk ( clk ), .r ({Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_1484, n1980}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2114 ( .a ({new_AGEMA_signal_1152, n1985}), .b ({new_AGEMA_signal_5538, new_AGEMA_signal_5537}), .clk ( clk ), .r ({Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864]}), .c ({new_AGEMA_signal_1329, n1986}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2124 ( .a ({new_AGEMA_signal_1330, n1994}), .b ({new_AGEMA_signal_5540, new_AGEMA_signal_5539}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868]}), .c ({new_AGEMA_signal_1486, n1997}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2137 ( .a ({new_AGEMA_signal_5542, new_AGEMA_signal_5541}), .b ({new_AGEMA_signal_1332, n2137}), .clk ( clk ), .r ({Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_1487, n2012}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2145 ( .a ({new_AGEMA_signal_1333, n2006}), .b ({new_AGEMA_signal_1334, n2005}), .clk ( clk ), .r ({Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876]}), .c ({new_AGEMA_signal_1488, n2007}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2161 ( .s ({new_AGEMA_signal_5544, new_AGEMA_signal_5543}), .b ({new_AGEMA_signal_1165, n2020}), .a ({new_AGEMA_signal_5548, new_AGEMA_signal_5546}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880]}), .c ({new_AGEMA_signal_1336, n2021}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2176 ( .a ({new_AGEMA_signal_5550, new_AGEMA_signal_5549}), .b ({new_AGEMA_signal_1338, n2031}), .clk ( clk ), .r ({Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_1490, n2032}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2185 ( .a ({new_AGEMA_signal_5552, new_AGEMA_signal_5551}), .b ({new_AGEMA_signal_1339, n2040}), .clk ( clk ), .r ({Fresh[1891], Fresh[1890], Fresh[1889], Fresh[1888]}), .c ({new_AGEMA_signal_1491, n2041}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2189 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_5554, new_AGEMA_signal_5553}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892]}), .c ({new_AGEMA_signal_1492, n2043}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2194 ( .a ({new_AGEMA_signal_5556, new_AGEMA_signal_5555}), .b ({new_AGEMA_signal_1340, n2045}), .clk ( clk ), .r ({Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_1493, n2046}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2204 ( .s ({new_AGEMA_signal_5544, new_AGEMA_signal_5543}), .b ({new_AGEMA_signal_1342, n2056}), .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557}), .clk ( clk ), .r ({Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900]}), .c ({new_AGEMA_signal_1494, n2058}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2210 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559}), .b ({new_AGEMA_signal_1343, n2060}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904]}), .c ({new_AGEMA_signal_1495, n2063}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2218 ( .a ({new_AGEMA_signal_1344, n2066}), .b ({new_AGEMA_signal_1345, n2065}), .clk ( clk ), .r ({Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_1496, n2652}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2227 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561}), .b ({new_AGEMA_signal_1347, n2074}), .clk ( clk ), .r ({Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912]}), .c ({new_AGEMA_signal_1497, n2076}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2236 ( .a ({new_AGEMA_signal_5566, new_AGEMA_signal_5564}), .b ({new_AGEMA_signal_1348, n2082}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916]}), .c ({new_AGEMA_signal_1498, n2105}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2241 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567}), .b ({new_AGEMA_signal_1349, n2084}), .clk ( clk ), .r ({Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_1499, n2099}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2243 ( .a ({new_AGEMA_signal_1350, n2085}), .b ({new_AGEMA_signal_5570, new_AGEMA_signal_5569}), .clk ( clk ), .r ({Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924]}), .c ({new_AGEMA_signal_1500, n2091}) ) ;
    and_GHPC #(.low_latency(1), .pipeline(1)) U2246 ( .a ({new_AGEMA_signal_5572, new_AGEMA_signal_5571}), .b ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928]}), .c ({new_AGEMA_signal_1501, n2090}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2253 ( .a ({new_AGEMA_signal_5574, new_AGEMA_signal_5573}), .b ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .r ({Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_1502, n2093}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2262 ( .a ({new_AGEMA_signal_5576, new_AGEMA_signal_5575}), .b ({new_AGEMA_signal_1356, n2160}), .clk ( clk ), .r ({Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936]}), .c ({new_AGEMA_signal_1503, n2102}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2266 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_5580, new_AGEMA_signal_5578}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940]}), .c ({new_AGEMA_signal_1357, n2106}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2272 ( .a ({new_AGEMA_signal_5582, new_AGEMA_signal_5581}), .b ({new_AGEMA_signal_1504, n2114}), .clk ( clk ), .r ({Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_1606, n2116}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2282 ( .a ({new_AGEMA_signal_1358, n2291}), .b ({new_AGEMA_signal_1192, n2119}), .clk ( clk ), .r ({Fresh[1951], Fresh[1950], Fresh[1949], Fresh[1948]}), .c ({new_AGEMA_signal_1505, n2120}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2293 ( .a ({new_AGEMA_signal_1195, n2130}), .b ({new_AGEMA_signal_1196, n2129}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952]}), .c ({new_AGEMA_signal_1359, n2155}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2296 ( .a ({new_AGEMA_signal_5584, new_AGEMA_signal_5583}), .b ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .r ({Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_1506, n2543}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2299 ( .a ({new_AGEMA_signal_1198, n2133}), .b ({new_AGEMA_signal_5586, new_AGEMA_signal_5585}), .clk ( clk ), .r ({Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960]}), .c ({new_AGEMA_signal_1360, n2134}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2303 ( .a ({new_AGEMA_signal_1332, n2137}), .b ({new_AGEMA_signal_1361, n2136}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964]}), .c ({new_AGEMA_signal_1508, n2143}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2308 ( .a ({new_AGEMA_signal_1362, n2139}), .b ({new_AGEMA_signal_5590, new_AGEMA_signal_5588}), .clk ( clk ), .r ({Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_1509, n2140}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2324 ( .a ({new_AGEMA_signal_1366, n2157}), .b ({new_AGEMA_signal_5592, new_AGEMA_signal_5591}), .clk ( clk ), .r ({Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972]}), .c ({new_AGEMA_signal_1510, n2159}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2326 ( .a ({new_AGEMA_signal_1356, n2160}), .b ({new_AGEMA_signal_5594, new_AGEMA_signal_5593}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976]}), .c ({new_AGEMA_signal_1511, n2161}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2330 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5520}), .b ({new_AGEMA_signal_1203, n2163}), .clk ( clk ), .r ({Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_1367, n2164}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2345 ( .a ({new_AGEMA_signal_5596, new_AGEMA_signal_5595}), .b ({new_AGEMA_signal_1370, n2177}), .clk ( clk ), .r ({Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984]}), .c ({new_AGEMA_signal_1513, n2179}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2359 ( .a ({new_AGEMA_signal_5600, new_AGEMA_signal_5598}), .b ({new_AGEMA_signal_1373, n2191}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988]}), .c ({new_AGEMA_signal_1514, n2192}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2370 ( .a ({new_AGEMA_signal_1374, n2201}), .b ({new_AGEMA_signal_1515, n2200}), .clk ( clk ), .r ({Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_1613, n2203}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2382 ( .a ({new_AGEMA_signal_1376, n2217}), .b ({new_AGEMA_signal_1210, n2216}), .clk ( clk ), .r ({Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996]}), .c ({new_AGEMA_signal_1517, n2224}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2388 ( .a ({new_AGEMA_signal_1377, n2222}), .b ({new_AGEMA_signal_1378, n2221}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000]}), .c ({new_AGEMA_signal_1518, n2223}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2392 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1213, n2226}), .clk ( clk ), .r ({Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_1379, n2229}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2399 ( .a ({new_AGEMA_signal_5524, new_AGEMA_signal_5523}), .b ({new_AGEMA_signal_1520, n2233}), .clk ( clk ), .r ({Fresh[2011], Fresh[2010], Fresh[2009], Fresh[2008]}), .c ({new_AGEMA_signal_1616, n2234}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2410 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525}), .b ({new_AGEMA_signal_1381, n2244}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012]}), .c ({new_AGEMA_signal_1521, n2246}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2418 ( .a ({new_AGEMA_signal_5602, new_AGEMA_signal_5601}), .b ({new_AGEMA_signal_1383, n2253}), .clk ( clk ), .r ({Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_1522, n2254}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2425 ( .a ({new_AGEMA_signal_5604, new_AGEMA_signal_5603}), .b ({new_AGEMA_signal_1384, n2260}), .clk ( clk ), .r ({Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020]}), .c ({new_AGEMA_signal_1523, n2263}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2434 ( .a ({new_AGEMA_signal_5606, new_AGEMA_signal_5605}), .b ({new_AGEMA_signal_1223, n2265}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024]}), .c ({new_AGEMA_signal_1385, n2267}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2438 ( .a ({new_AGEMA_signal_5524, new_AGEMA_signal_5523}), .b ({new_AGEMA_signal_1224, n2269}), .clk ( clk ), .r ({Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_1386, n2270}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2445 ( .a ({new_AGEMA_signal_5608, new_AGEMA_signal_5607}), .b ({new_AGEMA_signal_1226, n2277}), .clk ( clk ), .r ({Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032]}), .c ({new_AGEMA_signal_1387, n2279}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2450 ( .a ({new_AGEMA_signal_5548, new_AGEMA_signal_5546}), .b ({new_AGEMA_signal_1227, n2282}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036]}), .c ({new_AGEMA_signal_1388, n2283}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2453 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567}), .b ({new_AGEMA_signal_1389, n2284}), .clk ( clk ), .r ({Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_1528, n2285}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2457 ( .a ({new_AGEMA_signal_5522, new_AGEMA_signal_5520}), .b ({new_AGEMA_signal_1390, n2459}), .clk ( clk ), .r ({Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044]}), .c ({new_AGEMA_signal_1529, n2686}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2460 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525}), .b ({new_AGEMA_signal_1391, n2288}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048]}), .c ({new_AGEMA_signal_1530, n2289}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2463 ( .a ({new_AGEMA_signal_1392, n2458}), .b ({new_AGEMA_signal_5610, new_AGEMA_signal_5609}), .clk ( clk ), .r ({Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_1531, n2297}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2465 ( .a ({new_AGEMA_signal_5612, new_AGEMA_signal_5611}), .b ({new_AGEMA_signal_1358, n2291}), .clk ( clk ), .r ({Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056]}), .c ({new_AGEMA_signal_1532, n2292}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2473 ( .a ({new_AGEMA_signal_5614, new_AGEMA_signal_5613}), .b ({new_AGEMA_signal_1394, n2300}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060]}), .c ({new_AGEMA_signal_1533, n2301}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2483 ( .a ({new_AGEMA_signal_5616, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_1396, n2314}), .clk ( clk ), .r ({Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_1534, n2321}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2487 ( .a ({new_AGEMA_signal_1097, n2319}), .b ({new_AGEMA_signal_5618, new_AGEMA_signal_5617}), .clk ( clk ), .r ({Fresh[2071], Fresh[2070], Fresh[2069], Fresh[2068]}), .c ({new_AGEMA_signal_1233, n2320}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2493 ( .a ({new_AGEMA_signal_1234, n2326}), .b ({new_AGEMA_signal_5620, new_AGEMA_signal_5619}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072]}), .c ({new_AGEMA_signal_1397, n2334}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2497 ( .a ({new_AGEMA_signal_1398, n2329}), .b ({new_AGEMA_signal_5548, new_AGEMA_signal_5546}), .clk ( clk ), .r ({Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_1535, n2332}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2498 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621}), .b ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .r ({Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080]}), .c ({new_AGEMA_signal_1536, n2331}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2502 ( .a ({new_AGEMA_signal_5624, new_AGEMA_signal_5623}), .b ({new_AGEMA_signal_1537, n2335}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084]}), .c ({new_AGEMA_signal_1626, n2336}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2508 ( .a ({new_AGEMA_signal_1399, n2341}), .b ({new_AGEMA_signal_1238, n2340}), .clk ( clk ), .r ({Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_1538, n2342}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2519 ( .a ({new_AGEMA_signal_1242, n2352}), .b ({new_AGEMA_signal_5626, new_AGEMA_signal_5625}), .clk ( clk ), .r ({Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092]}), .c ({new_AGEMA_signal_1400, n2367}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2523 ( .a ({new_AGEMA_signal_1401, n2354}), .b ({new_AGEMA_signal_5628, new_AGEMA_signal_5627}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096]}), .c ({new_AGEMA_signal_1539, n2358}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2547 ( .a ({new_AGEMA_signal_1247, n2385}), .b ({new_AGEMA_signal_1248, n2384}), .clk ( clk ), .r ({Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_1406, n2387}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2555 ( .a ({new_AGEMA_signal_1250, n2391}), .b ({new_AGEMA_signal_1408, n2390}), .clk ( clk ), .r ({Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104]}), .c ({new_AGEMA_signal_1542, n2392}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2566 ( .a ({new_AGEMA_signal_1252, n2403}), .b ({new_AGEMA_signal_5630, new_AGEMA_signal_5629}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108]}), .c ({new_AGEMA_signal_1410, n2404}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2570 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559}), .b ({new_AGEMA_signal_1411, n2408}), .clk ( clk ), .r ({Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_1544, n2409}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2575 ( .a ({new_AGEMA_signal_1412, n2574}), .b ({new_AGEMA_signal_1253, n2413}), .clk ( clk ), .r ({Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116]}), .c ({new_AGEMA_signal_1545, n2414}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2578 ( .a ({new_AGEMA_signal_5632, new_AGEMA_signal_5631}), .b ({new_AGEMA_signal_1254, n2416}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120]}), .c ({new_AGEMA_signal_1413, n2418}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2589 ( .a ({new_AGEMA_signal_1415, n2689}), .b ({new_AGEMA_signal_5634, new_AGEMA_signal_5633}), .clk ( clk ), .r ({Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_1547, n2432}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2592 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5637}), .b ({new_AGEMA_signal_1257, n2434}), .clk ( clk ), .r ({Fresh[2131], Fresh[2130], Fresh[2129], Fresh[2128]}), .c ({new_AGEMA_signal_1416, n2435}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2601 ( .a ({new_AGEMA_signal_1418, n2445}), .b ({new_AGEMA_signal_1419, n2444}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132]}), .c ({new_AGEMA_signal_1548, n2449}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2603 ( .a ({new_AGEMA_signal_5616, new_AGEMA_signal_5615}), .b ({new_AGEMA_signal_1420, n2447}), .clk ( clk ), .r ({Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_1549, n2448}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2609 ( .a ({new_AGEMA_signal_1421, n2454}), .b ({new_AGEMA_signal_5642, new_AGEMA_signal_5641}), .clk ( clk ), .r ({Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140]}), .c ({new_AGEMA_signal_1550, n2455}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2612 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_1392, n2458}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144]}), .c ({new_AGEMA_signal_1551, n2460}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2618 ( .a ({new_AGEMA_signal_5612, new_AGEMA_signal_5611}), .b ({new_AGEMA_signal_1260, n2465}), .clk ( clk ), .r ({Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_1422, n2466}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2629 ( .a ({new_AGEMA_signal_1262, n2476}), .b ({new_AGEMA_signal_5644, new_AGEMA_signal_5643}), .clk ( clk ), .r ({Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152]}), .c ({new_AGEMA_signal_1423, n2477}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2634 ( .a ({new_AGEMA_signal_5558, new_AGEMA_signal_5557}), .b ({new_AGEMA_signal_1424, n2481}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156]}), .c ({new_AGEMA_signal_1554, n2482}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2640 ( .a ({new_AGEMA_signal_5646, new_AGEMA_signal_5645}), .b ({new_AGEMA_signal_1265, n2486}), .clk ( clk ), .r ({Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_1425, n2490}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2648 ( .a ({new_AGEMA_signal_1268, n2495}), .b ({new_AGEMA_signal_1426, n2494}), .clk ( clk ), .r ({Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164]}), .c ({new_AGEMA_signal_1556, n2496}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2654 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1557, n2503}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168]}), .c ({new_AGEMA_signal_1643, n2507}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2664 ( .a ({new_AGEMA_signal_1428, n2518}), .b ({new_AGEMA_signal_1558, n2517}), .clk ( clk ), .r ({Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_1644, n2525}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2669 ( .a ({new_AGEMA_signal_1429, n2523}), .b ({new_AGEMA_signal_1430, n2522}), .clk ( clk ), .r ({Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176]}), .c ({new_AGEMA_signal_1559, n2524}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2676 ( .a ({new_AGEMA_signal_1431, n2532}), .b ({new_AGEMA_signal_5650, new_AGEMA_signal_5648}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180]}), .c ({new_AGEMA_signal_1560, n2537}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2678 ( .a ({new_AGEMA_signal_5560, new_AGEMA_signal_5559}), .b ({new_AGEMA_signal_1432, n2534}), .clk ( clk ), .r ({Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_1561, n2536}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2684 ( .a ({new_AGEMA_signal_5652, new_AGEMA_signal_5651}), .b ({new_AGEMA_signal_1272, n2546}), .clk ( clk ), .r ({Fresh[2191], Fresh[2190], Fresh[2189], Fresh[2188]}), .c ({new_AGEMA_signal_1434, n2547}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2693 ( .a ({new_AGEMA_signal_5654, new_AGEMA_signal_5653}), .b ({new_AGEMA_signal_1437, n2556}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192]}), .c ({new_AGEMA_signal_1562, n2557}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2699 ( .a ({new_AGEMA_signal_1439, n2715}), .b ({new_AGEMA_signal_5656, new_AGEMA_signal_5655}), .clk ( clk ), .r ({Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_1563, n2565}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2704 ( .a ({new_AGEMA_signal_1412, n2574}), .b ({new_AGEMA_signal_1440, n2573}), .clk ( clk ), .r ({Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200]}), .c ({new_AGEMA_signal_1564, n2591}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2709 ( .a ({new_AGEMA_signal_1442, n2579}), .b ({new_AGEMA_signal_1277, n2578}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204]}), .c ({new_AGEMA_signal_1565, n2580}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2727 ( .a ({new_AGEMA_signal_1118, n2601}), .b ({new_AGEMA_signal_5660, new_AGEMA_signal_5658}), .clk ( clk ), .r ({Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_1282, n2602}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2738 ( .a ({new_AGEMA_signal_1448, n2618}), .b ({new_AGEMA_signal_5662, new_AGEMA_signal_5661}), .clk ( clk ), .r ({Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212]}), .c ({new_AGEMA_signal_1567, n2619}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2744 ( .a ({new_AGEMA_signal_5570, new_AGEMA_signal_5569}), .b ({new_AGEMA_signal_1449, n2626}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216]}), .c ({new_AGEMA_signal_1568, n2628}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2753 ( .a ({new_AGEMA_signal_1450, n2644}), .b ({new_AGEMA_signal_5584, new_AGEMA_signal_5583}), .clk ( clk ), .r ({Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_1569, n2649}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2755 ( .a ({new_AGEMA_signal_5664, new_AGEMA_signal_5663}), .b ({new_AGEMA_signal_1288, n2646}), .clk ( clk ), .r ({Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224]}), .c ({new_AGEMA_signal_1451, n2648}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2765 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525}), .b ({new_AGEMA_signal_1453, n2663}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228]}), .c ({new_AGEMA_signal_1570, n2664}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2771 ( .a ({new_AGEMA_signal_1290, n2675}), .b ({new_AGEMA_signal_5666, new_AGEMA_signal_5665}), .clk ( clk ), .r ({Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_1571, n2681}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2773 ( .a ({new_AGEMA_signal_5592, new_AGEMA_signal_5591}), .b ({new_AGEMA_signal_1291, n2678}), .clk ( clk ), .r ({Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236]}), .c ({new_AGEMA_signal_1454, n2680}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2776 ( .a ({new_AGEMA_signal_1325, n2684}), .b ({new_AGEMA_signal_5668, new_AGEMA_signal_5667}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240]}), .c ({new_AGEMA_signal_1572, n2685}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2778 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651}), .clk ( clk ), .r ({Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_1573, n2698}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2779 ( .a ({new_AGEMA_signal_1415, n2689}), .b ({new_AGEMA_signal_5654, new_AGEMA_signal_5653}), .clk ( clk ), .r ({Fresh[2251], Fresh[2250], Fresh[2249], Fresh[2248]}), .c ({new_AGEMA_signal_1574, n2692}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2793 ( .a ({new_AGEMA_signal_1439, n2715}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252]}), .c ({new_AGEMA_signal_1575, n2716}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2800 ( .a ({new_AGEMA_signal_1296, n2727}), .b ({new_AGEMA_signal_5672, new_AGEMA_signal_5671}), .clk ( clk ), .r ({Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_1457, n2728}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2804 ( .a ({new_AGEMA_signal_5674, new_AGEMA_signal_5673}), .b ({new_AGEMA_signal_1458, n2733}), .clk ( clk ), .r ({Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260]}), .c ({new_AGEMA_signal_1577, n2735}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2808 ( .a ({new_AGEMA_signal_5538, new_AGEMA_signal_5537}), .b ({new_AGEMA_signal_1459, n2740}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264]}), .c ({new_AGEMA_signal_1578, n2743}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2813 ( .a ({new_AGEMA_signal_5678, new_AGEMA_signal_5676}), .b ({new_AGEMA_signal_1299, n2749}), .clk ( clk ), .r ({Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_1460, n2751}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2817 ( .a ({new_AGEMA_signal_1461, n2757}), .b ({new_AGEMA_signal_1300, n2756}), .clk ( clk ), .r ({Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272]}), .c ({new_AGEMA_signal_1579, n2758}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2820 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679}), .b ({new_AGEMA_signal_1462, n2762}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276]}), .c ({new_AGEMA_signal_1580, n2764}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2827 ( .a ({new_AGEMA_signal_1464, n2776}), .b ({new_AGEMA_signal_1465, n2775}), .clk ( clk ), .r ({Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_1581, n2800}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2831 ( .a ({new_AGEMA_signal_5682, new_AGEMA_signal_5681}), .b ({new_AGEMA_signal_1302, n2783}), .clk ( clk ), .r ({Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284]}), .c ({new_AGEMA_signal_1466, n2788}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2837 ( .a ({new_AGEMA_signal_5686, new_AGEMA_signal_5684}), .b ({new_AGEMA_signal_1467, n2795}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288]}), .c ({new_AGEMA_signal_1583, n2797}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2846 ( .a ({new_AGEMA_signal_1468, n2814}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543}), .clk ( clk ), .r ({Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_1584, n2822}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2849 ( .a ({new_AGEMA_signal_5688, new_AGEMA_signal_5687}), .b ({new_AGEMA_signal_1307, n2819}), .clk ( clk ), .r ({Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296]}), .c ({new_AGEMA_signal_1469, n2821}) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C ( clk ), .D ( new_AGEMA_signal_5689 ), .Q ( new_AGEMA_signal_5690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C ( clk ), .D ( new_AGEMA_signal_5691 ), .Q ( new_AGEMA_signal_5692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C ( clk ), .D ( new_AGEMA_signal_5693 ), .Q ( new_AGEMA_signal_5694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C ( clk ), .D ( new_AGEMA_signal_5695 ), .Q ( new_AGEMA_signal_5696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C ( clk ), .D ( new_AGEMA_signal_5651 ), .Q ( new_AGEMA_signal_5697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C ( clk ), .D ( new_AGEMA_signal_5652 ), .Q ( new_AGEMA_signal_5698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C ( clk ), .D ( n1966 ), .Q ( new_AGEMA_signal_5699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C ( clk ), .D ( new_AGEMA_signal_1321 ), .Q ( new_AGEMA_signal_5700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C ( clk ), .D ( new_AGEMA_signal_5701 ), .Q ( new_AGEMA_signal_5702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C ( clk ), .D ( new_AGEMA_signal_5703 ), .Q ( new_AGEMA_signal_5704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C ( clk ), .D ( new_AGEMA_signal_5615 ), .Q ( new_AGEMA_signal_5705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C ( clk ), .D ( new_AGEMA_signal_5616 ), .Q ( new_AGEMA_signal_5706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C ( clk ), .D ( new_AGEMA_signal_5707 ), .Q ( new_AGEMA_signal_5708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C ( clk ), .D ( new_AGEMA_signal_5709 ), .Q ( new_AGEMA_signal_5710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C ( clk ), .D ( n1996 ), .Q ( new_AGEMA_signal_5711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C ( clk ), .D ( new_AGEMA_signal_1331 ), .Q ( new_AGEMA_signal_5712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C ( clk ), .D ( new_AGEMA_signal_5713 ), .Q ( new_AGEMA_signal_5714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C ( clk ), .D ( new_AGEMA_signal_5715 ), .Q ( new_AGEMA_signal_5716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C ( clk ), .D ( new_AGEMA_signal_5717 ), .Q ( new_AGEMA_signal_5718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C ( clk ), .D ( new_AGEMA_signal_5719 ), .Q ( new_AGEMA_signal_5720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C ( clk ), .D ( n2033 ), .Q ( new_AGEMA_signal_5721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C ( clk ), .D ( new_AGEMA_signal_1337 ), .Q ( new_AGEMA_signal_5722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C ( clk ), .D ( new_AGEMA_signal_5571 ), .Q ( new_AGEMA_signal_5723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C ( clk ), .D ( new_AGEMA_signal_5572 ), .Q ( new_AGEMA_signal_5724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C ( clk ), .D ( new_AGEMA_signal_5581 ), .Q ( new_AGEMA_signal_5725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C ( clk ), .D ( new_AGEMA_signal_5582 ), .Q ( new_AGEMA_signal_5726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C ( clk ), .D ( new_AGEMA_signal_5609 ), .Q ( new_AGEMA_signal_5727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C ( clk ), .D ( new_AGEMA_signal_5610 ), .Q ( new_AGEMA_signal_5728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C ( clk ), .D ( new_AGEMA_signal_5729 ), .Q ( new_AGEMA_signal_5730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C ( clk ), .D ( new_AGEMA_signal_5731 ), .Q ( new_AGEMA_signal_5732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C ( clk ), .D ( new_AGEMA_signal_5733 ), .Q ( new_AGEMA_signal_5734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C ( clk ), .D ( new_AGEMA_signal_5735 ), .Q ( new_AGEMA_signal_5736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C ( clk ), .D ( new_AGEMA_signal_5737 ), .Q ( new_AGEMA_signal_5738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C ( clk ), .D ( new_AGEMA_signal_5739 ), .Q ( new_AGEMA_signal_5740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C ( clk ), .D ( n2089 ), .Q ( new_AGEMA_signal_5741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C ( clk ), .D ( new_AGEMA_signal_1352 ), .Q ( new_AGEMA_signal_5742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C ( clk ), .D ( n2092 ), .Q ( new_AGEMA_signal_5743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_5744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C ( clk ), .D ( n2115 ), .Q ( new_AGEMA_signal_5745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C ( clk ), .D ( new_AGEMA_signal_1190 ), .Q ( new_AGEMA_signal_5746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C ( clk ), .D ( new_AGEMA_signal_5747 ), .Q ( new_AGEMA_signal_5748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C ( clk ), .D ( new_AGEMA_signal_5749 ), .Q ( new_AGEMA_signal_5750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C ( clk ), .D ( n2687 ), .Q ( new_AGEMA_signal_5751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C ( clk ), .D ( new_AGEMA_signal_1320 ), .Q ( new_AGEMA_signal_5752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C ( clk ), .D ( new_AGEMA_signal_5753 ), .Q ( new_AGEMA_signal_5754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C ( clk ), .D ( new_AGEMA_signal_5755 ), .Q ( new_AGEMA_signal_5756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C ( clk ), .D ( new_AGEMA_signal_5758 ), .Q ( new_AGEMA_signal_5759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C ( clk ), .D ( new_AGEMA_signal_5761 ), .Q ( new_AGEMA_signal_5762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C ( clk ), .D ( new_AGEMA_signal_5763 ), .Q ( new_AGEMA_signal_5764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C ( clk ), .D ( new_AGEMA_signal_5765 ), .Q ( new_AGEMA_signal_5766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C ( clk ), .D ( new_AGEMA_signal_5767 ), .Q ( new_AGEMA_signal_5768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C ( clk ), .D ( new_AGEMA_signal_5769 ), .Q ( new_AGEMA_signal_5770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C ( clk ), .D ( n2193 ), .Q ( new_AGEMA_signal_5771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_5772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C ( clk ), .D ( n2202 ), .Q ( new_AGEMA_signal_5773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C ( clk ), .D ( new_AGEMA_signal_1516 ), .Q ( new_AGEMA_signal_5774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C ( clk ), .D ( n2228 ), .Q ( new_AGEMA_signal_5775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C ( clk ), .D ( new_AGEMA_signal_1214 ), .Q ( new_AGEMA_signal_5776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C ( clk ), .D ( n2235 ), .Q ( new_AGEMA_signal_5777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C ( clk ), .D ( new_AGEMA_signal_1315 ), .Q ( new_AGEMA_signal_5778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C ( clk ), .D ( new_AGEMA_signal_5779 ), .Q ( new_AGEMA_signal_5780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C ( clk ), .D ( new_AGEMA_signal_5781 ), .Q ( new_AGEMA_signal_5782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C ( clk ), .D ( new_AGEMA_signal_5784 ), .Q ( new_AGEMA_signal_5785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C ( clk ), .D ( new_AGEMA_signal_5787 ), .Q ( new_AGEMA_signal_5788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C ( clk ), .D ( new_AGEMA_signal_5789 ), .Q ( new_AGEMA_signal_5790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C ( clk ), .D ( new_AGEMA_signal_5791 ), .Q ( new_AGEMA_signal_5792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C ( clk ), .D ( n2752 ), .Q ( new_AGEMA_signal_5793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C ( clk ), .D ( new_AGEMA_signal_1525 ), .Q ( new_AGEMA_signal_5794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C ( clk ), .D ( new_AGEMA_signal_5637 ), .Q ( new_AGEMA_signal_5795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C ( clk ), .D ( new_AGEMA_signal_5640 ), .Q ( new_AGEMA_signal_5796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C ( clk ), .D ( n2293 ), .Q ( new_AGEMA_signal_5797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C ( clk ), .D ( new_AGEMA_signal_1393 ), .Q ( new_AGEMA_signal_5798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C ( clk ), .D ( new_AGEMA_signal_5799 ), .Q ( new_AGEMA_signal_5800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C ( clk ), .D ( new_AGEMA_signal_5801 ), .Q ( new_AGEMA_signal_5802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C ( clk ), .D ( n2357 ), .Q ( new_AGEMA_signal_5803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C ( clk ), .D ( new_AGEMA_signal_1402 ), .Q ( new_AGEMA_signal_5804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C ( clk ), .D ( n2386 ), .Q ( new_AGEMA_signal_5805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C ( clk ), .D ( new_AGEMA_signal_1407 ), .Q ( new_AGEMA_signal_5806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C ( clk ), .D ( new_AGEMA_signal_5807 ), .Q ( new_AGEMA_signal_5808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C ( clk ), .D ( new_AGEMA_signal_5809 ), .Q ( new_AGEMA_signal_5810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C ( clk ), .D ( new_AGEMA_signal_5811 ), .Q ( new_AGEMA_signal_5812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C ( clk ), .D ( new_AGEMA_signal_5813 ), .Q ( new_AGEMA_signal_5814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C ( clk ), .D ( new_AGEMA_signal_5815 ), .Q ( new_AGEMA_signal_5816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C ( clk ), .D ( new_AGEMA_signal_5817 ), .Q ( new_AGEMA_signal_5818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C ( clk ), .D ( new_AGEMA_signal_5819 ), .Q ( new_AGEMA_signal_5820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C ( clk ), .D ( new_AGEMA_signal_5821 ), .Q ( new_AGEMA_signal_5822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C ( clk ), .D ( new_AGEMA_signal_5823 ), .Q ( new_AGEMA_signal_5824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C ( clk ), .D ( new_AGEMA_signal_5825 ), .Q ( new_AGEMA_signal_5826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C ( clk ), .D ( n2433 ), .Q ( new_AGEMA_signal_5827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C ( clk ), .D ( new_AGEMA_signal_1414 ), .Q ( new_AGEMA_signal_5828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C ( clk ), .D ( new_AGEMA_signal_5578 ), .Q ( new_AGEMA_signal_5829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C ( clk ), .D ( new_AGEMA_signal_5580 ), .Q ( new_AGEMA_signal_5830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C ( clk ), .D ( n2459 ), .Q ( new_AGEMA_signal_5831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C ( clk ), .D ( new_AGEMA_signal_1390 ), .Q ( new_AGEMA_signal_5832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C ( clk ), .D ( n2467 ), .Q ( new_AGEMA_signal_5833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C ( clk ), .D ( new_AGEMA_signal_1246 ), .Q ( new_AGEMA_signal_5834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C ( clk ), .D ( new_AGEMA_signal_5835 ), .Q ( new_AGEMA_signal_5836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C ( clk ), .D ( new_AGEMA_signal_5837 ), .Q ( new_AGEMA_signal_5838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C ( clk ), .D ( new_AGEMA_signal_5839 ), .Q ( new_AGEMA_signal_5840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C ( clk ), .D ( new_AGEMA_signal_5841 ), .Q ( new_AGEMA_signal_5842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C ( clk ), .D ( n2489 ), .Q ( new_AGEMA_signal_5843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C ( clk ), .D ( new_AGEMA_signal_1266 ), .Q ( new_AGEMA_signal_5844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C ( clk ), .D ( n2497 ), .Q ( new_AGEMA_signal_5845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C ( clk ), .D ( new_AGEMA_signal_1267 ), .Q ( new_AGEMA_signal_5846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C ( clk ), .D ( n2506 ), .Q ( new_AGEMA_signal_5847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C ( clk ), .D ( new_AGEMA_signal_1427 ), .Q ( new_AGEMA_signal_5848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C ( clk ), .D ( n2542 ), .Q ( new_AGEMA_signal_5849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C ( clk ), .D ( new_AGEMA_signal_1433 ), .Q ( new_AGEMA_signal_5850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C ( clk ), .D ( n2558 ), .Q ( new_AGEMA_signal_5851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C ( clk ), .D ( new_AGEMA_signal_1436 ), .Q ( new_AGEMA_signal_5852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C ( clk ), .D ( n2566 ), .Q ( new_AGEMA_signal_5853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_5854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C ( clk ), .D ( n2581 ), .Q ( new_AGEMA_signal_5855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C ( clk ), .D ( new_AGEMA_signal_1276 ), .Q ( new_AGEMA_signal_5856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C ( clk ), .D ( n2603 ), .Q ( new_AGEMA_signal_5857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_5858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C ( clk ), .D ( n2620 ), .Q ( new_AGEMA_signal_5859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C ( clk ), .D ( new_AGEMA_signal_1447 ), .Q ( new_AGEMA_signal_5860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C ( clk ), .D ( new_AGEMA_signal_5861 ), .Q ( new_AGEMA_signal_5862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C ( clk ), .D ( new_AGEMA_signal_5863 ), .Q ( new_AGEMA_signal_5864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C ( clk ), .D ( n2653 ), .Q ( new_AGEMA_signal_5865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C ( clk ), .D ( new_AGEMA_signal_1289 ), .Q ( new_AGEMA_signal_5866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C ( clk ), .D ( n2665 ), .Q ( new_AGEMA_signal_5867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C ( clk ), .D ( new_AGEMA_signal_1313 ), .Q ( new_AGEMA_signal_5868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C ( clk ), .D ( n2691 ), .Q ( new_AGEMA_signal_5869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C ( clk ), .D ( new_AGEMA_signal_1292 ), .Q ( new_AGEMA_signal_5870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C ( clk ), .D ( n2717 ), .Q ( new_AGEMA_signal_5871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C ( clk ), .D ( new_AGEMA_signal_1456 ), .Q ( new_AGEMA_signal_5872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C ( clk ), .D ( n2729 ), .Q ( new_AGEMA_signal_5873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C ( clk ), .D ( new_AGEMA_signal_1576 ), .Q ( new_AGEMA_signal_5874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C ( clk ), .D ( new_AGEMA_signal_5875 ), .Q ( new_AGEMA_signal_5876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C ( clk ), .D ( new_AGEMA_signal_5877 ), .Q ( new_AGEMA_signal_5878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C ( clk ), .D ( new_AGEMA_signal_5879 ), .Q ( new_AGEMA_signal_5880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C ( clk ), .D ( new_AGEMA_signal_5881 ), .Q ( new_AGEMA_signal_5882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C ( clk ), .D ( new_AGEMA_signal_5883 ), .Q ( new_AGEMA_signal_5884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C ( clk ), .D ( new_AGEMA_signal_5885 ), .Q ( new_AGEMA_signal_5886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C ( clk ), .D ( new_AGEMA_signal_5887 ), .Q ( new_AGEMA_signal_5888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C ( clk ), .D ( new_AGEMA_signal_5889 ), .Q ( new_AGEMA_signal_5890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C ( clk ), .D ( new_AGEMA_signal_5623 ), .Q ( new_AGEMA_signal_5891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C ( clk ), .D ( new_AGEMA_signal_5624 ), .Q ( new_AGEMA_signal_5893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C ( clk ), .D ( n1956 ), .Q ( new_AGEMA_signal_5895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C ( clk ), .D ( new_AGEMA_signal_1317 ), .Q ( new_AGEMA_signal_5897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C ( clk ), .D ( new_AGEMA_signal_5900 ), .Q ( new_AGEMA_signal_5901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C ( clk ), .D ( new_AGEMA_signal_5904 ), .Q ( new_AGEMA_signal_5905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C ( clk ), .D ( new_AGEMA_signal_5910 ), .Q ( new_AGEMA_signal_5911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C ( clk ), .D ( new_AGEMA_signal_5914 ), .Q ( new_AGEMA_signal_5915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C ( clk ), .D ( new_AGEMA_signal_5917 ), .Q ( new_AGEMA_signal_5918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C ( clk ), .D ( new_AGEMA_signal_5920 ), .Q ( new_AGEMA_signal_5921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C ( clk ), .D ( n2023 ), .Q ( new_AGEMA_signal_5923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C ( clk ), .D ( new_AGEMA_signal_1166 ), .Q ( new_AGEMA_signal_5925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C ( clk ), .D ( new_AGEMA_signal_5927 ), .Q ( new_AGEMA_signal_5928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C ( clk ), .D ( new_AGEMA_signal_5930 ), .Q ( new_AGEMA_signal_5931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C ( clk ), .D ( new_AGEMA_signal_5935 ), .Q ( new_AGEMA_signal_5936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C ( clk ), .D ( new_AGEMA_signal_5938 ), .Q ( new_AGEMA_signal_5939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C ( clk ), .D ( new_AGEMA_signal_5941 ), .Q ( new_AGEMA_signal_5942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C ( clk ), .D ( new_AGEMA_signal_5944 ), .Q ( new_AGEMA_signal_5945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C ( clk ), .D ( n2094 ), .Q ( new_AGEMA_signal_5949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C ( clk ), .D ( new_AGEMA_signal_1355 ), .Q ( new_AGEMA_signal_5951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C ( clk ), .D ( new_AGEMA_signal_5953 ), .Q ( new_AGEMA_signal_5954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C ( clk ), .D ( new_AGEMA_signal_5956 ), .Q ( new_AGEMA_signal_5957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C ( clk ), .D ( new_AGEMA_signal_5959 ), .Q ( new_AGEMA_signal_5960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C ( clk ), .D ( new_AGEMA_signal_5962 ), .Q ( new_AGEMA_signal_5963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C ( clk ), .D ( new_AGEMA_signal_5967 ), .Q ( new_AGEMA_signal_5968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C ( clk ), .D ( new_AGEMA_signal_5970 ), .Q ( new_AGEMA_signal_5971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C ( clk ), .D ( n2181 ), .Q ( new_AGEMA_signal_5975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C ( clk ), .D ( new_AGEMA_signal_1369 ), .Q ( new_AGEMA_signal_5977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C ( clk ), .D ( n2195 ), .Q ( new_AGEMA_signal_5979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C ( clk ), .D ( new_AGEMA_signal_1371 ), .Q ( new_AGEMA_signal_5981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C ( clk ), .D ( new_AGEMA_signal_5986 ), .Q ( new_AGEMA_signal_5987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C ( clk ), .D ( new_AGEMA_signal_5990 ), .Q ( new_AGEMA_signal_5991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C ( clk ), .D ( new_AGEMA_signal_5993 ), .Q ( new_AGEMA_signal_5994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C ( clk ), .D ( new_AGEMA_signal_5996 ), .Q ( new_AGEMA_signal_5997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C ( clk ), .D ( n2237 ), .Q ( new_AGEMA_signal_5999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C ( clk ), .D ( new_AGEMA_signal_1215 ), .Q ( new_AGEMA_signal_6001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C ( clk ), .D ( n2248 ), .Q ( new_AGEMA_signal_6003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C ( clk ), .D ( new_AGEMA_signal_1380 ), .Q ( new_AGEMA_signal_6005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C ( clk ), .D ( n2294 ), .Q ( new_AGEMA_signal_6011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C ( clk ), .D ( new_AGEMA_signal_1230 ), .Q ( new_AGEMA_signal_6013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C ( clk ), .D ( n2323 ), .Q ( new_AGEMA_signal_6015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C ( clk ), .D ( new_AGEMA_signal_1395 ), .Q ( new_AGEMA_signal_6017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C ( clk ), .D ( new_AGEMA_signal_6021 ), .Q ( new_AGEMA_signal_6022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C ( clk ), .D ( new_AGEMA_signal_6024 ), .Q ( new_AGEMA_signal_6025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C ( clk ), .D ( n2360 ), .Q ( new_AGEMA_signal_6027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C ( clk ), .D ( new_AGEMA_signal_1403 ), .Q ( new_AGEMA_signal_6029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C ( clk ), .D ( n2394 ), .Q ( new_AGEMA_signal_6033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C ( clk ), .D ( new_AGEMA_signal_1249 ), .Q ( new_AGEMA_signal_6035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C ( clk ), .D ( n2406 ), .Q ( new_AGEMA_signal_6037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C ( clk ), .D ( new_AGEMA_signal_1409 ), .Q ( new_AGEMA_signal_6039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C ( clk ), .D ( new_AGEMA_signal_5523 ), .Q ( new_AGEMA_signal_6041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C ( clk ), .D ( new_AGEMA_signal_5524 ), .Q ( new_AGEMA_signal_6043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C ( clk ), .D ( new_AGEMA_signal_5525 ), .Q ( new_AGEMA_signal_6047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C ( clk ), .D ( new_AGEMA_signal_5526 ), .Q ( new_AGEMA_signal_6049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C ( clk ), .D ( new_AGEMA_signal_6053 ), .Q ( new_AGEMA_signal_6054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C ( clk ), .D ( new_AGEMA_signal_6056 ), .Q ( new_AGEMA_signal_6057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C ( clk ), .D ( new_AGEMA_signal_6059 ), .Q ( new_AGEMA_signal_6060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C ( clk ), .D ( new_AGEMA_signal_6062 ), .Q ( new_AGEMA_signal_6063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C ( clk ), .D ( n2499 ), .Q ( new_AGEMA_signal_6065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C ( clk ), .D ( new_AGEMA_signal_1269 ), .Q ( new_AGEMA_signal_6067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C ( clk ), .D ( new_AGEMA_signal_6072 ), .Q ( new_AGEMA_signal_6073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C ( clk ), .D ( new_AGEMA_signal_6076 ), .Q ( new_AGEMA_signal_6077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C ( clk ), .D ( n2582 ), .Q ( new_AGEMA_signal_6081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C ( clk ), .D ( new_AGEMA_signal_1443 ), .Q ( new_AGEMA_signal_6083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C ( clk ), .D ( n2605 ), .Q ( new_AGEMA_signal_6085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C ( clk ), .D ( new_AGEMA_signal_1445 ), .Q ( new_AGEMA_signal_6087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C ( clk ), .D ( n2632 ), .Q ( new_AGEMA_signal_6089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C ( clk ), .D ( new_AGEMA_signal_1286 ), .Q ( new_AGEMA_signal_6091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C ( clk ), .D ( n2655 ), .Q ( new_AGEMA_signal_6093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C ( clk ), .D ( new_AGEMA_signal_1452 ), .Q ( new_AGEMA_signal_6095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C ( clk ), .D ( n2695 ), .Q ( new_AGEMA_signal_6097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C ( clk ), .D ( new_AGEMA_signal_1455 ), .Q ( new_AGEMA_signal_6099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C ( clk ), .D ( new_AGEMA_signal_6102 ), .Q ( new_AGEMA_signal_6103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C ( clk ), .D ( new_AGEMA_signal_6106 ), .Q ( new_AGEMA_signal_6107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C ( clk ), .D ( n2770 ), .Q ( new_AGEMA_signal_6111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C ( clk ), .D ( new_AGEMA_signal_1463 ), .Q ( new_AGEMA_signal_6113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C ( clk ), .D ( new_AGEMA_signal_6117 ), .Q ( new_AGEMA_signal_6118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C ( clk ), .D ( new_AGEMA_signal_6120 ), .Q ( new_AGEMA_signal_6121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C ( clk ), .D ( new_AGEMA_signal_6125 ), .Q ( new_AGEMA_signal_6126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C ( clk ), .D ( new_AGEMA_signal_6129 ), .Q ( new_AGEMA_signal_6130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C ( clk ), .D ( new_AGEMA_signal_6139 ), .Q ( new_AGEMA_signal_6140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C ( clk ), .D ( new_AGEMA_signal_6143 ), .Q ( new_AGEMA_signal_6144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C ( clk ), .D ( n2050 ), .Q ( new_AGEMA_signal_6149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C ( clk ), .D ( new_AGEMA_signal_1171 ), .Q ( new_AGEMA_signal_6152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C ( clk ), .D ( new_AGEMA_signal_6159 ), .Q ( new_AGEMA_signal_6160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C ( clk ), .D ( new_AGEMA_signal_6163 ), .Q ( new_AGEMA_signal_6164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C ( clk ), .D ( n2183 ), .Q ( new_AGEMA_signal_6171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C ( clk ), .D ( new_AGEMA_signal_1086 ), .Q ( new_AGEMA_signal_6174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C ( clk ), .D ( n2196 ), .Q ( new_AGEMA_signal_6177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C ( clk ), .D ( new_AGEMA_signal_1209 ), .Q ( new_AGEMA_signal_6180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C ( clk ), .D ( n2238 ), .Q ( new_AGEMA_signal_6183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C ( clk ), .D ( new_AGEMA_signal_1216 ), .Q ( new_AGEMA_signal_6186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C ( clk ), .D ( n2249 ), .Q ( new_AGEMA_signal_6189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C ( clk ), .D ( new_AGEMA_signal_1382 ), .Q ( new_AGEMA_signal_6192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C ( clk ), .D ( n2273 ), .Q ( new_AGEMA_signal_6195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C ( clk ), .D ( new_AGEMA_signal_1524 ), .Q ( new_AGEMA_signal_6198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C ( clk ), .D ( new_AGEMA_signal_6205 ), .Q ( new_AGEMA_signal_6206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C ( clk ), .D ( new_AGEMA_signal_6209 ), .Q ( new_AGEMA_signal_6210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C ( clk ), .D ( n2349 ), .Q ( new_AGEMA_signal_6217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C ( clk ), .D ( new_AGEMA_signal_1240 ), .Q ( new_AGEMA_signal_6220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C ( clk ), .D ( new_AGEMA_signal_6223 ), .Q ( new_AGEMA_signal_6224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C ( clk ), .D ( new_AGEMA_signal_6227 ), .Q ( new_AGEMA_signal_6228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C ( clk ), .D ( n2396 ), .Q ( new_AGEMA_signal_6233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C ( clk ), .D ( new_AGEMA_signal_1251 ), .Q ( new_AGEMA_signal_6236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C ( clk ), .D ( n2439 ), .Q ( new_AGEMA_signal_6243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C ( clk ), .D ( new_AGEMA_signal_1417 ), .Q ( new_AGEMA_signal_6246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C ( clk ), .D ( n2470 ), .Q ( new_AGEMA_signal_6249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C ( clk ), .D ( new_AGEMA_signal_1261 ), .Q ( new_AGEMA_signal_6252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C ( clk ), .D ( new_AGEMA_signal_6255 ), .Q ( new_AGEMA_signal_6256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C ( clk ), .D ( new_AGEMA_signal_6259 ), .Q ( new_AGEMA_signal_6260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C ( clk ), .D ( new_AGEMA_signal_6263 ), .Q ( new_AGEMA_signal_6264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C ( clk ), .D ( new_AGEMA_signal_6267 ), .Q ( new_AGEMA_signal_6268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C ( clk ), .D ( n2585 ), .Q ( new_AGEMA_signal_6271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C ( clk ), .D ( new_AGEMA_signal_1441 ), .Q ( new_AGEMA_signal_6274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C ( clk ), .D ( n2607 ), .Q ( new_AGEMA_signal_6277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C ( clk ), .D ( new_AGEMA_signal_1279 ), .Q ( new_AGEMA_signal_6280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C ( clk ), .D ( n2013 ), .Q ( new_AGEMA_signal_6311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C ( clk ), .D ( new_AGEMA_signal_1335 ), .Q ( new_AGEMA_signal_6315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C ( clk ), .D ( n2028 ), .Q ( new_AGEMA_signal_6319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C ( clk ), .D ( new_AGEMA_signal_1071 ), .Q ( new_AGEMA_signal_6323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C ( clk ), .D ( n2051 ), .Q ( new_AGEMA_signal_6327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C ( clk ), .D ( new_AGEMA_signal_1341 ), .Q ( new_AGEMA_signal_6331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C ( clk ), .D ( n2069 ), .Q ( new_AGEMA_signal_6335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C ( clk ), .D ( new_AGEMA_signal_1346 ), .Q ( new_AGEMA_signal_6339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C ( clk ), .D ( new_AGEMA_signal_6349 ), .Q ( new_AGEMA_signal_6350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C ( clk ), .D ( new_AGEMA_signal_6354 ), .Q ( new_AGEMA_signal_6355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C ( clk ), .D ( n2144 ), .Q ( new_AGEMA_signal_6359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C ( clk ), .D ( new_AGEMA_signal_1363 ), .Q ( new_AGEMA_signal_6363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C ( clk ), .D ( n2170 ), .Q ( new_AGEMA_signal_6367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C ( clk ), .D ( new_AGEMA_signal_1365 ), .Q ( new_AGEMA_signal_6371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C ( clk ), .D ( n2186 ), .Q ( new_AGEMA_signal_6375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_6379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C ( clk ), .D ( new_AGEMA_signal_6399 ), .Q ( new_AGEMA_signal_6400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C ( clk ), .D ( new_AGEMA_signal_6404 ), .Q ( new_AGEMA_signal_6405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C ( clk ), .D ( new_AGEMA_signal_5653 ), .Q ( new_AGEMA_signal_6409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C ( clk ), .D ( new_AGEMA_signal_5654 ), .Q ( new_AGEMA_signal_6413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C ( clk ), .D ( n2551 ), .Q ( new_AGEMA_signal_6423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C ( clk ), .D ( new_AGEMA_signal_1435 ), .Q ( new_AGEMA_signal_6427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C ( clk ), .D ( n2588 ), .Q ( new_AGEMA_signal_6431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C ( clk ), .D ( new_AGEMA_signal_1444 ), .Q ( new_AGEMA_signal_6435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C ( clk ), .D ( n2701 ), .Q ( new_AGEMA_signal_6449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C ( clk ), .D ( new_AGEMA_signal_1293 ), .Q ( new_AGEMA_signal_6453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C ( clk ), .D ( n2172 ), .Q ( new_AGEMA_signal_6515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C ( clk ), .D ( new_AGEMA_signal_1368 ), .Q ( new_AGEMA_signal_6520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C ( clk ), .D ( n2150 ), .Q ( new_AGEMA_signal_6711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C ( clk ), .D ( new_AGEMA_signal_1197 ), .Q ( new_AGEMA_signal_6718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C ( clk ), .D ( n2369 ), .Q ( new_AGEMA_signal_6733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C ( clk ), .D ( new_AGEMA_signal_1540 ), .Q ( new_AGEMA_signal_6740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C ( clk ), .D ( n2152 ), .Q ( new_AGEMA_signal_6769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C ( clk ), .D ( new_AGEMA_signal_1364 ), .Q ( new_AGEMA_signal_6777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C ( clk ), .D ( n2372 ), .Q ( new_AGEMA_signal_6791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C ( clk ), .D ( new_AGEMA_signal_1404 ), .Q ( new_AGEMA_signal_6799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C ( clk ), .D ( n2375 ), .Q ( new_AGEMA_signal_6867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C ( clk ), .D ( new_AGEMA_signal_1241 ), .Q ( new_AGEMA_signal_6876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C ( clk ), .D ( n2377 ), .Q ( new_AGEMA_signal_6917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C ( clk ), .D ( new_AGEMA_signal_1405 ), .Q ( new_AGEMA_signal_6927 ) ) ;

    /* cells in depth 5 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1983 ( .a ({new_AGEMA_signal_5692, new_AGEMA_signal_5690}), .b ({new_AGEMA_signal_1471, n1928}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300]}), .c ({new_AGEMA_signal_1585, n1934}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U1998 ( .a ({new_AGEMA_signal_1472, n1931}), .b ({new_AGEMA_signal_5696, new_AGEMA_signal_5694}), .clk ( clk ), .r ({Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_1586, n1932}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2015 ( .a ({new_AGEMA_signal_1473, n1939}), .b ({new_AGEMA_signal_5698, new_AGEMA_signal_5697}), .clk ( clk ), .r ({Fresh[2311], Fresh[2310], Fresh[2309], Fresh[2308]}), .c ({new_AGEMA_signal_1587, n1940}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2033 ( .a ({new_AGEMA_signal_1474, n1948}), .b ({new_AGEMA_signal_1475, n1947}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312]}), .c ({new_AGEMA_signal_1588, n1961}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2050 ( .a ({new_AGEMA_signal_1476, n1954}), .b ({new_AGEMA_signal_1477, n1953}), .clk ( clk ), .r ({Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_1589, n1955}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2066 ( .a ({new_AGEMA_signal_5700, new_AGEMA_signal_5699}), .b ({new_AGEMA_signal_1322, n1965}), .clk ( clk ), .r ({Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320]}), .c ({new_AGEMA_signal_1479, n1967}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2085 ( .a ({new_AGEMA_signal_1591, n1970}), .b ({new_AGEMA_signal_1481, n1969}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324]}), .c ({new_AGEMA_signal_1669, n1984}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2103 ( .a ({new_AGEMA_signal_5704, new_AGEMA_signal_5702}), .b ({new_AGEMA_signal_1483, n1975}), .clk ( clk ), .r ({Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_1592, n1977}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2108 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705}), .b ({new_AGEMA_signal_1484, n1980}), .clk ( clk ), .r ({Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332]}), .c ({new_AGEMA_signal_1593, n1981}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2115 ( .a ({new_AGEMA_signal_5710, new_AGEMA_signal_5708}), .b ({new_AGEMA_signal_1329, n1986}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336]}), .c ({new_AGEMA_signal_1485, n1987}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2127 ( .a ({new_AGEMA_signal_1486, n1997}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711}), .clk ( clk ), .r ({Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_1594, n1998}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2146 ( .a ({new_AGEMA_signal_5716, new_AGEMA_signal_5714}), .b ({new_AGEMA_signal_1488, n2007}), .clk ( clk ), .r ({Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344]}), .c ({new_AGEMA_signal_1595, n2010}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2162 ( .a ({new_AGEMA_signal_5720, new_AGEMA_signal_5718}), .b ({new_AGEMA_signal_1336, n2021}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348]}), .c ({new_AGEMA_signal_1489, n2024}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2177 ( .a ({new_AGEMA_signal_5722, new_AGEMA_signal_5721}), .b ({new_AGEMA_signal_1490, n2032}), .clk ( clk ), .r ({Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_1597, n2035}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2186 ( .a ({new_AGEMA_signal_1491, n2041}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723}), .clk ( clk ), .r ({Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356]}), .c ({new_AGEMA_signal_1598, n2054}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2190 ( .a ({new_AGEMA_signal_5726, new_AGEMA_signal_5725}), .b ({new_AGEMA_signal_1492, n2043}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360]}), .c ({new_AGEMA_signal_1599, n2048}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2195 ( .a ({new_AGEMA_signal_1493, n2046}), .b ({new_AGEMA_signal_5728, new_AGEMA_signal_5727}), .clk ( clk ), .r ({Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_1600, n2047}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2206 ( .a ({new_AGEMA_signal_1494, n2058}), .b ({new_AGEMA_signal_5732, new_AGEMA_signal_5730}), .clk ( clk ), .r ({Fresh[2371], Fresh[2370], Fresh[2369], Fresh[2368]}), .c ({new_AGEMA_signal_1601, n2059}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2213 ( .a ({new_AGEMA_signal_1495, n2063}), .b ({new_AGEMA_signal_5736, new_AGEMA_signal_5734}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372]}), .c ({new_AGEMA_signal_1602, n2064}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2229 ( .a ({new_AGEMA_signal_1497, n2076}), .b ({new_AGEMA_signal_5740, new_AGEMA_signal_5738}), .clk ( clk ), .r ({Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_1603, n2077}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2249 ( .a ({new_AGEMA_signal_1501, n2090}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741}), .clk ( clk ), .r ({Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380]}), .c ({new_AGEMA_signal_1604, n2158}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2255 ( .a ({new_AGEMA_signal_1502, n2093}), .b ({new_AGEMA_signal_5744, new_AGEMA_signal_5743}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384]}), .c ({new_AGEMA_signal_1605, n2095}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2274 ( .a ({new_AGEMA_signal_1606, n2116}), .b ({new_AGEMA_signal_5746, new_AGEMA_signal_5745}), .clk ( clk ), .r ({Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_1681, n2117}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2283 ( .a ({new_AGEMA_signal_5750, new_AGEMA_signal_5748}), .b ({new_AGEMA_signal_1505, n2120}), .clk ( clk ), .r ({Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392]}), .c ({new_AGEMA_signal_1607, n2123}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2300 ( .a ({new_AGEMA_signal_5752, new_AGEMA_signal_5751}), .b ({new_AGEMA_signal_1360, n2134}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396]}), .c ({new_AGEMA_signal_1507, n2135}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2309 ( .a ({new_AGEMA_signal_5756, new_AGEMA_signal_5754}), .b ({new_AGEMA_signal_1509, n2140}), .clk ( clk ), .r ({Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_1609, n2141}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2327 ( .a ({new_AGEMA_signal_5762, new_AGEMA_signal_5759}), .b ({new_AGEMA_signal_1511, n2161}), .clk ( clk ), .r ({Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404]}), .c ({new_AGEMA_signal_1610, n2166}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2331 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5764}), .b ({new_AGEMA_signal_1367, n2164}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408]}), .c ({new_AGEMA_signal_1512, n2165}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2346 ( .a ({new_AGEMA_signal_1513, n2179}), .b ({new_AGEMA_signal_5770, new_AGEMA_signal_5768}), .clk ( clk ), .r ({Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_1611, n2180}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2360 ( .a ({new_AGEMA_signal_5772, new_AGEMA_signal_5771}), .b ({new_AGEMA_signal_1514, n2192}), .clk ( clk ), .r ({Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416]}), .c ({new_AGEMA_signal_1612, n2194}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2372 ( .a ({new_AGEMA_signal_1613, n2203}), .b ({new_AGEMA_signal_5774, new_AGEMA_signal_5773}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420]}), .c ({new_AGEMA_signal_1688, n2204}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2389 ( .a ({new_AGEMA_signal_1517, n2224}), .b ({new_AGEMA_signal_1518, n2223}), .clk ( clk ), .r ({Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_1614, n2225}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2394 ( .a ({new_AGEMA_signal_1379, n2229}), .b ({new_AGEMA_signal_5776, new_AGEMA_signal_5775}), .clk ( clk ), .r ({Fresh[2431], Fresh[2430], Fresh[2429], Fresh[2428]}), .c ({new_AGEMA_signal_1519, n2230}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2400 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777}), .b ({new_AGEMA_signal_1616, n2234}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432]}), .c ({new_AGEMA_signal_1690, n2236}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2412 ( .a ({new_AGEMA_signal_1521, n2246}), .b ({new_AGEMA_signal_5782, new_AGEMA_signal_5780}), .clk ( clk ), .r ({Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_1617, n2247}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2419 ( .a ({new_AGEMA_signal_1522, n2254}), .b ({new_AGEMA_signal_5788, new_AGEMA_signal_5785}), .clk ( clk ), .r ({Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440]}), .c ({new_AGEMA_signal_1618, n2255}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2427 ( .a ({new_AGEMA_signal_1523, n2263}), .b ({new_AGEMA_signal_5792, new_AGEMA_signal_5790}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444]}), .c ({new_AGEMA_signal_1619, n2264}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2435 ( .a ({new_AGEMA_signal_5794, new_AGEMA_signal_5793}), .b ({new_AGEMA_signal_1385, n2267}), .clk ( clk ), .r ({Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_1620, n2271}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2446 ( .a ({new_AGEMA_signal_5710, new_AGEMA_signal_5708}), .b ({new_AGEMA_signal_1387, n2279}), .clk ( clk ), .r ({Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452]}), .c ({new_AGEMA_signal_1526, n2280}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2451 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795}), .b ({new_AGEMA_signal_1388, n2283}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456]}), .c ({new_AGEMA_signal_1527, n2286}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2461 ( .a ({new_AGEMA_signal_1529, n2686}), .b ({new_AGEMA_signal_1530, n2289}), .clk ( clk ), .r ({Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_1622, n2304}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2466 ( .a ({new_AGEMA_signal_5798, new_AGEMA_signal_5797}), .b ({new_AGEMA_signal_1532, n2292}), .clk ( clk ), .r ({Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464]}), .c ({new_AGEMA_signal_1623, n2295}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2488 ( .a ({new_AGEMA_signal_1534, n2321}), .b ({new_AGEMA_signal_1233, n2320}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468]}), .c ({new_AGEMA_signal_1624, n2322}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2499 ( .a ({new_AGEMA_signal_1535, n2332}), .b ({new_AGEMA_signal_1536, n2331}), .clk ( clk ), .r ({Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_1625, n2333}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2509 ( .a ({new_AGEMA_signal_5802, new_AGEMA_signal_5800}), .b ({new_AGEMA_signal_1538, n2342}), .clk ( clk ), .r ({Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476]}), .c ({new_AGEMA_signal_1627, n2345}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2526 ( .a ({new_AGEMA_signal_1539, n2358}), .b ({new_AGEMA_signal_5804, new_AGEMA_signal_5803}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480]}), .c ({new_AGEMA_signal_1628, n2361}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2549 ( .a ({new_AGEMA_signal_1406, n2387}), .b ({new_AGEMA_signal_5806, new_AGEMA_signal_5805}), .clk ( clk ), .r ({Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_1541, n2388}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2556 ( .a ({new_AGEMA_signal_5810, new_AGEMA_signal_5808}), .b ({new_AGEMA_signal_1542, n2392}), .clk ( clk ), .r ({Fresh[2491], Fresh[2490], Fresh[2489], Fresh[2488]}), .c ({new_AGEMA_signal_1630, n2393}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2567 ( .a ({new_AGEMA_signal_5814, new_AGEMA_signal_5812}), .b ({new_AGEMA_signal_1410, n2404}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492]}), .c ({new_AGEMA_signal_1543, n2405}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2571 ( .a ({new_AGEMA_signal_1544, n2409}), .b ({new_AGEMA_signal_5818, new_AGEMA_signal_5816}), .clk ( clk ), .r ({Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_1632, n2410}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2576 ( .a ({new_AGEMA_signal_5822, new_AGEMA_signal_5820}), .b ({new_AGEMA_signal_1545, n2414}), .clk ( clk ), .r ({Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500]}), .c ({new_AGEMA_signal_1633, n2421}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2579 ( .a ({new_AGEMA_signal_1413, n2418}), .b ({new_AGEMA_signal_5826, new_AGEMA_signal_5824}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504]}), .c ({new_AGEMA_signal_1546, n2419}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2590 ( .a ({new_AGEMA_signal_5828, new_AGEMA_signal_5827}), .b ({new_AGEMA_signal_1547, n2432}), .clk ( clk ), .r ({Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_1635, n2436}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2604 ( .a ({new_AGEMA_signal_1548, n2449}), .b ({new_AGEMA_signal_1549, n2448}), .clk ( clk ), .r ({Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512]}), .c ({new_AGEMA_signal_1636, n2450}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2610 ( .a ({new_AGEMA_signal_5830, new_AGEMA_signal_5829}), .b ({new_AGEMA_signal_1550, n2455}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516]}), .c ({new_AGEMA_signal_1637, n2456}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2613 ( .a ({new_AGEMA_signal_1551, n2460}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831}), .clk ( clk ), .r ({Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_1638, n2461}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2619 ( .a ({new_AGEMA_signal_5834, new_AGEMA_signal_5833}), .b ({new_AGEMA_signal_1422, n2466}), .clk ( clk ), .r ({Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524]}), .c ({new_AGEMA_signal_1552, n2469}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2630 ( .a ({new_AGEMA_signal_5838, new_AGEMA_signal_5836}), .b ({new_AGEMA_signal_1423, n2477}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528]}), .c ({new_AGEMA_signal_1553, n2478}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2635 ( .a ({new_AGEMA_signal_5842, new_AGEMA_signal_5840}), .b ({new_AGEMA_signal_1554, n2482}), .clk ( clk ), .r ({Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_1640, n2484}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2643 ( .a ({new_AGEMA_signal_1425, n2490}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843}), .clk ( clk ), .r ({Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536]}), .c ({new_AGEMA_signal_1555, n2491}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2649 ( .a ({new_AGEMA_signal_5846, new_AGEMA_signal_5845}), .b ({new_AGEMA_signal_1556, n2496}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540]}), .c ({new_AGEMA_signal_1642, n2500}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2656 ( .a ({new_AGEMA_signal_1643, n2507}), .b ({new_AGEMA_signal_5848, new_AGEMA_signal_5847}), .clk ( clk ), .r ({Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_1708, n2508}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2670 ( .a ({new_AGEMA_signal_1644, n2525}), .b ({new_AGEMA_signal_1559, n2524}), .clk ( clk ), .r ({Fresh[2551], Fresh[2550], Fresh[2549], Fresh[2548]}), .c ({new_AGEMA_signal_1709, n2526}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2679 ( .a ({new_AGEMA_signal_1560, n2537}), .b ({new_AGEMA_signal_1561, n2536}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552]}), .c ({new_AGEMA_signal_1645, n2539}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2682 ( .a ({new_AGEMA_signal_1506, n2543}), .b ({new_AGEMA_signal_5850, new_AGEMA_signal_5849}), .clk ( clk ), .r ({Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_1646, n2548}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2694 ( .a ({new_AGEMA_signal_5852, new_AGEMA_signal_5851}), .b ({new_AGEMA_signal_1562, n2557}), .clk ( clk ), .r ({Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560]}), .c ({new_AGEMA_signal_1647, n2568}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2700 ( .a ({new_AGEMA_signal_5854, new_AGEMA_signal_5853}), .b ({new_AGEMA_signal_1563, n2565}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564]}), .c ({new_AGEMA_signal_1648, n2567}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2710 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855}), .b ({new_AGEMA_signal_1565, n2580}), .clk ( clk ), .r ({Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_1649, n2583}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2728 ( .a ({new_AGEMA_signal_5858, new_AGEMA_signal_5857}), .b ({new_AGEMA_signal_1282, n2602}), .clk ( clk ), .r ({Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572]}), .c ({new_AGEMA_signal_1566, n2604}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2739 ( .a ({new_AGEMA_signal_5860, new_AGEMA_signal_5859}), .b ({new_AGEMA_signal_1567, n2619}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576]}), .c ({new_AGEMA_signal_1651, n2621}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2745 ( .a ({new_AGEMA_signal_5864, new_AGEMA_signal_5862}), .b ({new_AGEMA_signal_1568, n2628}), .clk ( clk ), .r ({Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_1652, n2633}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2756 ( .a ({new_AGEMA_signal_1569, n2649}), .b ({new_AGEMA_signal_1451, n2648}), .clk ( clk ), .r ({Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584]}), .c ({new_AGEMA_signal_1653, n2660}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2759 ( .a ({new_AGEMA_signal_5866, new_AGEMA_signal_5865}), .b ({new_AGEMA_signal_1496, n2652}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588]}), .c ({new_AGEMA_signal_1654, n2656}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2766 ( .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867}), .b ({new_AGEMA_signal_1570, n2664}), .clk ( clk ), .r ({Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_1655, n2666}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2774 ( .a ({new_AGEMA_signal_1571, n2681}), .b ({new_AGEMA_signal_1454, n2680}), .clk ( clk ), .r ({Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596]}), .c ({new_AGEMA_signal_1656, n2706}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2777 ( .a ({new_AGEMA_signal_1529, n2686}), .b ({new_AGEMA_signal_1572, n2685}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600]}), .c ({new_AGEMA_signal_1657, n2704}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2781 ( .a ({new_AGEMA_signal_1574, n2692}), .b ({new_AGEMA_signal_5870, new_AGEMA_signal_5869}), .clk ( clk ), .r ({Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_1658, n2696}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2794 ( .a ({new_AGEMA_signal_5872, new_AGEMA_signal_5871}), .b ({new_AGEMA_signal_1575, n2716}), .clk ( clk ), .r ({Fresh[2611], Fresh[2610], Fresh[2609], Fresh[2608]}), .c ({new_AGEMA_signal_1659, n2718}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2801 ( .a ({new_AGEMA_signal_5874, new_AGEMA_signal_5873}), .b ({new_AGEMA_signal_1457, n2728}), .clk ( clk ), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612]}), .c ({new_AGEMA_signal_1660, n2730}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2805 ( .a ({new_AGEMA_signal_5878, new_AGEMA_signal_5876}), .b ({new_AGEMA_signal_1577, n2735}), .clk ( clk ), .r ({Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_1661, n2745}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2809 ( .a ({new_AGEMA_signal_1578, n2743}), .b ({new_AGEMA_signal_5882, new_AGEMA_signal_5880}), .clk ( clk ), .r ({Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620]}), .c ({new_AGEMA_signal_1662, n2744}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2814 ( .a ({new_AGEMA_signal_5794, new_AGEMA_signal_5793}), .b ({new_AGEMA_signal_1460, n2751}), .clk ( clk ), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624]}), .c ({new_AGEMA_signal_1663, n2759}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2821 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5884}), .b ({new_AGEMA_signal_1580, n2764}), .clk ( clk ), .r ({Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_1664, n2771}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2833 ( .a ({new_AGEMA_signal_1466, n2788}), .b ({new_AGEMA_signal_5890, new_AGEMA_signal_5888}), .clk ( clk ), .r ({Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632]}), .c ({new_AGEMA_signal_1582, n2798}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2850 ( .a ({new_AGEMA_signal_1584, n2822}), .b ({new_AGEMA_signal_1469, n2821}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636]}), .c ({new_AGEMA_signal_1666, n2826}) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C ( clk ), .D ( new_AGEMA_signal_5891 ), .Q ( new_AGEMA_signal_5892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C ( clk ), .D ( new_AGEMA_signal_5893 ), .Q ( new_AGEMA_signal_5894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C ( clk ), .D ( new_AGEMA_signal_5895 ), .Q ( new_AGEMA_signal_5896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C ( clk ), .D ( new_AGEMA_signal_5897 ), .Q ( new_AGEMA_signal_5898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C ( clk ), .D ( new_AGEMA_signal_5901 ), .Q ( new_AGEMA_signal_5902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C ( clk ), .D ( new_AGEMA_signal_5905 ), .Q ( new_AGEMA_signal_5906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C ( clk ), .D ( n1978 ), .Q ( new_AGEMA_signal_5907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C ( clk ), .D ( new_AGEMA_signal_1482 ), .Q ( new_AGEMA_signal_5908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C ( clk ), .D ( new_AGEMA_signal_5911 ), .Q ( new_AGEMA_signal_5912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C ( clk ), .D ( new_AGEMA_signal_5915 ), .Q ( new_AGEMA_signal_5916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C ( clk ), .D ( new_AGEMA_signal_5918 ), .Q ( new_AGEMA_signal_5919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C ( clk ), .D ( new_AGEMA_signal_5921 ), .Q ( new_AGEMA_signal_5922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C ( clk ), .D ( new_AGEMA_signal_5923 ), .Q ( new_AGEMA_signal_5924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C ( clk ), .D ( new_AGEMA_signal_5925 ), .Q ( new_AGEMA_signal_5926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C ( clk ), .D ( new_AGEMA_signal_5928 ), .Q ( new_AGEMA_signal_5929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C ( clk ), .D ( new_AGEMA_signal_5931 ), .Q ( new_AGEMA_signal_5932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C ( clk ), .D ( new_AGEMA_signal_5836 ), .Q ( new_AGEMA_signal_5933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C ( clk ), .D ( new_AGEMA_signal_5838 ), .Q ( new_AGEMA_signal_5934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C ( clk ), .D ( new_AGEMA_signal_5936 ), .Q ( new_AGEMA_signal_5937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C ( clk ), .D ( new_AGEMA_signal_5939 ), .Q ( new_AGEMA_signal_5940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C ( clk ), .D ( new_AGEMA_signal_5942 ), .Q ( new_AGEMA_signal_5943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C ( clk ), .D ( new_AGEMA_signal_5945 ), .Q ( new_AGEMA_signal_5946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C ( clk ), .D ( n2091 ), .Q ( new_AGEMA_signal_5947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C ( clk ), .D ( new_AGEMA_signal_1500 ), .Q ( new_AGEMA_signal_5948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C ( clk ), .D ( new_AGEMA_signal_5949 ), .Q ( new_AGEMA_signal_5950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C ( clk ), .D ( new_AGEMA_signal_5951 ), .Q ( new_AGEMA_signal_5952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C ( clk ), .D ( new_AGEMA_signal_5954 ), .Q ( new_AGEMA_signal_5955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C ( clk ), .D ( new_AGEMA_signal_5957 ), .Q ( new_AGEMA_signal_5958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C ( clk ), .D ( new_AGEMA_signal_5960 ), .Q ( new_AGEMA_signal_5961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C ( clk ), .D ( new_AGEMA_signal_5963 ), .Q ( new_AGEMA_signal_5964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C ( clk ), .D ( n2543 ), .Q ( new_AGEMA_signal_5965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C ( clk ), .D ( new_AGEMA_signal_1506 ), .Q ( new_AGEMA_signal_5966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C ( clk ), .D ( new_AGEMA_signal_5968 ), .Q ( new_AGEMA_signal_5969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C ( clk ), .D ( new_AGEMA_signal_5971 ), .Q ( new_AGEMA_signal_5972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C ( clk ), .D ( n2159 ), .Q ( new_AGEMA_signal_5973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C ( clk ), .D ( new_AGEMA_signal_1510 ), .Q ( new_AGEMA_signal_5974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C ( clk ), .D ( new_AGEMA_signal_5975 ), .Q ( new_AGEMA_signal_5976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C ( clk ), .D ( new_AGEMA_signal_5977 ), .Q ( new_AGEMA_signal_5978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C ( clk ), .D ( new_AGEMA_signal_5979 ), .Q ( new_AGEMA_signal_5980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C ( clk ), .D ( new_AGEMA_signal_5981 ), .Q ( new_AGEMA_signal_5982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C ( clk ), .D ( new_AGEMA_signal_5829 ), .Q ( new_AGEMA_signal_5983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C ( clk ), .D ( new_AGEMA_signal_5830 ), .Q ( new_AGEMA_signal_5984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C ( clk ), .D ( new_AGEMA_signal_5987 ), .Q ( new_AGEMA_signal_5988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C ( clk ), .D ( new_AGEMA_signal_5991 ), .Q ( new_AGEMA_signal_5992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C ( clk ), .D ( new_AGEMA_signal_5994 ), .Q ( new_AGEMA_signal_5995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C ( clk ), .D ( new_AGEMA_signal_5997 ), .Q ( new_AGEMA_signal_5998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C ( clk ), .D ( new_AGEMA_signal_5999 ), .Q ( new_AGEMA_signal_6000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C ( clk ), .D ( new_AGEMA_signal_6001 ), .Q ( new_AGEMA_signal_6002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C ( clk ), .D ( new_AGEMA_signal_6003 ), .Q ( new_AGEMA_signal_6004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C ( clk ), .D ( new_AGEMA_signal_6005 ), .Q ( new_AGEMA_signal_6006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C ( clk ), .D ( n2270 ), .Q ( new_AGEMA_signal_6007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C ( clk ), .D ( new_AGEMA_signal_1386 ), .Q ( new_AGEMA_signal_6008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C ( clk ), .D ( n2285 ), .Q ( new_AGEMA_signal_6009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C ( clk ), .D ( new_AGEMA_signal_1528 ), .Q ( new_AGEMA_signal_6010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C ( clk ), .D ( new_AGEMA_signal_6011 ), .Q ( new_AGEMA_signal_6012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C ( clk ), .D ( new_AGEMA_signal_6013 ), .Q ( new_AGEMA_signal_6014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C ( clk ), .D ( new_AGEMA_signal_6015 ), .Q ( new_AGEMA_signal_6016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C ( clk ), .D ( new_AGEMA_signal_6017 ), .Q ( new_AGEMA_signal_6018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C ( clk ), .D ( n2334 ), .Q ( new_AGEMA_signal_6019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C ( clk ), .D ( new_AGEMA_signal_1397 ), .Q ( new_AGEMA_signal_6020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C ( clk ), .D ( new_AGEMA_signal_6022 ), .Q ( new_AGEMA_signal_6023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C ( clk ), .D ( new_AGEMA_signal_6025 ), .Q ( new_AGEMA_signal_6026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C ( clk ), .D ( new_AGEMA_signal_6027 ), .Q ( new_AGEMA_signal_6028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C ( clk ), .D ( new_AGEMA_signal_6029 ), .Q ( new_AGEMA_signal_6030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C ( clk ), .D ( new_AGEMA_signal_5833 ), .Q ( new_AGEMA_signal_6031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C ( clk ), .D ( new_AGEMA_signal_5834 ), .Q ( new_AGEMA_signal_6032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C ( clk ), .D ( new_AGEMA_signal_6033 ), .Q ( new_AGEMA_signal_6034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C ( clk ), .D ( new_AGEMA_signal_6035 ), .Q ( new_AGEMA_signal_6036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C ( clk ), .D ( new_AGEMA_signal_6037 ), .Q ( new_AGEMA_signal_6038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C ( clk ), .D ( new_AGEMA_signal_6039 ), .Q ( new_AGEMA_signal_6040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C ( clk ), .D ( new_AGEMA_signal_6041 ), .Q ( new_AGEMA_signal_6042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C ( clk ), .D ( new_AGEMA_signal_6043 ), .Q ( new_AGEMA_signal_6044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C ( clk ), .D ( n2435 ), .Q ( new_AGEMA_signal_6045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C ( clk ), .D ( new_AGEMA_signal_1416 ), .Q ( new_AGEMA_signal_6046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C ( clk ), .D ( new_AGEMA_signal_6047 ), .Q ( new_AGEMA_signal_6048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C ( clk ), .D ( new_AGEMA_signal_6049 ), .Q ( new_AGEMA_signal_6050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C ( clk ), .D ( new_AGEMA_signal_5795 ), .Q ( new_AGEMA_signal_6051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C ( clk ), .D ( new_AGEMA_signal_5796 ), .Q ( new_AGEMA_signal_6052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C ( clk ), .D ( new_AGEMA_signal_6054 ), .Q ( new_AGEMA_signal_6055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C ( clk ), .D ( new_AGEMA_signal_6057 ), .Q ( new_AGEMA_signal_6058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C ( clk ), .D ( new_AGEMA_signal_6060 ), .Q ( new_AGEMA_signal_6061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C ( clk ), .D ( new_AGEMA_signal_6063 ), .Q ( new_AGEMA_signal_6064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C ( clk ), .D ( new_AGEMA_signal_6065 ), .Q ( new_AGEMA_signal_6066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C ( clk ), .D ( new_AGEMA_signal_6067 ), .Q ( new_AGEMA_signal_6068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C ( clk ), .D ( new_AGEMA_signal_5785 ), .Q ( new_AGEMA_signal_6069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C ( clk ), .D ( new_AGEMA_signal_5788 ), .Q ( new_AGEMA_signal_6070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C ( clk ), .D ( new_AGEMA_signal_6073 ), .Q ( new_AGEMA_signal_6074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C ( clk ), .D ( new_AGEMA_signal_6077 ), .Q ( new_AGEMA_signal_6078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C ( clk ), .D ( n2547 ), .Q ( new_AGEMA_signal_6079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C ( clk ), .D ( new_AGEMA_signal_1434 ), .Q ( new_AGEMA_signal_6080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C ( clk ), .D ( new_AGEMA_signal_6081 ), .Q ( new_AGEMA_signal_6082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C ( clk ), .D ( new_AGEMA_signal_6083 ), .Q ( new_AGEMA_signal_6084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C ( clk ), .D ( new_AGEMA_signal_6085 ), .Q ( new_AGEMA_signal_6086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C ( clk ), .D ( new_AGEMA_signal_6087 ), .Q ( new_AGEMA_signal_6088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C ( clk ), .D ( new_AGEMA_signal_6089 ), .Q ( new_AGEMA_signal_6090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C ( clk ), .D ( new_AGEMA_signal_6091 ), .Q ( new_AGEMA_signal_6092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C ( clk ), .D ( new_AGEMA_signal_6093 ), .Q ( new_AGEMA_signal_6094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C ( clk ), .D ( new_AGEMA_signal_6095 ), .Q ( new_AGEMA_signal_6096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C ( clk ), .D ( new_AGEMA_signal_6097 ), .Q ( new_AGEMA_signal_6098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C ( clk ), .D ( new_AGEMA_signal_6099 ), .Q ( new_AGEMA_signal_6100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C ( clk ), .D ( new_AGEMA_signal_6103 ), .Q ( new_AGEMA_signal_6104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C ( clk ), .D ( new_AGEMA_signal_6107 ), .Q ( new_AGEMA_signal_6108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C ( clk ), .D ( n2758 ), .Q ( new_AGEMA_signal_6109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C ( clk ), .D ( new_AGEMA_signal_1579 ), .Q ( new_AGEMA_signal_6110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C ( clk ), .D ( new_AGEMA_signal_6111 ), .Q ( new_AGEMA_signal_6112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C ( clk ), .D ( new_AGEMA_signal_6113 ), .Q ( new_AGEMA_signal_6114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C ( clk ), .D ( n2797 ), .Q ( new_AGEMA_signal_6115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C ( clk ), .D ( new_AGEMA_signal_1583 ), .Q ( new_AGEMA_signal_6116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C ( clk ), .D ( new_AGEMA_signal_6118 ), .Q ( new_AGEMA_signal_6119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C ( clk ), .D ( new_AGEMA_signal_6121 ), .Q ( new_AGEMA_signal_6122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C ( clk ), .D ( new_AGEMA_signal_6126 ), .Q ( new_AGEMA_signal_6127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C ( clk ), .D ( new_AGEMA_signal_6130 ), .Q ( new_AGEMA_signal_6131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C ( clk ), .D ( n2012 ), .Q ( new_AGEMA_signal_6135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C ( clk ), .D ( new_AGEMA_signal_1487 ), .Q ( new_AGEMA_signal_6137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C ( clk ), .D ( new_AGEMA_signal_6140 ), .Q ( new_AGEMA_signal_6141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C ( clk ), .D ( new_AGEMA_signal_6144 ), .Q ( new_AGEMA_signal_6145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C ( clk ), .D ( new_AGEMA_signal_6149 ), .Q ( new_AGEMA_signal_6150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C ( clk ), .D ( new_AGEMA_signal_6152 ), .Q ( new_AGEMA_signal_6153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C ( clk ), .D ( n2652 ), .Q ( new_AGEMA_signal_6155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C ( clk ), .D ( new_AGEMA_signal_1496 ), .Q ( new_AGEMA_signal_6157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C ( clk ), .D ( new_AGEMA_signal_6160 ), .Q ( new_AGEMA_signal_6161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C ( clk ), .D ( new_AGEMA_signal_6164 ), .Q ( new_AGEMA_signal_6165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C ( clk ), .D ( n2143 ), .Q ( new_AGEMA_signal_6167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C ( clk ), .D ( new_AGEMA_signal_1508 ), .Q ( new_AGEMA_signal_6169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C ( clk ), .D ( new_AGEMA_signal_6171 ), .Q ( new_AGEMA_signal_6172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C ( clk ), .D ( new_AGEMA_signal_6174 ), .Q ( new_AGEMA_signal_6175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C ( clk ), .D ( new_AGEMA_signal_6177 ), .Q ( new_AGEMA_signal_6178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C ( clk ), .D ( new_AGEMA_signal_6180 ), .Q ( new_AGEMA_signal_6181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C ( clk ), .D ( new_AGEMA_signal_6183 ), .Q ( new_AGEMA_signal_6184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C ( clk ), .D ( new_AGEMA_signal_6186 ), .Q ( new_AGEMA_signal_6187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C ( clk ), .D ( new_AGEMA_signal_6189 ), .Q ( new_AGEMA_signal_6190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C ( clk ), .D ( new_AGEMA_signal_6192 ), .Q ( new_AGEMA_signal_6193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C ( clk ), .D ( new_AGEMA_signal_6195 ), .Q ( new_AGEMA_signal_6196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C ( clk ), .D ( new_AGEMA_signal_6198 ), .Q ( new_AGEMA_signal_6199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C ( clk ), .D ( n2297 ), .Q ( new_AGEMA_signal_6201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C ( clk ), .D ( new_AGEMA_signal_1531 ), .Q ( new_AGEMA_signal_6203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C ( clk ), .D ( new_AGEMA_signal_6206 ), .Q ( new_AGEMA_signal_6207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C ( clk ), .D ( new_AGEMA_signal_6210 ), .Q ( new_AGEMA_signal_6211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C ( clk ), .D ( n2336 ), .Q ( new_AGEMA_signal_6213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C ( clk ), .D ( new_AGEMA_signal_1626 ), .Q ( new_AGEMA_signal_6215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C ( clk ), .D ( new_AGEMA_signal_6217 ), .Q ( new_AGEMA_signal_6218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C ( clk ), .D ( new_AGEMA_signal_6220 ), .Q ( new_AGEMA_signal_6221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C ( clk ), .D ( new_AGEMA_signal_6224 ), .Q ( new_AGEMA_signal_6225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C ( clk ), .D ( new_AGEMA_signal_6228 ), .Q ( new_AGEMA_signal_6229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C ( clk ), .D ( new_AGEMA_signal_6233 ), .Q ( new_AGEMA_signal_6234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C ( clk ), .D ( new_AGEMA_signal_6236 ), .Q ( new_AGEMA_signal_6237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C ( clk ), .D ( new_AGEMA_signal_6243 ), .Q ( new_AGEMA_signal_6244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C ( clk ), .D ( new_AGEMA_signal_6246 ), .Q ( new_AGEMA_signal_6247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C ( clk ), .D ( new_AGEMA_signal_6249 ), .Q ( new_AGEMA_signal_6250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C ( clk ), .D ( new_AGEMA_signal_6252 ), .Q ( new_AGEMA_signal_6253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C ( clk ), .D ( new_AGEMA_signal_6256 ), .Q ( new_AGEMA_signal_6257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C ( clk ), .D ( new_AGEMA_signal_6260 ), .Q ( new_AGEMA_signal_6261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C ( clk ), .D ( new_AGEMA_signal_6264 ), .Q ( new_AGEMA_signal_6265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C ( clk ), .D ( new_AGEMA_signal_6268 ), .Q ( new_AGEMA_signal_6269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C ( clk ), .D ( new_AGEMA_signal_6271 ), .Q ( new_AGEMA_signal_6272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C ( clk ), .D ( new_AGEMA_signal_6274 ), .Q ( new_AGEMA_signal_6275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C ( clk ), .D ( new_AGEMA_signal_6277 ), .Q ( new_AGEMA_signal_6278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C ( clk ), .D ( new_AGEMA_signal_6280 ), .Q ( new_AGEMA_signal_6281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C ( clk ), .D ( n2658 ), .Q ( new_AGEMA_signal_6285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C ( clk ), .D ( new_AGEMA_signal_1478 ), .Q ( new_AGEMA_signal_6287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C ( clk ), .D ( n2698 ), .Q ( new_AGEMA_signal_6289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C ( clk ), .D ( new_AGEMA_signal_1573 ), .Q ( new_AGEMA_signal_6291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C ( clk ), .D ( n2800 ), .Q ( new_AGEMA_signal_6293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C ( clk ), .D ( new_AGEMA_signal_1581 ), .Q ( new_AGEMA_signal_6295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C ( clk ), .D ( n1936 ), .Q ( new_AGEMA_signal_6299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C ( clk ), .D ( new_AGEMA_signal_1470 ), .Q ( new_AGEMA_signal_6302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C ( clk ), .D ( new_AGEMA_signal_6311 ), .Q ( new_AGEMA_signal_6312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C ( clk ), .D ( new_AGEMA_signal_6315 ), .Q ( new_AGEMA_signal_6316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C ( clk ), .D ( new_AGEMA_signal_6319 ), .Q ( new_AGEMA_signal_6320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C ( clk ), .D ( new_AGEMA_signal_6323 ), .Q ( new_AGEMA_signal_6324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C ( clk ), .D ( new_AGEMA_signal_6327 ), .Q ( new_AGEMA_signal_6328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C ( clk ), .D ( new_AGEMA_signal_6331 ), .Q ( new_AGEMA_signal_6332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C ( clk ), .D ( new_AGEMA_signal_6335 ), .Q ( new_AGEMA_signal_6336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C ( clk ), .D ( new_AGEMA_signal_6339 ), .Q ( new_AGEMA_signal_6340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C ( clk ), .D ( n2099 ), .Q ( new_AGEMA_signal_6343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C ( clk ), .D ( new_AGEMA_signal_1499 ), .Q ( new_AGEMA_signal_6346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C ( clk ), .D ( new_AGEMA_signal_6350 ), .Q ( new_AGEMA_signal_6351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C ( clk ), .D ( new_AGEMA_signal_6355 ), .Q ( new_AGEMA_signal_6356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C ( clk ), .D ( new_AGEMA_signal_6359 ), .Q ( new_AGEMA_signal_6360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C ( clk ), .D ( new_AGEMA_signal_6363 ), .Q ( new_AGEMA_signal_6364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C ( clk ), .D ( new_AGEMA_signal_6367 ), .Q ( new_AGEMA_signal_6368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C ( clk ), .D ( new_AGEMA_signal_6371 ), .Q ( new_AGEMA_signal_6372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C ( clk ), .D ( new_AGEMA_signal_6375 ), .Q ( new_AGEMA_signal_6376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C ( clk ), .D ( new_AGEMA_signal_6379 ), .Q ( new_AGEMA_signal_6380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C ( clk ), .D ( n2301 ), .Q ( new_AGEMA_signal_6389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C ( clk ), .D ( new_AGEMA_signal_1533 ), .Q ( new_AGEMA_signal_6392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C ( clk ), .D ( new_AGEMA_signal_6400 ), .Q ( new_AGEMA_signal_6401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C ( clk ), .D ( new_AGEMA_signal_6405 ), .Q ( new_AGEMA_signal_6406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C ( clk ), .D ( new_AGEMA_signal_6409 ), .Q ( new_AGEMA_signal_6410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C ( clk ), .D ( new_AGEMA_signal_6413 ), .Q ( new_AGEMA_signal_6414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C ( clk ), .D ( new_AGEMA_signal_6423 ), .Q ( new_AGEMA_signal_6424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C ( clk ), .D ( new_AGEMA_signal_6427 ), .Q ( new_AGEMA_signal_6428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C ( clk ), .D ( new_AGEMA_signal_6431 ), .Q ( new_AGEMA_signal_6432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C ( clk ), .D ( new_AGEMA_signal_6435 ), .Q ( new_AGEMA_signal_6436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C ( clk ), .D ( new_AGEMA_signal_5768 ), .Q ( new_AGEMA_signal_6439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C ( clk ), .D ( new_AGEMA_signal_5770 ), .Q ( new_AGEMA_signal_6442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C ( clk ), .D ( new_AGEMA_signal_6449 ), .Q ( new_AGEMA_signal_6450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C ( clk ), .D ( new_AGEMA_signal_6453 ), .Q ( new_AGEMA_signal_6454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C ( clk ), .D ( new_AGEMA_signal_5880 ), .Q ( new_AGEMA_signal_6481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C ( clk ), .D ( new_AGEMA_signal_5882 ), .Q ( new_AGEMA_signal_6485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C ( clk ), .D ( n2102 ), .Q ( new_AGEMA_signal_6499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C ( clk ), .D ( new_AGEMA_signal_1503 ), .Q ( new_AGEMA_signal_6503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C ( clk ), .D ( new_AGEMA_signal_5727 ), .Q ( new_AGEMA_signal_6507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C ( clk ), .D ( new_AGEMA_signal_5728 ), .Q ( new_AGEMA_signal_6511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C ( clk ), .D ( new_AGEMA_signal_6515 ), .Q ( new_AGEMA_signal_6516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C ( clk ), .D ( new_AGEMA_signal_6520 ), .Q ( new_AGEMA_signal_6521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C ( clk ), .D ( new_AGEMA_signal_5820 ), .Q ( new_AGEMA_signal_6525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C ( clk ), .D ( new_AGEMA_signal_5822 ), .Q ( new_AGEMA_signal_6529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C ( clk ), .D ( n2367 ), .Q ( new_AGEMA_signal_6549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C ( clk ), .D ( new_AGEMA_signal_1400 ), .Q ( new_AGEMA_signal_6553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C ( clk ), .D ( n2591 ), .Q ( new_AGEMA_signal_6565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C ( clk ), .D ( new_AGEMA_signal_1564 ), .Q ( new_AGEMA_signal_6569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C ( clk ), .D ( n2105 ), .Q ( new_AGEMA_signal_6609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C ( clk ), .D ( new_AGEMA_signal_1498 ), .Q ( new_AGEMA_signal_6614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C ( clk ), .D ( n2106 ), .Q ( new_AGEMA_signal_6699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C ( clk ), .D ( new_AGEMA_signal_1357 ), .Q ( new_AGEMA_signal_6705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C ( clk ), .D ( new_AGEMA_signal_6711 ), .Q ( new_AGEMA_signal_6712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C ( clk ), .D ( new_AGEMA_signal_6718 ), .Q ( new_AGEMA_signal_6719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C ( clk ), .D ( new_AGEMA_signal_6733 ), .Q ( new_AGEMA_signal_6734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C ( clk ), .D ( new_AGEMA_signal_6740 ), .Q ( new_AGEMA_signal_6741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C ( clk ), .D ( new_AGEMA_signal_6769 ), .Q ( new_AGEMA_signal_6770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C ( clk ), .D ( new_AGEMA_signal_6777 ), .Q ( new_AGEMA_signal_6778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C ( clk ), .D ( new_AGEMA_signal_6791 ), .Q ( new_AGEMA_signal_6792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C ( clk ), .D ( new_AGEMA_signal_6799 ), .Q ( new_AGEMA_signal_6800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C ( clk ), .D ( n2155 ), .Q ( new_AGEMA_signal_6841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C ( clk ), .D ( new_AGEMA_signal_1359 ), .Q ( new_AGEMA_signal_6849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C ( clk ), .D ( new_AGEMA_signal_6867 ), .Q ( new_AGEMA_signal_6868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C ( clk ), .D ( new_AGEMA_signal_6876 ), .Q ( new_AGEMA_signal_6877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C ( clk ), .D ( new_AGEMA_signal_6917 ), .Q ( new_AGEMA_signal_6918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C ( clk ), .D ( new_AGEMA_signal_6927 ), .Q ( new_AGEMA_signal_6928 ) ) ;

    /* cells in depth 6 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2001 ( .a ({new_AGEMA_signal_1586, n1932}), .b ({new_AGEMA_signal_5894, new_AGEMA_signal_5892}), .clk ( clk ), .r ({Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_1667, n1933}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2051 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5896}), .b ({new_AGEMA_signal_1589, n1955}), .clk ( clk ), .r ({Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644]}), .c ({new_AGEMA_signal_1668, n1958}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2067 ( .a ({new_AGEMA_signal_1479, n1967}), .b ({new_AGEMA_signal_5906, new_AGEMA_signal_5902}), .clk ( clk ), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648]}), .c ({new_AGEMA_signal_1590, n1990}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2104 ( .a ({new_AGEMA_signal_5908, new_AGEMA_signal_5907}), .b ({new_AGEMA_signal_1592, n1977}), .clk ( clk ), .r ({Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_1670, n1982}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2128 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5912}), .b ({new_AGEMA_signal_1594, n1998}), .clk ( clk ), .r ({Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656]}), .c ({new_AGEMA_signal_1671, n1999}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2148 ( .a ({new_AGEMA_signal_1595, n2010}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5919}), .clk ( clk ), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660]}), .c ({new_AGEMA_signal_1672, n2011}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2165 ( .a ({new_AGEMA_signal_1489, n2024}), .b ({new_AGEMA_signal_5926, new_AGEMA_signal_5924}), .clk ( clk ), .r ({Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_1596, n2025}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2179 ( .a ({new_AGEMA_signal_1597, n2035}), .b ({new_AGEMA_signal_5932, new_AGEMA_signal_5929}), .clk ( clk ), .r ({Fresh[2671], Fresh[2670], Fresh[2669], Fresh[2668]}), .c ({new_AGEMA_signal_1674, n2036}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2196 ( .a ({new_AGEMA_signal_1599, n2048}), .b ({new_AGEMA_signal_1600, n2047}), .clk ( clk ), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672]}), .c ({new_AGEMA_signal_1675, n2049}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2207 ( .a ({new_AGEMA_signal_5934, new_AGEMA_signal_5933}), .b ({new_AGEMA_signal_1601, n2059}), .clk ( clk ), .r ({Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_1676, n2072}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2214 ( .a ({new_AGEMA_signal_5940, new_AGEMA_signal_5937}), .b ({new_AGEMA_signal_1602, n2064}), .clk ( clk ), .r ({Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680]}), .c ({new_AGEMA_signal_1677, n2067}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2230 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5943}), .b ({new_AGEMA_signal_1603, n2077}), .clk ( clk ), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684]}), .c ({new_AGEMA_signal_1678, n2078}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2250 ( .a ({new_AGEMA_signal_5948, new_AGEMA_signal_5947}), .b ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .r ({Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_1679, n2097}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2257 ( .a ({new_AGEMA_signal_1605, n2095}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5950}), .clk ( clk ), .r ({Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692]}), .c ({new_AGEMA_signal_1680, n2096}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2275 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5955}), .b ({new_AGEMA_signal_1681, n2117}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696]}), .c ({new_AGEMA_signal_1735, n2128}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2285 ( .a ({new_AGEMA_signal_1607, n2123}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5961}), .clk ( clk ), .r ({Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_1682, n2124}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2301 ( .a ({new_AGEMA_signal_5966, new_AGEMA_signal_5965}), .b ({new_AGEMA_signal_1507, n2135}), .clk ( clk ), .r ({Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704]}), .c ({new_AGEMA_signal_1608, n2148}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2310 ( .a ({new_AGEMA_signal_5972, new_AGEMA_signal_5969}), .b ({new_AGEMA_signal_1609, n2141}), .clk ( clk ), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708]}), .c ({new_AGEMA_signal_1683, n2142}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2325 ( .a ({new_AGEMA_signal_5974, new_AGEMA_signal_5973}), .b ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .r ({Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_1684, n2168}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2332 ( .a ({new_AGEMA_signal_1610, n2166}), .b ({new_AGEMA_signal_1512, n2165}), .clk ( clk ), .r ({Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716]}), .c ({new_AGEMA_signal_1685, n2167}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2347 ( .a ({new_AGEMA_signal_5978, new_AGEMA_signal_5976}), .b ({new_AGEMA_signal_1611, n2180}), .clk ( clk ), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720]}), .c ({new_AGEMA_signal_1686, n2184}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2361 ( .a ({new_AGEMA_signal_5982, new_AGEMA_signal_5980}), .b ({new_AGEMA_signal_1612, n2194}), .clk ( clk ), .r ({Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_1687, n2197}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2373 ( .a ({new_AGEMA_signal_5984, new_AGEMA_signal_5983}), .b ({new_AGEMA_signal_1688, n2204}), .clk ( clk ), .r ({Fresh[2731], Fresh[2730], Fresh[2729], Fresh[2728]}), .c ({new_AGEMA_signal_1741, n2205}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2390 ( .a ({new_AGEMA_signal_5992, new_AGEMA_signal_5988}), .b ({new_AGEMA_signal_1614, n2225}), .clk ( clk ), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732]}), .c ({new_AGEMA_signal_1689, n2232}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2395 ( .a ({new_AGEMA_signal_1519, n2230}), .b ({new_AGEMA_signal_5998, new_AGEMA_signal_5995}), .clk ( clk ), .r ({Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_1615, n2231}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2401 ( .a ({new_AGEMA_signal_6002, new_AGEMA_signal_6000}), .b ({new_AGEMA_signal_1690, n2236}), .clk ( clk ), .r ({Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740]}), .c ({new_AGEMA_signal_1743, n2239}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2413 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6004}), .b ({new_AGEMA_signal_1617, n2247}), .clk ( clk ), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744]}), .c ({new_AGEMA_signal_1691, n2250}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2428 ( .a ({new_AGEMA_signal_5934, new_AGEMA_signal_5933}), .b ({new_AGEMA_signal_1619, n2264}), .clk ( clk ), .r ({Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_1692, n2276}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2439 ( .a ({new_AGEMA_signal_1620, n2271}), .b ({new_AGEMA_signal_6008, new_AGEMA_signal_6007}), .clk ( clk ), .r ({Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752]}), .c ({new_AGEMA_signal_1693, n2272}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2454 ( .a ({new_AGEMA_signal_1527, n2286}), .b ({new_AGEMA_signal_6010, new_AGEMA_signal_6009}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756]}), .c ({new_AGEMA_signal_1621, n2306}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2468 ( .a ({new_AGEMA_signal_1623, n2295}), .b ({new_AGEMA_signal_6014, new_AGEMA_signal_6012}), .clk ( clk ), .r ({Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_1694, n2296}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2489 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6016}), .b ({new_AGEMA_signal_1624, n2322}), .clk ( clk ), .r ({Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764]}), .c ({new_AGEMA_signal_1695, n2324}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2500 ( .a ({new_AGEMA_signal_6020, new_AGEMA_signal_6019}), .b ({new_AGEMA_signal_1625, n2333}), .clk ( clk ), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768]}), .c ({new_AGEMA_signal_1696, n2337}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2511 ( .a ({new_AGEMA_signal_1627, n2345}), .b ({new_AGEMA_signal_6026, new_AGEMA_signal_6023}), .clk ( clk ), .r ({Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_1697, n2350}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2528 ( .a ({new_AGEMA_signal_1628, n2361}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6028}), .clk ( clk ), .r ({Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776]}), .c ({new_AGEMA_signal_1698, n2362}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2550 ( .a ({new_AGEMA_signal_6032, new_AGEMA_signal_6031}), .b ({new_AGEMA_signal_1541, n2388}), .clk ( clk ), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780]}), .c ({new_AGEMA_signal_1629, n2389}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2557 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6034}), .b ({new_AGEMA_signal_1630, n2393}), .clk ( clk ), .r ({Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_1700, n2397}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2568 ( .a ({new_AGEMA_signal_6040, new_AGEMA_signal_6038}), .b ({new_AGEMA_signal_1543, n2405}), .clk ( clk ), .r ({Fresh[2791], Fresh[2790], Fresh[2789], Fresh[2788]}), .c ({new_AGEMA_signal_1631, n2411}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2580 ( .a ({new_AGEMA_signal_6044, new_AGEMA_signal_6042}), .b ({new_AGEMA_signal_1546, n2419}), .clk ( clk ), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792]}), .c ({new_AGEMA_signal_1634, n2420}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2593 ( .a ({new_AGEMA_signal_1635, n2436}), .b ({new_AGEMA_signal_6046, new_AGEMA_signal_6045}), .clk ( clk ), .r ({Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_1703, n2440}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2614 ( .a ({new_AGEMA_signal_6050, new_AGEMA_signal_6048}), .b ({new_AGEMA_signal_1638, n2461}), .clk ( clk ), .r ({Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800]}), .c ({new_AGEMA_signal_1704, n2516}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2621 ( .s ({new_AGEMA_signal_6052, new_AGEMA_signal_6051}), .b ({new_AGEMA_signal_1552, n2469}), .a ({new_AGEMA_signal_6058, new_AGEMA_signal_6055}), .clk ( clk ), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804]}), .c ({new_AGEMA_signal_1639, n2471}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2636 ( .a ({new_AGEMA_signal_6064, new_AGEMA_signal_6061}), .b ({new_AGEMA_signal_1640, n2484}), .clk ( clk ), .r ({Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_1706, n2485}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2644 ( .a ({new_AGEMA_signal_5940, new_AGEMA_signal_5937}), .b ({new_AGEMA_signal_1555, n2491}), .clk ( clk ), .r ({Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812]}), .c ({new_AGEMA_signal_1641, n2502}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2651 ( .a ({new_AGEMA_signal_1642, n2500}), .b ({new_AGEMA_signal_6068, new_AGEMA_signal_6066}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816]}), .c ({new_AGEMA_signal_1707, n2501}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2657 ( .a ({new_AGEMA_signal_6044, new_AGEMA_signal_6042}), .b ({new_AGEMA_signal_1708, n2508}), .clk ( clk ), .r ({Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_1757, n2509}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2671 ( .a ({new_AGEMA_signal_6070, new_AGEMA_signal_6069}), .b ({new_AGEMA_signal_1709, n2526}), .clk ( clk ), .r ({Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824]}), .c ({new_AGEMA_signal_1758, n2527}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2680 ( .a ({new_AGEMA_signal_1645, n2539}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6074}), .clk ( clk ), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828]}), .c ({new_AGEMA_signal_1710, n2550}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2685 ( .a ({new_AGEMA_signal_1646, n2548}), .b ({new_AGEMA_signal_6080, new_AGEMA_signal_6079}), .clk ( clk ), .r ({Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_1711, n2549}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2701 ( .a ({new_AGEMA_signal_1647, n2568}), .b ({new_AGEMA_signal_1648, n2567}), .clk ( clk ), .r ({Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836]}), .c ({new_AGEMA_signal_1712, n2569}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2712 ( .a ({new_AGEMA_signal_1649, n2583}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6082}), .clk ( clk ), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840]}), .c ({new_AGEMA_signal_1713, n2584}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2729 ( .a ({new_AGEMA_signal_6088, new_AGEMA_signal_6086}), .b ({new_AGEMA_signal_1566, n2604}), .clk ( clk ), .r ({Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_1650, n2606}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2740 ( .a ({new_AGEMA_signal_5940, new_AGEMA_signal_5937}), .b ({new_AGEMA_signal_1651, n2621}), .clk ( clk ), .r ({Fresh[2851], Fresh[2850], Fresh[2849], Fresh[2848]}), .c ({new_AGEMA_signal_1715, n2622}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2747 ( .a ({new_AGEMA_signal_1652, n2633}), .b ({new_AGEMA_signal_6092, new_AGEMA_signal_6090}), .clk ( clk ), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852]}), .c ({new_AGEMA_signal_1716, n2634}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2761 ( .a ({new_AGEMA_signal_1654, n2656}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6094}), .clk ( clk ), .r ({Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_1717, n2657}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2783 ( .a ({new_AGEMA_signal_1658, n2696}), .b ({new_AGEMA_signal_6100, new_AGEMA_signal_6098}), .clk ( clk ), .r ({Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860]}), .c ({new_AGEMA_signal_1718, n2697}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2795 ( .a ({new_AGEMA_signal_5934, new_AGEMA_signal_5933}), .b ({new_AGEMA_signal_1659, n2718}), .clk ( clk ), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864]}), .c ({new_AGEMA_signal_1719, n2808}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2802 ( .a ({new_AGEMA_signal_1660, n2730}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6104}), .clk ( clk ), .r ({Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_1720, n2747}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2810 ( .a ({new_AGEMA_signal_1661, n2745}), .b ({new_AGEMA_signal_1662, n2744}), .clk ( clk ), .r ({Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872]}), .c ({new_AGEMA_signal_1721, n2746}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2818 ( .a ({new_AGEMA_signal_1663, n2759}), .b ({new_AGEMA_signal_6110, new_AGEMA_signal_6109}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876]}), .c ({new_AGEMA_signal_1722, n2804}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2824 ( .a ({new_AGEMA_signal_1664, n2771}), .b ({new_AGEMA_signal_6114, new_AGEMA_signal_6112}), .clk ( clk ), .r ({Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_1723, n2802}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2838 ( .a ({new_AGEMA_signal_1582, n2798}), .b ({new_AGEMA_signal_6116, new_AGEMA_signal_6115}), .clk ( clk ), .r ({Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884]}), .c ({new_AGEMA_signal_1665, n2799}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2852 ( .a ({new_AGEMA_signal_1666, n2826}), .b ({new_AGEMA_signal_6122, new_AGEMA_signal_6119}), .clk ( clk ), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888]}), .c ({new_AGEMA_signal_1725, n2827}) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C ( clk ), .D ( n1934 ), .Q ( new_AGEMA_signal_6123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C ( clk ), .D ( new_AGEMA_signal_1585 ), .Q ( new_AGEMA_signal_6124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C ( clk ), .D ( new_AGEMA_signal_6127 ), .Q ( new_AGEMA_signal_6128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C ( clk ), .D ( new_AGEMA_signal_6131 ), .Q ( new_AGEMA_signal_6132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C ( clk ), .D ( n1981 ), .Q ( new_AGEMA_signal_6133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C ( clk ), .D ( new_AGEMA_signal_1593 ), .Q ( new_AGEMA_signal_6134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C ( clk ), .D ( new_AGEMA_signal_6135 ), .Q ( new_AGEMA_signal_6136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C ( clk ), .D ( new_AGEMA_signal_6137 ), .Q ( new_AGEMA_signal_6138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C ( clk ), .D ( new_AGEMA_signal_6141 ), .Q ( new_AGEMA_signal_6142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C ( clk ), .D ( new_AGEMA_signal_6145 ), .Q ( new_AGEMA_signal_6146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C ( clk ), .D ( new_AGEMA_signal_5912 ), .Q ( new_AGEMA_signal_6147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C ( clk ), .D ( new_AGEMA_signal_5916 ), .Q ( new_AGEMA_signal_6148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C ( clk ), .D ( new_AGEMA_signal_6150 ), .Q ( new_AGEMA_signal_6151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C ( clk ), .D ( new_AGEMA_signal_6153 ), .Q ( new_AGEMA_signal_6154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C ( clk ), .D ( new_AGEMA_signal_6155 ), .Q ( new_AGEMA_signal_6156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C ( clk ), .D ( new_AGEMA_signal_6157 ), .Q ( new_AGEMA_signal_6158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C ( clk ), .D ( new_AGEMA_signal_6161 ), .Q ( new_AGEMA_signal_6162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C ( clk ), .D ( new_AGEMA_signal_6165 ), .Q ( new_AGEMA_signal_6166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C ( clk ), .D ( new_AGEMA_signal_6167 ), .Q ( new_AGEMA_signal_6168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C ( clk ), .D ( new_AGEMA_signal_6169 ), .Q ( new_AGEMA_signal_6170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C ( clk ), .D ( new_AGEMA_signal_6172 ), .Q ( new_AGEMA_signal_6173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C ( clk ), .D ( new_AGEMA_signal_6175 ), .Q ( new_AGEMA_signal_6176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C ( clk ), .D ( new_AGEMA_signal_6178 ), .Q ( new_AGEMA_signal_6179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C ( clk ), .D ( new_AGEMA_signal_6181 ), .Q ( new_AGEMA_signal_6182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C ( clk ), .D ( new_AGEMA_signal_6184 ), .Q ( new_AGEMA_signal_6185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C ( clk ), .D ( new_AGEMA_signal_6187 ), .Q ( new_AGEMA_signal_6188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C ( clk ), .D ( new_AGEMA_signal_6190 ), .Q ( new_AGEMA_signal_6191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C ( clk ), .D ( new_AGEMA_signal_6193 ), .Q ( new_AGEMA_signal_6194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C ( clk ), .D ( new_AGEMA_signal_6196 ), .Q ( new_AGEMA_signal_6197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C ( clk ), .D ( new_AGEMA_signal_6199 ), .Q ( new_AGEMA_signal_6200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C ( clk ), .D ( new_AGEMA_signal_6201 ), .Q ( new_AGEMA_signal_6202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C ( clk ), .D ( new_AGEMA_signal_6203 ), .Q ( new_AGEMA_signal_6204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C ( clk ), .D ( new_AGEMA_signal_6207 ), .Q ( new_AGEMA_signal_6208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C ( clk ), .D ( new_AGEMA_signal_6211 ), .Q ( new_AGEMA_signal_6212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C ( clk ), .D ( new_AGEMA_signal_6213 ), .Q ( new_AGEMA_signal_6214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C ( clk ), .D ( new_AGEMA_signal_6215 ), .Q ( new_AGEMA_signal_6216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C ( clk ), .D ( new_AGEMA_signal_6218 ), .Q ( new_AGEMA_signal_6219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C ( clk ), .D ( new_AGEMA_signal_6221 ), .Q ( new_AGEMA_signal_6222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C ( clk ), .D ( new_AGEMA_signal_6225 ), .Q ( new_AGEMA_signal_6226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C ( clk ), .D ( new_AGEMA_signal_6229 ), .Q ( new_AGEMA_signal_6230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C ( clk ), .D ( new_AGEMA_signal_6051 ), .Q ( new_AGEMA_signal_6231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C ( clk ), .D ( new_AGEMA_signal_6052 ), .Q ( new_AGEMA_signal_6232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C ( clk ), .D ( new_AGEMA_signal_6234 ), .Q ( new_AGEMA_signal_6235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C ( clk ), .D ( new_AGEMA_signal_6237 ), .Q ( new_AGEMA_signal_6238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C ( clk ), .D ( n2410 ), .Q ( new_AGEMA_signal_6239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C ( clk ), .D ( new_AGEMA_signal_1632 ), .Q ( new_AGEMA_signal_6240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C ( clk ), .D ( n2421 ), .Q ( new_AGEMA_signal_6241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C ( clk ), .D ( new_AGEMA_signal_1633 ), .Q ( new_AGEMA_signal_6242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C ( clk ), .D ( new_AGEMA_signal_6244 ), .Q ( new_AGEMA_signal_6245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C ( clk ), .D ( new_AGEMA_signal_6247 ), .Q ( new_AGEMA_signal_6248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C ( clk ), .D ( new_AGEMA_signal_6250 ), .Q ( new_AGEMA_signal_6251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C ( clk ), .D ( new_AGEMA_signal_6253 ), .Q ( new_AGEMA_signal_6254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C ( clk ), .D ( new_AGEMA_signal_6257 ), .Q ( new_AGEMA_signal_6258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C ( clk ), .D ( new_AGEMA_signal_6261 ), .Q ( new_AGEMA_signal_6262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C ( clk ), .D ( new_AGEMA_signal_6265 ), .Q ( new_AGEMA_signal_6266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C ( clk ), .D ( new_AGEMA_signal_6269 ), .Q ( new_AGEMA_signal_6270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C ( clk ), .D ( new_AGEMA_signal_6272 ), .Q ( new_AGEMA_signal_6273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C ( clk ), .D ( new_AGEMA_signal_6275 ), .Q ( new_AGEMA_signal_6276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C ( clk ), .D ( new_AGEMA_signal_6278 ), .Q ( new_AGEMA_signal_6279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C ( clk ), .D ( new_AGEMA_signal_6281 ), .Q ( new_AGEMA_signal_6282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C ( clk ), .D ( new_AGEMA_signal_6042 ), .Q ( new_AGEMA_signal_6283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C ( clk ), .D ( new_AGEMA_signal_6044 ), .Q ( new_AGEMA_signal_6284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C ( clk ), .D ( new_AGEMA_signal_6285 ), .Q ( new_AGEMA_signal_6286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C ( clk ), .D ( new_AGEMA_signal_6287 ), .Q ( new_AGEMA_signal_6288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C ( clk ), .D ( new_AGEMA_signal_6289 ), .Q ( new_AGEMA_signal_6290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C ( clk ), .D ( new_AGEMA_signal_6291 ), .Q ( new_AGEMA_signal_6292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C ( clk ), .D ( new_AGEMA_signal_6293 ), .Q ( new_AGEMA_signal_6294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C ( clk ), .D ( new_AGEMA_signal_6295 ), .Q ( new_AGEMA_signal_6296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C ( clk ), .D ( new_AGEMA_signal_5988 ), .Q ( new_AGEMA_signal_6297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C ( clk ), .D ( new_AGEMA_signal_5992 ), .Q ( new_AGEMA_signal_6298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C ( clk ), .D ( new_AGEMA_signal_6299 ), .Q ( new_AGEMA_signal_6300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C ( clk ), .D ( new_AGEMA_signal_6302 ), .Q ( new_AGEMA_signal_6303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C ( clk ), .D ( n1984 ), .Q ( new_AGEMA_signal_6307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C ( clk ), .D ( new_AGEMA_signal_1669 ), .Q ( new_AGEMA_signal_6309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C ( clk ), .D ( new_AGEMA_signal_6312 ), .Q ( new_AGEMA_signal_6313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C ( clk ), .D ( new_AGEMA_signal_6316 ), .Q ( new_AGEMA_signal_6317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C ( clk ), .D ( new_AGEMA_signal_6320 ), .Q ( new_AGEMA_signal_6321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C ( clk ), .D ( new_AGEMA_signal_6324 ), .Q ( new_AGEMA_signal_6325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C ( clk ), .D ( new_AGEMA_signal_6328 ), .Q ( new_AGEMA_signal_6329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C ( clk ), .D ( new_AGEMA_signal_6332 ), .Q ( new_AGEMA_signal_6333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C ( clk ), .D ( new_AGEMA_signal_6336 ), .Q ( new_AGEMA_signal_6337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C ( clk ), .D ( new_AGEMA_signal_6340 ), .Q ( new_AGEMA_signal_6341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C ( clk ), .D ( new_AGEMA_signal_6343 ), .Q ( new_AGEMA_signal_6344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C ( clk ), .D ( new_AGEMA_signal_6346 ), .Q ( new_AGEMA_signal_6347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C ( clk ), .D ( new_AGEMA_signal_6351 ), .Q ( new_AGEMA_signal_6352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C ( clk ), .D ( new_AGEMA_signal_6356 ), .Q ( new_AGEMA_signal_6357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C ( clk ), .D ( new_AGEMA_signal_6360 ), .Q ( new_AGEMA_signal_6361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C ( clk ), .D ( new_AGEMA_signal_6364 ), .Q ( new_AGEMA_signal_6365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C ( clk ), .D ( new_AGEMA_signal_6368 ), .Q ( new_AGEMA_signal_6369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C ( clk ), .D ( new_AGEMA_signal_6372 ), .Q ( new_AGEMA_signal_6373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C ( clk ), .D ( new_AGEMA_signal_6376 ), .Q ( new_AGEMA_signal_6377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C ( clk ), .D ( new_AGEMA_signal_6380 ), .Q ( new_AGEMA_signal_6381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C ( clk ), .D ( new_AGEMA_signal_6048 ), .Q ( new_AGEMA_signal_6385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C ( clk ), .D ( new_AGEMA_signal_6050 ), .Q ( new_AGEMA_signal_6387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C ( clk ), .D ( new_AGEMA_signal_6389 ), .Q ( new_AGEMA_signal_6390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C ( clk ), .D ( new_AGEMA_signal_6392 ), .Q ( new_AGEMA_signal_6393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C ( clk ), .D ( new_AGEMA_signal_5937 ), .Q ( new_AGEMA_signal_6395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C ( clk ), .D ( new_AGEMA_signal_5940 ), .Q ( new_AGEMA_signal_6397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C ( clk ), .D ( new_AGEMA_signal_6401 ), .Q ( new_AGEMA_signal_6402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C ( clk ), .D ( new_AGEMA_signal_6406 ), .Q ( new_AGEMA_signal_6407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C ( clk ), .D ( new_AGEMA_signal_6410 ), .Q ( new_AGEMA_signal_6411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C ( clk ), .D ( new_AGEMA_signal_6414 ), .Q ( new_AGEMA_signal_6415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C ( clk ), .D ( n2478 ), .Q ( new_AGEMA_signal_6417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C ( clk ), .D ( new_AGEMA_signal_1553 ), .Q ( new_AGEMA_signal_6419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C ( clk ), .D ( new_AGEMA_signal_6424 ), .Q ( new_AGEMA_signal_6425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C ( clk ), .D ( new_AGEMA_signal_6428 ), .Q ( new_AGEMA_signal_6429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C ( clk ), .D ( new_AGEMA_signal_6432 ), .Q ( new_AGEMA_signal_6433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C ( clk ), .D ( new_AGEMA_signal_6436 ), .Q ( new_AGEMA_signal_6437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C ( clk ), .D ( new_AGEMA_signal_6439 ), .Q ( new_AGEMA_signal_6440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C ( clk ), .D ( new_AGEMA_signal_6442 ), .Q ( new_AGEMA_signal_6443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C ( clk ), .D ( n2660 ), .Q ( new_AGEMA_signal_6445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_6447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C ( clk ), .D ( new_AGEMA_signal_6450 ), .Q ( new_AGEMA_signal_6451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C ( clk ), .D ( new_AGEMA_signal_6454 ), .Q ( new_AGEMA_signal_6455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C ( clk ), .D ( n1940 ), .Q ( new_AGEMA_signal_6459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C ( clk ), .D ( new_AGEMA_signal_1587 ), .Q ( new_AGEMA_signal_6462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C ( clk ), .D ( n1961 ), .Q ( new_AGEMA_signal_6465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C ( clk ), .D ( new_AGEMA_signal_1588 ), .Q ( new_AGEMA_signal_6468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C ( clk ), .D ( n1987 ), .Q ( new_AGEMA_signal_6471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C ( clk ), .D ( new_AGEMA_signal_1485 ), .Q ( new_AGEMA_signal_6474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C ( clk ), .D ( new_AGEMA_signal_6481 ), .Q ( new_AGEMA_signal_6482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C ( clk ), .D ( new_AGEMA_signal_6485 ), .Q ( new_AGEMA_signal_6486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C ( clk ), .D ( n2054 ), .Q ( new_AGEMA_signal_6489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C ( clk ), .D ( new_AGEMA_signal_1598 ), .Q ( new_AGEMA_signal_6492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C ( clk ), .D ( new_AGEMA_signal_6499 ), .Q ( new_AGEMA_signal_6500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C ( clk ), .D ( new_AGEMA_signal_6503 ), .Q ( new_AGEMA_signal_6504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C ( clk ), .D ( new_AGEMA_signal_6507 ), .Q ( new_AGEMA_signal_6508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C ( clk ), .D ( new_AGEMA_signal_6511 ), .Q ( new_AGEMA_signal_6512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C ( clk ), .D ( new_AGEMA_signal_6516 ), .Q ( new_AGEMA_signal_6517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C ( clk ), .D ( new_AGEMA_signal_6521 ), .Q ( new_AGEMA_signal_6522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C ( clk ), .D ( new_AGEMA_signal_6525 ), .Q ( new_AGEMA_signal_6526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C ( clk ), .D ( new_AGEMA_signal_6529 ), .Q ( new_AGEMA_signal_6530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C ( clk ), .D ( n2255 ), .Q ( new_AGEMA_signal_6533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C ( clk ), .D ( new_AGEMA_signal_1618 ), .Q ( new_AGEMA_signal_6536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C ( clk ), .D ( n2304 ), .Q ( new_AGEMA_signal_6543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C ( clk ), .D ( new_AGEMA_signal_1622 ), .Q ( new_AGEMA_signal_6546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C ( clk ), .D ( new_AGEMA_signal_6549 ), .Q ( new_AGEMA_signal_6550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C ( clk ), .D ( new_AGEMA_signal_6553 ), .Q ( new_AGEMA_signal_6554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C ( clk ), .D ( n2450 ), .Q ( new_AGEMA_signal_6557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C ( clk ), .D ( new_AGEMA_signal_1636 ), .Q ( new_AGEMA_signal_6560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C ( clk ), .D ( new_AGEMA_signal_6565 ), .Q ( new_AGEMA_signal_6566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C ( clk ), .D ( new_AGEMA_signal_6569 ), .Q ( new_AGEMA_signal_6570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C ( clk ), .D ( n2666 ), .Q ( new_AGEMA_signal_6577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C ( clk ), .D ( new_AGEMA_signal_1655 ), .Q ( new_AGEMA_signal_6580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C ( clk ), .D ( n2704 ), .Q ( new_AGEMA_signal_6583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C ( clk ), .D ( new_AGEMA_signal_1657 ), .Q ( new_AGEMA_signal_6586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C ( clk ), .D ( new_AGEMA_signal_6609 ), .Q ( new_AGEMA_signal_6610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C ( clk ), .D ( new_AGEMA_signal_6614 ), .Q ( new_AGEMA_signal_6615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C ( clk ), .D ( n2280 ), .Q ( new_AGEMA_signal_6639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C ( clk ), .D ( new_AGEMA_signal_1526 ), .Q ( new_AGEMA_signal_6643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C ( clk ), .D ( new_AGEMA_signal_5933 ), .Q ( new_AGEMA_signal_6653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C ( clk ), .D ( new_AGEMA_signal_5934 ), .Q ( new_AGEMA_signal_6657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C ( clk ), .D ( n2456 ), .Q ( new_AGEMA_signal_6661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C ( clk ), .D ( new_AGEMA_signal_1637 ), .Q ( new_AGEMA_signal_6665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C ( clk ), .D ( n2706 ), .Q ( new_AGEMA_signal_6679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C ( clk ), .D ( new_AGEMA_signal_1656 ), .Q ( new_AGEMA_signal_6683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C ( clk ), .D ( new_AGEMA_signal_6699 ), .Q ( new_AGEMA_signal_6700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C ( clk ), .D ( new_AGEMA_signal_6705 ), .Q ( new_AGEMA_signal_6706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C ( clk ), .D ( new_AGEMA_signal_6712 ), .Q ( new_AGEMA_signal_6713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C ( clk ), .D ( new_AGEMA_signal_6719 ), .Q ( new_AGEMA_signal_6720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C ( clk ), .D ( new_AGEMA_signal_6734 ), .Q ( new_AGEMA_signal_6735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C ( clk ), .D ( new_AGEMA_signal_6741 ), .Q ( new_AGEMA_signal_6742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C ( clk ), .D ( new_AGEMA_signal_6770 ), .Q ( new_AGEMA_signal_6771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C ( clk ), .D ( new_AGEMA_signal_6778 ), .Q ( new_AGEMA_signal_6779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C ( clk ), .D ( new_AGEMA_signal_6792 ), .Q ( new_AGEMA_signal_6793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C ( clk ), .D ( new_AGEMA_signal_6800 ), .Q ( new_AGEMA_signal_6801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C ( clk ), .D ( new_AGEMA_signal_6841 ), .Q ( new_AGEMA_signal_6842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C ( clk ), .D ( new_AGEMA_signal_6849 ), .Q ( new_AGEMA_signal_6850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C ( clk ), .D ( new_AGEMA_signal_6868 ), .Q ( new_AGEMA_signal_6869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C ( clk ), .D ( new_AGEMA_signal_6877 ), .Q ( new_AGEMA_signal_6878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C ( clk ), .D ( new_AGEMA_signal_6918 ), .Q ( new_AGEMA_signal_6919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C ( clk ), .D ( new_AGEMA_signal_6928 ), .Q ( new_AGEMA_signal_6929 ) ) ;

    /* cells in depth 7 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2002 ( .a ({new_AGEMA_signal_6124, new_AGEMA_signal_6123}), .b ({new_AGEMA_signal_1667, n1933}), .clk ( clk ), .r ({Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_1726, n1935}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2054 ( .a ({new_AGEMA_signal_1668, n1958}), .b ({new_AGEMA_signal_6132, new_AGEMA_signal_6128}), .clk ( clk ), .r ({Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896]}), .c ({new_AGEMA_signal_1727, n1959}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2109 ( .a ({new_AGEMA_signal_1670, n1982}), .b ({new_AGEMA_signal_6134, new_AGEMA_signal_6133}), .clk ( clk ), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900]}), .c ({new_AGEMA_signal_1728, n1983}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2149 ( .a ({new_AGEMA_signal_6138, new_AGEMA_signal_6136}), .b ({new_AGEMA_signal_1672, n2011}), .clk ( clk ), .r ({Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_1729, n2014}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2166 ( .a ({new_AGEMA_signal_6146, new_AGEMA_signal_6142}), .b ({new_AGEMA_signal_1596, n2025}), .clk ( clk ), .r ({Fresh[2911], Fresh[2910], Fresh[2909], Fresh[2908]}), .c ({new_AGEMA_signal_1673, n2029}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2180 ( .a ({new_AGEMA_signal_6148, new_AGEMA_signal_6147}), .b ({new_AGEMA_signal_1674, n2036}), .clk ( clk ), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912]}), .c ({new_AGEMA_signal_1731, n2037}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2197 ( .a ({new_AGEMA_signal_6154, new_AGEMA_signal_6151}), .b ({new_AGEMA_signal_1675, n2049}), .clk ( clk ), .r ({Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_1732, n2052}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2219 ( .a ({new_AGEMA_signal_1677, n2067}), .b ({new_AGEMA_signal_6158, new_AGEMA_signal_6156}), .clk ( clk ), .r ({Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920]}), .c ({new_AGEMA_signal_1733, n2070}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2258 ( .a ({new_AGEMA_signal_1679, n2097}), .b ({new_AGEMA_signal_1680, n2096}), .clk ( clk ), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924]}), .c ({new_AGEMA_signal_1734, n2098}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2287 ( .a ({new_AGEMA_signal_1682, n2124}), .b ({new_AGEMA_signal_6166, new_AGEMA_signal_6162}), .clk ( clk ), .r ({Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_1736, n2125}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2311 ( .a ({new_AGEMA_signal_6170, new_AGEMA_signal_6168}), .b ({new_AGEMA_signal_1683, n2142}), .clk ( clk ), .r ({Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932]}), .c ({new_AGEMA_signal_1737, n2145}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2333 ( .a ({new_AGEMA_signal_1684, n2168}), .b ({new_AGEMA_signal_1685, n2167}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936]}), .c ({new_AGEMA_signal_1738, n2169}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2350 ( .a ({new_AGEMA_signal_1686, n2184}), .b ({new_AGEMA_signal_6176, new_AGEMA_signal_6173}), .clk ( clk ), .r ({Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_1739, n2185}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2365 ( .a ({new_AGEMA_signal_1687, n2197}), .b ({new_AGEMA_signal_6182, new_AGEMA_signal_6179}), .clk ( clk ), .r ({Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944]}), .c ({new_AGEMA_signal_1740, n2198}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2396 ( .a ({new_AGEMA_signal_1689, n2232}), .b ({new_AGEMA_signal_1615, n2231}), .clk ( clk ), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948]}), .c ({new_AGEMA_signal_1742, n2312}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2404 ( .a ({new_AGEMA_signal_1743, n2239}), .b ({new_AGEMA_signal_6188, new_AGEMA_signal_6185}), .clk ( clk ), .r ({Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_1781, n2258}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2415 ( .a ({new_AGEMA_signal_1691, n2250}), .b ({new_AGEMA_signal_6194, new_AGEMA_signal_6191}), .clk ( clk ), .r ({Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956]}), .c ({new_AGEMA_signal_1744, n2251}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2440 ( .a ({new_AGEMA_signal_6200, new_AGEMA_signal_6197}), .b ({new_AGEMA_signal_1693, n2272}), .clk ( clk ), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960]}), .c ({new_AGEMA_signal_1745, n2274}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2469 ( .a ({new_AGEMA_signal_6204, new_AGEMA_signal_6202}), .b ({new_AGEMA_signal_1694, n2296}), .clk ( clk ), .r ({Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_1746, n2302}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2490 ( .a ({new_AGEMA_signal_1695, n2324}), .b ({new_AGEMA_signal_6212, new_AGEMA_signal_6208}), .clk ( clk ), .r ({Fresh[2971], Fresh[2970], Fresh[2969], Fresh[2968]}), .c ({new_AGEMA_signal_1747, n2339}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2503 ( .a ({new_AGEMA_signal_1696, n2337}), .b ({new_AGEMA_signal_6216, new_AGEMA_signal_6214}), .clk ( clk ), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972]}), .c ({new_AGEMA_signal_1748, n2338}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2515 ( .a ({new_AGEMA_signal_1697, n2350}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6219}), .clk ( clk ), .r ({Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_1749, n2351}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2529 ( .a ({new_AGEMA_signal_6230, new_AGEMA_signal_6226}), .b ({new_AGEMA_signal_1698, n2362}), .clk ( clk ), .r ({Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980]}), .c ({new_AGEMA_signal_1750, n2365}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2551 ( .a ({new_AGEMA_signal_1629, n2389}), .b ({new_AGEMA_signal_6232, new_AGEMA_signal_6231}), .clk ( clk ), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984]}), .c ({new_AGEMA_signal_1699, n2399}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2560 ( .a ({new_AGEMA_signal_1700, n2397}), .b ({new_AGEMA_signal_6238, new_AGEMA_signal_6235}), .clk ( clk ), .r ({Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_1751, n2398}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2572 ( .a ({new_AGEMA_signal_1631, n2411}), .b ({new_AGEMA_signal_6240, new_AGEMA_signal_6239}), .clk ( clk ), .r ({Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992]}), .c ({new_AGEMA_signal_1701, n2423}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2581 ( .a ({new_AGEMA_signal_6242, new_AGEMA_signal_6241}), .b ({new_AGEMA_signal_1634, n2420}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996]}), .c ({new_AGEMA_signal_1702, n2422}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2596 ( .a ({new_AGEMA_signal_1703, n2440}), .b ({new_AGEMA_signal_6248, new_AGEMA_signal_6245}), .clk ( clk ), .r ({Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_1753, n2441}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2623 ( .a ({new_AGEMA_signal_1639, n2471}), .b ({new_AGEMA_signal_6254, new_AGEMA_signal_6251}), .clk ( clk ), .r ({Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004]}), .c ({new_AGEMA_signal_1705, n2479}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2637 ( .a ({new_AGEMA_signal_1706, n2485}), .b ({new_AGEMA_signal_6262, new_AGEMA_signal_6258}), .clk ( clk ), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008]}), .c ({new_AGEMA_signal_1755, n2512}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2652 ( .a ({new_AGEMA_signal_1641, n2502}), .b ({new_AGEMA_signal_1707, n2501}), .clk ( clk ), .r ({Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_1756, n2510}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2686 ( .a ({new_AGEMA_signal_1710, n2550}), .b ({new_AGEMA_signal_1711, n2549}), .clk ( clk ), .r ({Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016]}), .c ({new_AGEMA_signal_1759, n2552}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2702 ( .a ({new_AGEMA_signal_6270, new_AGEMA_signal_6266}), .b ({new_AGEMA_signal_1712, n2569}), .clk ( clk ), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020]}), .c ({new_AGEMA_signal_1760, n2593}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2713 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6273}), .b ({new_AGEMA_signal_1713, n2584}), .clk ( clk ), .r ({Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_1761, n2589}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2730 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6279}), .b ({new_AGEMA_signal_1650, n2606}), .clk ( clk ), .r ({Fresh[3031], Fresh[3030], Fresh[3029], Fresh[3028]}), .c ({new_AGEMA_signal_1714, n2608}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2748 ( .a ({new_AGEMA_signal_6284, new_AGEMA_signal_6283}), .b ({new_AGEMA_signal_1716, n2634}), .clk ( clk ), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032]}), .c ({new_AGEMA_signal_1763, n2636}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2762 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6286}), .b ({new_AGEMA_signal_1717, n2657}), .clk ( clk ), .r ({Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_1764, n2659}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2784 ( .a ({new_AGEMA_signal_6292, new_AGEMA_signal_6290}), .b ({new_AGEMA_signal_1718, n2697}), .clk ( clk ), .r ({Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040]}), .c ({new_AGEMA_signal_1765, n2702}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2811 ( .a ({new_AGEMA_signal_1720, n2747}), .b ({new_AGEMA_signal_1721, n2746}), .clk ( clk ), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044]}), .c ({new_AGEMA_signal_1766, n2806}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2839 ( .a ({new_AGEMA_signal_6296, new_AGEMA_signal_6294}), .b ({new_AGEMA_signal_1665, n2799}), .clk ( clk ), .r ({Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_1724, n2801}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2853 ( .a ({new_AGEMA_signal_6298, new_AGEMA_signal_6297}), .b ({new_AGEMA_signal_1725, n2827}), .clk ( clk ), .r ({Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052]}), .c ({new_AGEMA_signal_1768, n2829}) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C ( clk ), .D ( new_AGEMA_signal_6300 ), .Q ( new_AGEMA_signal_6301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C ( clk ), .D ( new_AGEMA_signal_6303 ), .Q ( new_AGEMA_signal_6304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C ( clk ), .D ( new_AGEMA_signal_6286 ), .Q ( new_AGEMA_signal_6305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C ( clk ), .D ( new_AGEMA_signal_6288 ), .Q ( new_AGEMA_signal_6306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C ( clk ), .D ( new_AGEMA_signal_6307 ), .Q ( new_AGEMA_signal_6308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C ( clk ), .D ( new_AGEMA_signal_6309 ), .Q ( new_AGEMA_signal_6310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C ( clk ), .D ( new_AGEMA_signal_6313 ), .Q ( new_AGEMA_signal_6314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C ( clk ), .D ( new_AGEMA_signal_6317 ), .Q ( new_AGEMA_signal_6318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C ( clk ), .D ( new_AGEMA_signal_6321 ), .Q ( new_AGEMA_signal_6322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C ( clk ), .D ( new_AGEMA_signal_6325 ), .Q ( new_AGEMA_signal_6326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C ( clk ), .D ( new_AGEMA_signal_6329 ), .Q ( new_AGEMA_signal_6330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C ( clk ), .D ( new_AGEMA_signal_6333 ), .Q ( new_AGEMA_signal_6334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C ( clk ), .D ( new_AGEMA_signal_6337 ), .Q ( new_AGEMA_signal_6338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C ( clk ), .D ( new_AGEMA_signal_6341 ), .Q ( new_AGEMA_signal_6342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C ( clk ), .D ( new_AGEMA_signal_6344 ), .Q ( new_AGEMA_signal_6345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C ( clk ), .D ( new_AGEMA_signal_6347 ), .Q ( new_AGEMA_signal_6348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C ( clk ), .D ( new_AGEMA_signal_6352 ), .Q ( new_AGEMA_signal_6353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C ( clk ), .D ( new_AGEMA_signal_6357 ), .Q ( new_AGEMA_signal_6358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C ( clk ), .D ( new_AGEMA_signal_6361 ), .Q ( new_AGEMA_signal_6362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C ( clk ), .D ( new_AGEMA_signal_6365 ), .Q ( new_AGEMA_signal_6366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C ( clk ), .D ( new_AGEMA_signal_6369 ), .Q ( new_AGEMA_signal_6370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C ( clk ), .D ( new_AGEMA_signal_6373 ), .Q ( new_AGEMA_signal_6374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C ( clk ), .D ( new_AGEMA_signal_6377 ), .Q ( new_AGEMA_signal_6378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C ( clk ), .D ( new_AGEMA_signal_6381 ), .Q ( new_AGEMA_signal_6382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C ( clk ), .D ( new_AGEMA_signal_6147 ), .Q ( new_AGEMA_signal_6383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C ( clk ), .D ( new_AGEMA_signal_6148 ), .Q ( new_AGEMA_signal_6384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C ( clk ), .D ( new_AGEMA_signal_6385 ), .Q ( new_AGEMA_signal_6386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C ( clk ), .D ( new_AGEMA_signal_6387 ), .Q ( new_AGEMA_signal_6388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C ( clk ), .D ( new_AGEMA_signal_6390 ), .Q ( new_AGEMA_signal_6391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C ( clk ), .D ( new_AGEMA_signal_6393 ), .Q ( new_AGEMA_signal_6394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C ( clk ), .D ( new_AGEMA_signal_6395 ), .Q ( new_AGEMA_signal_6396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C ( clk ), .D ( new_AGEMA_signal_6397 ), .Q ( new_AGEMA_signal_6398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C ( clk ), .D ( new_AGEMA_signal_6402 ), .Q ( new_AGEMA_signal_6403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C ( clk ), .D ( new_AGEMA_signal_6407 ), .Q ( new_AGEMA_signal_6408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C ( clk ), .D ( new_AGEMA_signal_6411 ), .Q ( new_AGEMA_signal_6412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C ( clk ), .D ( new_AGEMA_signal_6415 ), .Q ( new_AGEMA_signal_6416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C ( clk ), .D ( new_AGEMA_signal_6417 ), .Q ( new_AGEMA_signal_6418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C ( clk ), .D ( new_AGEMA_signal_6419 ), .Q ( new_AGEMA_signal_6420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C ( clk ), .D ( n2509 ), .Q ( new_AGEMA_signal_6421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C ( clk ), .D ( new_AGEMA_signal_1757 ), .Q ( new_AGEMA_signal_6422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C ( clk ), .D ( new_AGEMA_signal_6425 ), .Q ( new_AGEMA_signal_6426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C ( clk ), .D ( new_AGEMA_signal_6429 ), .Q ( new_AGEMA_signal_6430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C ( clk ), .D ( new_AGEMA_signal_6433 ), .Q ( new_AGEMA_signal_6434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C ( clk ), .D ( new_AGEMA_signal_6437 ), .Q ( new_AGEMA_signal_6438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C ( clk ), .D ( new_AGEMA_signal_6440 ), .Q ( new_AGEMA_signal_6441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C ( clk ), .D ( new_AGEMA_signal_6443 ), .Q ( new_AGEMA_signal_6444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C ( clk ), .D ( new_AGEMA_signal_6445 ), .Q ( new_AGEMA_signal_6446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C ( clk ), .D ( new_AGEMA_signal_6447 ), .Q ( new_AGEMA_signal_6448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C ( clk ), .D ( new_AGEMA_signal_6451 ), .Q ( new_AGEMA_signal_6452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C ( clk ), .D ( new_AGEMA_signal_6455 ), .Q ( new_AGEMA_signal_6456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C ( clk ), .D ( n2802 ), .Q ( new_AGEMA_signal_6457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C ( clk ), .D ( new_AGEMA_signal_1723 ), .Q ( new_AGEMA_signal_6458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C ( clk ), .D ( new_AGEMA_signal_6459 ), .Q ( new_AGEMA_signal_6460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C ( clk ), .D ( new_AGEMA_signal_6462 ), .Q ( new_AGEMA_signal_6463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C ( clk ), .D ( new_AGEMA_signal_6465 ), .Q ( new_AGEMA_signal_6466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C ( clk ), .D ( new_AGEMA_signal_6468 ), .Q ( new_AGEMA_signal_6469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C ( clk ), .D ( new_AGEMA_signal_6471 ), .Q ( new_AGEMA_signal_6472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C ( clk ), .D ( new_AGEMA_signal_6474 ), .Q ( new_AGEMA_signal_6475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C ( clk ), .D ( new_AGEMA_signal_6297 ), .Q ( new_AGEMA_signal_6477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C ( clk ), .D ( new_AGEMA_signal_6298 ), .Q ( new_AGEMA_signal_6479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C ( clk ), .D ( new_AGEMA_signal_6482 ), .Q ( new_AGEMA_signal_6483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C ( clk ), .D ( new_AGEMA_signal_6486 ), .Q ( new_AGEMA_signal_6487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C ( clk ), .D ( new_AGEMA_signal_6489 ), .Q ( new_AGEMA_signal_6490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C ( clk ), .D ( new_AGEMA_signal_6492 ), .Q ( new_AGEMA_signal_6493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C ( clk ), .D ( n2072 ), .Q ( new_AGEMA_signal_6495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C ( clk ), .D ( new_AGEMA_signal_1676 ), .Q ( new_AGEMA_signal_6497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C ( clk ), .D ( new_AGEMA_signal_6500 ), .Q ( new_AGEMA_signal_6501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C ( clk ), .D ( new_AGEMA_signal_6504 ), .Q ( new_AGEMA_signal_6505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C ( clk ), .D ( new_AGEMA_signal_6508 ), .Q ( new_AGEMA_signal_6509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C ( clk ), .D ( new_AGEMA_signal_6512 ), .Q ( new_AGEMA_signal_6513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C ( clk ), .D ( new_AGEMA_signal_6517 ), .Q ( new_AGEMA_signal_6518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C ( clk ), .D ( new_AGEMA_signal_6522 ), .Q ( new_AGEMA_signal_6523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C ( clk ), .D ( new_AGEMA_signal_6526 ), .Q ( new_AGEMA_signal_6527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C ( clk ), .D ( new_AGEMA_signal_6530 ), .Q ( new_AGEMA_signal_6531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C ( clk ), .D ( new_AGEMA_signal_6533 ), .Q ( new_AGEMA_signal_6534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C ( clk ), .D ( new_AGEMA_signal_6536 ), .Q ( new_AGEMA_signal_6537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C ( clk ), .D ( n2276 ), .Q ( new_AGEMA_signal_6539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C ( clk ), .D ( new_AGEMA_signal_1692 ), .Q ( new_AGEMA_signal_6541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C ( clk ), .D ( new_AGEMA_signal_6543 ), .Q ( new_AGEMA_signal_6544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C ( clk ), .D ( new_AGEMA_signal_6546 ), .Q ( new_AGEMA_signal_6547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C ( clk ), .D ( new_AGEMA_signal_6550 ), .Q ( new_AGEMA_signal_6551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C ( clk ), .D ( new_AGEMA_signal_6554 ), .Q ( new_AGEMA_signal_6555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C ( clk ), .D ( new_AGEMA_signal_6557 ), .Q ( new_AGEMA_signal_6558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C ( clk ), .D ( new_AGEMA_signal_6560 ), .Q ( new_AGEMA_signal_6561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C ( clk ), .D ( new_AGEMA_signal_6566 ), .Q ( new_AGEMA_signal_6567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C ( clk ), .D ( new_AGEMA_signal_6570 ), .Q ( new_AGEMA_signal_6571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C ( clk ), .D ( n2622 ), .Q ( new_AGEMA_signal_6573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C ( clk ), .D ( new_AGEMA_signal_1715 ), .Q ( new_AGEMA_signal_6575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C ( clk ), .D ( new_AGEMA_signal_6577 ), .Q ( new_AGEMA_signal_6578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C ( clk ), .D ( new_AGEMA_signal_6580 ), .Q ( new_AGEMA_signal_6581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C ( clk ), .D ( new_AGEMA_signal_6583 ), .Q ( new_AGEMA_signal_6584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C ( clk ), .D ( new_AGEMA_signal_6586 ), .Q ( new_AGEMA_signal_6587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C ( clk ), .D ( n2804 ), .Q ( new_AGEMA_signal_6589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C ( clk ), .D ( new_AGEMA_signal_1722 ), .Q ( new_AGEMA_signal_6591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C ( clk ), .D ( n1990 ), .Q ( new_AGEMA_signal_6593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C ( clk ), .D ( new_AGEMA_signal_1590 ), .Q ( new_AGEMA_signal_6596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C ( clk ), .D ( n2078 ), .Q ( new_AGEMA_signal_6603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C ( clk ), .D ( new_AGEMA_signal_1678 ), .Q ( new_AGEMA_signal_6606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C ( clk ), .D ( new_AGEMA_signal_6610 ), .Q ( new_AGEMA_signal_6611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C ( clk ), .D ( new_AGEMA_signal_6615 ), .Q ( new_AGEMA_signal_6616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C ( clk ), .D ( n2128 ), .Q ( new_AGEMA_signal_6619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C ( clk ), .D ( new_AGEMA_signal_1735 ), .Q ( new_AGEMA_signal_6622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C ( clk ), .D ( n2148 ), .Q ( new_AGEMA_signal_6625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_6628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C ( clk ), .D ( new_AGEMA_signal_6639 ), .Q ( new_AGEMA_signal_6640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C ( clk ), .D ( new_AGEMA_signal_6643 ), .Q ( new_AGEMA_signal_6644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C ( clk ), .D ( n2306 ), .Q ( new_AGEMA_signal_6647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C ( clk ), .D ( new_AGEMA_signal_1621 ), .Q ( new_AGEMA_signal_6650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C ( clk ), .D ( new_AGEMA_signal_6653 ), .Q ( new_AGEMA_signal_6654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C ( clk ), .D ( new_AGEMA_signal_6657 ), .Q ( new_AGEMA_signal_6658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C ( clk ), .D ( new_AGEMA_signal_6661 ), .Q ( new_AGEMA_signal_6662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C ( clk ), .D ( new_AGEMA_signal_6665 ), .Q ( new_AGEMA_signal_6666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C ( clk ), .D ( new_AGEMA_signal_6679 ), .Q ( new_AGEMA_signal_6680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C ( clk ), .D ( new_AGEMA_signal_6683 ), .Q ( new_AGEMA_signal_6684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C ( clk ), .D ( n1999 ), .Q ( new_AGEMA_signal_6691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C ( clk ), .D ( new_AGEMA_signal_1671 ), .Q ( new_AGEMA_signal_6695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C ( clk ), .D ( new_AGEMA_signal_6700 ), .Q ( new_AGEMA_signal_6701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C ( clk ), .D ( new_AGEMA_signal_6706 ), .Q ( new_AGEMA_signal_6707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C ( clk ), .D ( new_AGEMA_signal_6713 ), .Q ( new_AGEMA_signal_6714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C ( clk ), .D ( new_AGEMA_signal_6720 ), .Q ( new_AGEMA_signal_6721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C ( clk ), .D ( n2205 ), .Q ( new_AGEMA_signal_6725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C ( clk ), .D ( new_AGEMA_signal_1741 ), .Q ( new_AGEMA_signal_6729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C ( clk ), .D ( new_AGEMA_signal_6735 ), .Q ( new_AGEMA_signal_6736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C ( clk ), .D ( new_AGEMA_signal_6742 ), .Q ( new_AGEMA_signal_6743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C ( clk ), .D ( n2516 ), .Q ( new_AGEMA_signal_6747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C ( clk ), .D ( new_AGEMA_signal_1704 ), .Q ( new_AGEMA_signal_6751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C ( clk ), .D ( n2808 ), .Q ( new_AGEMA_signal_6755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C ( clk ), .D ( new_AGEMA_signal_1719 ), .Q ( new_AGEMA_signal_6759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C ( clk ), .D ( new_AGEMA_signal_6771 ), .Q ( new_AGEMA_signal_6772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C ( clk ), .D ( new_AGEMA_signal_6779 ), .Q ( new_AGEMA_signal_6780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C ( clk ), .D ( new_AGEMA_signal_6793 ), .Q ( new_AGEMA_signal_6794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C ( clk ), .D ( new_AGEMA_signal_6801 ), .Q ( new_AGEMA_signal_6802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C ( clk ), .D ( n2527 ), .Q ( new_AGEMA_signal_6807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C ( clk ), .D ( new_AGEMA_signal_1758 ), .Q ( new_AGEMA_signal_6812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C ( clk ), .D ( new_AGEMA_signal_6842 ), .Q ( new_AGEMA_signal_6843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C ( clk ), .D ( new_AGEMA_signal_6850 ), .Q ( new_AGEMA_signal_6851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C ( clk ), .D ( new_AGEMA_signal_6869 ), .Q ( new_AGEMA_signal_6870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C ( clk ), .D ( new_AGEMA_signal_6878 ), .Q ( new_AGEMA_signal_6879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C ( clk ), .D ( new_AGEMA_signal_6919 ), .Q ( new_AGEMA_signal_6920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C ( clk ), .D ( new_AGEMA_signal_6929 ), .Q ( new_AGEMA_signal_6930 ) ) ;

    /* cells in depth 8 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2003 ( .a ({new_AGEMA_signal_6304, new_AGEMA_signal_6301}), .b ({new_AGEMA_signal_1726, n1935}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056]}), .c ({new_AGEMA_signal_1769, n1941}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2059 ( .a ({new_AGEMA_signal_1727, n1959}), .b ({new_AGEMA_signal_6306, new_AGEMA_signal_6305}), .clk ( clk ), .r ({Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_1770, n1960}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2110 ( .a ({new_AGEMA_signal_6310, new_AGEMA_signal_6308}), .b ({new_AGEMA_signal_1728, n1983}), .clk ( clk ), .r ({Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064]}), .c ({new_AGEMA_signal_1771, n1988}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2153 ( .a ({new_AGEMA_signal_1729, n2014}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6314}), .clk ( clk ), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068]}), .c ({new_AGEMA_signal_1772, n2015}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2169 ( .a ({new_AGEMA_signal_1673, n2029}), .b ({new_AGEMA_signal_6326, new_AGEMA_signal_6322}), .clk ( clk ), .r ({Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_1730, n2030}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2200 ( .a ({new_AGEMA_signal_1732, n2052}), .b ({new_AGEMA_signal_6334, new_AGEMA_signal_6330}), .clk ( clk ), .r ({Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076]}), .c ({new_AGEMA_signal_1774, n2053}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2222 ( .a ({new_AGEMA_signal_1733, n2070}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6338}), .clk ( clk ), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080]}), .c ({new_AGEMA_signal_1775, n2071}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2259 ( .a ({new_AGEMA_signal_6348, new_AGEMA_signal_6345}), .b ({new_AGEMA_signal_1734, n2098}), .clk ( clk ), .r ({Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_1776, n2103}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2288 ( .a ({new_AGEMA_signal_6358, new_AGEMA_signal_6353}), .b ({new_AGEMA_signal_1736, n2125}), .clk ( clk ), .r ({Fresh[3091], Fresh[3090], Fresh[3089], Fresh[3088]}), .c ({new_AGEMA_signal_1777, n2126}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2314 ( .a ({new_AGEMA_signal_1737, n2145}), .b ({new_AGEMA_signal_6366, new_AGEMA_signal_6362}), .clk ( clk ), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092]}), .c ({new_AGEMA_signal_1778, n2146}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2334 ( .a ({new_AGEMA_signal_6374, new_AGEMA_signal_6370}), .b ({new_AGEMA_signal_1738, n2169}), .clk ( clk ), .r ({Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_1779, n2173}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2351 ( .a ({new_AGEMA_signal_6382, new_AGEMA_signal_6378}), .b ({new_AGEMA_signal_1739, n2185}), .clk ( clk ), .r ({Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100]}), .c ({new_AGEMA_signal_1780, n2187}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2416 ( .a ({new_AGEMA_signal_6384, new_AGEMA_signal_6383}), .b ({new_AGEMA_signal_1744, n2251}), .clk ( clk ), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104]}), .c ({new_AGEMA_signal_1782, n2256}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2441 ( .a ({new_AGEMA_signal_1745, n2274}), .b ({new_AGEMA_signal_6388, new_AGEMA_signal_6386}), .clk ( clk ), .r ({Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_1783, n2275}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2474 ( .a ({new_AGEMA_signal_1746, n2302}), .b ({new_AGEMA_signal_6394, new_AGEMA_signal_6391}), .clk ( clk ), .r ({Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112]}), .c ({new_AGEMA_signal_1784, n2303}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2504 ( .a ({new_AGEMA_signal_1747, n2339}), .b ({new_AGEMA_signal_1748, n2338}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116]}), .c ({new_AGEMA_signal_1785, n2382}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2516 ( .a ({new_AGEMA_signal_1749, n2351}), .b ({new_AGEMA_signal_6398, new_AGEMA_signal_6396}), .clk ( clk ), .r ({Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_1786, n2380}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2531 ( .a ({new_AGEMA_signal_1750, n2365}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6403}), .clk ( clk ), .r ({Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124]}), .c ({new_AGEMA_signal_1787, n2366}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2561 ( .a ({new_AGEMA_signal_1699, n2399}), .b ({new_AGEMA_signal_1751, n2398}), .clk ( clk ), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128]}), .c ({new_AGEMA_signal_1788, n2425}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2582 ( .a ({new_AGEMA_signal_1701, n2423}), .b ({new_AGEMA_signal_1702, n2422}), .clk ( clk ), .r ({Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_1752, n2424}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2597 ( .a ({new_AGEMA_signal_6416, new_AGEMA_signal_6412}), .b ({new_AGEMA_signal_1753, n2441}), .clk ( clk ), .r ({Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136]}), .c ({new_AGEMA_signal_1789, n2451}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2631 ( .a ({new_AGEMA_signal_1705, n2479}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6418}), .clk ( clk ), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140]}), .c ({new_AGEMA_signal_1754, n2514}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2658 ( .a ({new_AGEMA_signal_1756, n2510}), .b ({new_AGEMA_signal_6422, new_AGEMA_signal_6421}), .clk ( clk ), .r ({Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_1790, n2511}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2688 ( .a ({new_AGEMA_signal_1759, n2552}), .b ({new_AGEMA_signal_6430, new_AGEMA_signal_6426}), .clk ( clk ), .r ({Fresh[3151], Fresh[3150], Fresh[3149], Fresh[3148]}), .c ({new_AGEMA_signal_1791, n2671}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2716 ( .a ({new_AGEMA_signal_1761, n2589}), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6434}), .clk ( clk ), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152]}), .c ({new_AGEMA_signal_1792, n2590}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2731 ( .a ({new_AGEMA_signal_1714, n2608}), .b ({new_AGEMA_signal_6444, new_AGEMA_signal_6441}), .clk ( clk ), .r ({Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_1762, n2623}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2763 ( .a ({new_AGEMA_signal_6448, new_AGEMA_signal_6446}), .b ({new_AGEMA_signal_1764, n2659}), .clk ( clk ), .r ({Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160]}), .c ({new_AGEMA_signal_1794, n2667}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2786 ( .a ({new_AGEMA_signal_1765, n2702}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6452}), .clk ( clk ), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164]}), .c ({new_AGEMA_signal_1795, n2703}) ) ;
    mux2_GHPC #(.low_latency(1), .pipeline(1)) U2840 ( .s ({new_AGEMA_signal_6388, new_AGEMA_signal_6386}), .b ({new_AGEMA_signal_6458, new_AGEMA_signal_6457}), .a ({new_AGEMA_signal_1724, n2801}), .clk ( clk ), .r ({Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_1767, n2803}) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C ( clk ), .D ( new_AGEMA_signal_6460 ), .Q ( new_AGEMA_signal_6461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C ( clk ), .D ( new_AGEMA_signal_6463 ), .Q ( new_AGEMA_signal_6464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C ( clk ), .D ( new_AGEMA_signal_6466 ), .Q ( new_AGEMA_signal_6467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C ( clk ), .D ( new_AGEMA_signal_6469 ), .Q ( new_AGEMA_signal_6470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C ( clk ), .D ( new_AGEMA_signal_6472 ), .Q ( new_AGEMA_signal_6473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C ( clk ), .D ( new_AGEMA_signal_6475 ), .Q ( new_AGEMA_signal_6476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C ( clk ), .D ( new_AGEMA_signal_6477 ), .Q ( new_AGEMA_signal_6478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C ( clk ), .D ( new_AGEMA_signal_6479 ), .Q ( new_AGEMA_signal_6480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C ( clk ), .D ( new_AGEMA_signal_6483 ), .Q ( new_AGEMA_signal_6484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C ( clk ), .D ( new_AGEMA_signal_6487 ), .Q ( new_AGEMA_signal_6488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C ( clk ), .D ( new_AGEMA_signal_6490 ), .Q ( new_AGEMA_signal_6491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C ( clk ), .D ( new_AGEMA_signal_6493 ), .Q ( new_AGEMA_signal_6494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C ( clk ), .D ( new_AGEMA_signal_6495 ), .Q ( new_AGEMA_signal_6496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C ( clk ), .D ( new_AGEMA_signal_6497 ), .Q ( new_AGEMA_signal_6498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C ( clk ), .D ( new_AGEMA_signal_6501 ), .Q ( new_AGEMA_signal_6502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C ( clk ), .D ( new_AGEMA_signal_6505 ), .Q ( new_AGEMA_signal_6506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C ( clk ), .D ( new_AGEMA_signal_6509 ), .Q ( new_AGEMA_signal_6510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C ( clk ), .D ( new_AGEMA_signal_6513 ), .Q ( new_AGEMA_signal_6514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C ( clk ), .D ( new_AGEMA_signal_6518 ), .Q ( new_AGEMA_signal_6519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C ( clk ), .D ( new_AGEMA_signal_6523 ), .Q ( new_AGEMA_signal_6524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C ( clk ), .D ( new_AGEMA_signal_6527 ), .Q ( new_AGEMA_signal_6528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C ( clk ), .D ( new_AGEMA_signal_6531 ), .Q ( new_AGEMA_signal_6532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C ( clk ), .D ( new_AGEMA_signal_6534 ), .Q ( new_AGEMA_signal_6535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C ( clk ), .D ( new_AGEMA_signal_6537 ), .Q ( new_AGEMA_signal_6538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C ( clk ), .D ( new_AGEMA_signal_6539 ), .Q ( new_AGEMA_signal_6540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C ( clk ), .D ( new_AGEMA_signal_6541 ), .Q ( new_AGEMA_signal_6542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C ( clk ), .D ( new_AGEMA_signal_6544 ), .Q ( new_AGEMA_signal_6545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C ( clk ), .D ( new_AGEMA_signal_6547 ), .Q ( new_AGEMA_signal_6548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C ( clk ), .D ( new_AGEMA_signal_6551 ), .Q ( new_AGEMA_signal_6552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C ( clk ), .D ( new_AGEMA_signal_6555 ), .Q ( new_AGEMA_signal_6556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C ( clk ), .D ( new_AGEMA_signal_6558 ), .Q ( new_AGEMA_signal_6559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C ( clk ), .D ( new_AGEMA_signal_6561 ), .Q ( new_AGEMA_signal_6562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C ( clk ), .D ( n2512 ), .Q ( new_AGEMA_signal_6563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C ( clk ), .D ( new_AGEMA_signal_1755 ), .Q ( new_AGEMA_signal_6564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C ( clk ), .D ( new_AGEMA_signal_6567 ), .Q ( new_AGEMA_signal_6568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C ( clk ), .D ( new_AGEMA_signal_6571 ), .Q ( new_AGEMA_signal_6572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C ( clk ), .D ( new_AGEMA_signal_6573 ), .Q ( new_AGEMA_signal_6574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C ( clk ), .D ( new_AGEMA_signal_6575 ), .Q ( new_AGEMA_signal_6576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C ( clk ), .D ( new_AGEMA_signal_6578 ), .Q ( new_AGEMA_signal_6579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C ( clk ), .D ( new_AGEMA_signal_6581 ), .Q ( new_AGEMA_signal_6582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C ( clk ), .D ( new_AGEMA_signal_6584 ), .Q ( new_AGEMA_signal_6585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C ( clk ), .D ( new_AGEMA_signal_6587 ), .Q ( new_AGEMA_signal_6588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C ( clk ), .D ( new_AGEMA_signal_6589 ), .Q ( new_AGEMA_signal_6590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C ( clk ), .D ( new_AGEMA_signal_6591 ), .Q ( new_AGEMA_signal_6592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C ( clk ), .D ( new_AGEMA_signal_6593 ), .Q ( new_AGEMA_signal_6594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C ( clk ), .D ( new_AGEMA_signal_6596 ), .Q ( new_AGEMA_signal_6597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C ( clk ), .D ( n2037 ), .Q ( new_AGEMA_signal_6599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C ( clk ), .D ( new_AGEMA_signal_1731 ), .Q ( new_AGEMA_signal_6601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C ( clk ), .D ( new_AGEMA_signal_6603 ), .Q ( new_AGEMA_signal_6604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C ( clk ), .D ( new_AGEMA_signal_6606 ), .Q ( new_AGEMA_signal_6607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C ( clk ), .D ( new_AGEMA_signal_6611 ), .Q ( new_AGEMA_signal_6612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C ( clk ), .D ( new_AGEMA_signal_6616 ), .Q ( new_AGEMA_signal_6617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C ( clk ), .D ( new_AGEMA_signal_6619 ), .Q ( new_AGEMA_signal_6620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C ( clk ), .D ( new_AGEMA_signal_6622 ), .Q ( new_AGEMA_signal_6623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C ( clk ), .D ( new_AGEMA_signal_6625 ), .Q ( new_AGEMA_signal_6626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C ( clk ), .D ( new_AGEMA_signal_6628 ), .Q ( new_AGEMA_signal_6629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C ( clk ), .D ( n2198 ), .Q ( new_AGEMA_signal_6631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C ( clk ), .D ( new_AGEMA_signal_1740 ), .Q ( new_AGEMA_signal_6633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C ( clk ), .D ( n2258 ), .Q ( new_AGEMA_signal_6635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C ( clk ), .D ( new_AGEMA_signal_1781 ), .Q ( new_AGEMA_signal_6637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C ( clk ), .D ( new_AGEMA_signal_6640 ), .Q ( new_AGEMA_signal_6641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C ( clk ), .D ( new_AGEMA_signal_6644 ), .Q ( new_AGEMA_signal_6645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C ( clk ), .D ( new_AGEMA_signal_6647 ), .Q ( new_AGEMA_signal_6648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C ( clk ), .D ( new_AGEMA_signal_6650 ), .Q ( new_AGEMA_signal_6651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C ( clk ), .D ( new_AGEMA_signal_6654 ), .Q ( new_AGEMA_signal_6655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C ( clk ), .D ( new_AGEMA_signal_6658 ), .Q ( new_AGEMA_signal_6659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C ( clk ), .D ( new_AGEMA_signal_6662 ), .Q ( new_AGEMA_signal_6663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C ( clk ), .D ( new_AGEMA_signal_6666 ), .Q ( new_AGEMA_signal_6667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C ( clk ), .D ( n2593 ), .Q ( new_AGEMA_signal_6671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C ( clk ), .D ( new_AGEMA_signal_1760 ), .Q ( new_AGEMA_signal_6673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C ( clk ), .D ( n2636 ), .Q ( new_AGEMA_signal_6675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_6677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C ( clk ), .D ( new_AGEMA_signal_6680 ), .Q ( new_AGEMA_signal_6681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C ( clk ), .D ( new_AGEMA_signal_6684 ), .Q ( new_AGEMA_signal_6685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C ( clk ), .D ( n2806 ), .Q ( new_AGEMA_signal_6687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_6689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C ( clk ), .D ( new_AGEMA_signal_6691 ), .Q ( new_AGEMA_signal_6692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C ( clk ), .D ( new_AGEMA_signal_6695 ), .Q ( new_AGEMA_signal_6696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C ( clk ), .D ( new_AGEMA_signal_6701 ), .Q ( new_AGEMA_signal_6702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C ( clk ), .D ( new_AGEMA_signal_6707 ), .Q ( new_AGEMA_signal_6708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C ( clk ), .D ( new_AGEMA_signal_6714 ), .Q ( new_AGEMA_signal_6715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C ( clk ), .D ( new_AGEMA_signal_6721 ), .Q ( new_AGEMA_signal_6722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C ( clk ), .D ( new_AGEMA_signal_6725 ), .Q ( new_AGEMA_signal_6726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C ( clk ), .D ( new_AGEMA_signal_6729 ), .Q ( new_AGEMA_signal_6730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C ( clk ), .D ( new_AGEMA_signal_6736 ), .Q ( new_AGEMA_signal_6737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C ( clk ), .D ( new_AGEMA_signal_6743 ), .Q ( new_AGEMA_signal_6744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C ( clk ), .D ( new_AGEMA_signal_6747 ), .Q ( new_AGEMA_signal_6748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C ( clk ), .D ( new_AGEMA_signal_6751 ), .Q ( new_AGEMA_signal_6752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C ( clk ), .D ( new_AGEMA_signal_6755 ), .Q ( new_AGEMA_signal_6756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C ( clk ), .D ( new_AGEMA_signal_6759 ), .Q ( new_AGEMA_signal_6760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C ( clk ), .D ( new_AGEMA_signal_6772 ), .Q ( new_AGEMA_signal_6773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C ( clk ), .D ( new_AGEMA_signal_6780 ), .Q ( new_AGEMA_signal_6781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C ( clk ), .D ( new_AGEMA_signal_6794 ), .Q ( new_AGEMA_signal_6795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C ( clk ), .D ( new_AGEMA_signal_6802 ), .Q ( new_AGEMA_signal_6803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C ( clk ), .D ( new_AGEMA_signal_6807 ), .Q ( new_AGEMA_signal_6808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C ( clk ), .D ( new_AGEMA_signal_6812 ), .Q ( new_AGEMA_signal_6813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C ( clk ), .D ( n2829 ), .Q ( new_AGEMA_signal_6821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C ( clk ), .D ( new_AGEMA_signal_1768 ), .Q ( new_AGEMA_signal_6825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C ( clk ), .D ( new_AGEMA_signal_6843 ), .Q ( new_AGEMA_signal_6844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C ( clk ), .D ( new_AGEMA_signal_6851 ), .Q ( new_AGEMA_signal_6852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C ( clk ), .D ( n2312 ), .Q ( new_AGEMA_signal_6857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C ( clk ), .D ( new_AGEMA_signal_1742 ), .Q ( new_AGEMA_signal_6862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C ( clk ), .D ( new_AGEMA_signal_6870 ), .Q ( new_AGEMA_signal_6871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C ( clk ), .D ( new_AGEMA_signal_6879 ), .Q ( new_AGEMA_signal_6880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C ( clk ), .D ( new_AGEMA_signal_6920 ), .Q ( new_AGEMA_signal_6921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C ( clk ), .D ( new_AGEMA_signal_6930 ), .Q ( new_AGEMA_signal_6931 ) ) ;

    /* cells in depth 9 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2016 ( .a ({new_AGEMA_signal_1769, n1941}), .b ({new_AGEMA_signal_6464, new_AGEMA_signal_6461}), .clk ( clk ), .r ({Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172]}), .c ({new_AGEMA_signal_1797, n2019}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2060 ( .a ({new_AGEMA_signal_6470, new_AGEMA_signal_6467}), .b ({new_AGEMA_signal_1770, n1960}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176]}), .c ({new_AGEMA_signal_1798, n2002}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2116 ( .a ({new_AGEMA_signal_1771, n1988}), .b ({new_AGEMA_signal_6476, new_AGEMA_signal_6473}), .clk ( clk ), .r ({Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_1799, n1989}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2154 ( .a ({new_AGEMA_signal_6480, new_AGEMA_signal_6478}), .b ({new_AGEMA_signal_1772, n2015}), .clk ( clk ), .r ({Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184]}), .c ({new_AGEMA_signal_1800, n2016}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2170 ( .a ({new_AGEMA_signal_6488, new_AGEMA_signal_6484}), .b ({new_AGEMA_signal_1730, n2030}), .clk ( clk ), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188]}), .c ({new_AGEMA_signal_1773, n2038}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2201 ( .a ({new_AGEMA_signal_6494, new_AGEMA_signal_6491}), .b ({new_AGEMA_signal_1774, n2053}), .clk ( clk ), .r ({Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_1802, n2111}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2223 ( .a ({new_AGEMA_signal_6498, new_AGEMA_signal_6496}), .b ({new_AGEMA_signal_1775, n2071}), .clk ( clk ), .r ({Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196]}), .c ({new_AGEMA_signal_1803, n2079}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2263 ( .a ({new_AGEMA_signal_1776, n2103}), .b ({new_AGEMA_signal_6506, new_AGEMA_signal_6502}), .clk ( clk ), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200]}), .c ({new_AGEMA_signal_1804, n2104}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2289 ( .a ({new_AGEMA_signal_6514, new_AGEMA_signal_6510}), .b ({new_AGEMA_signal_1777, n2126}), .clk ( clk ), .r ({Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_1805, n2127}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2315 ( .a ({new_AGEMA_signal_6480, new_AGEMA_signal_6478}), .b ({new_AGEMA_signal_1778, n2146}), .clk ( clk ), .r ({Fresh[3211], Fresh[3210], Fresh[3209], Fresh[3208]}), .c ({new_AGEMA_signal_1806, n2147}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2336 ( .a ({new_AGEMA_signal_1779, n2173}), .b ({new_AGEMA_signal_6524, new_AGEMA_signal_6519}), .clk ( clk ), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212]}), .c ({new_AGEMA_signal_1807, n2208}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2352 ( .a ({new_AGEMA_signal_1780, n2187}), .b ({new_AGEMA_signal_6532, new_AGEMA_signal_6528}), .clk ( clk ), .r ({Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_1808, n2199}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2420 ( .a ({new_AGEMA_signal_1782, n2256}), .b ({new_AGEMA_signal_6538, new_AGEMA_signal_6535}), .clk ( clk ), .r ({Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220]}), .c ({new_AGEMA_signal_1809, n2257}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2442 ( .a ({new_AGEMA_signal_6542, new_AGEMA_signal_6540}), .b ({new_AGEMA_signal_1783, n2275}), .clk ( clk ), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224]}), .c ({new_AGEMA_signal_1810, n2281}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2475 ( .a ({new_AGEMA_signal_6548, new_AGEMA_signal_6545}), .b ({new_AGEMA_signal_1784, n2303}), .clk ( clk ), .r ({Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_1811, n2305}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2532 ( .a ({new_AGEMA_signal_6556, new_AGEMA_signal_6552}), .b ({new_AGEMA_signal_1787, n2366}), .clk ( clk ), .r ({Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232]}), .c ({new_AGEMA_signal_1812, n2368}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2583 ( .a ({new_AGEMA_signal_1788, n2425}), .b ({new_AGEMA_signal_1752, n2424}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236]}), .c ({new_AGEMA_signal_1813, n2426}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2605 ( .a ({new_AGEMA_signal_1789, n2451}), .b ({new_AGEMA_signal_6562, new_AGEMA_signal_6559}), .clk ( clk ), .r ({Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_1814, n2457}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2659 ( .a ({new_AGEMA_signal_6564, new_AGEMA_signal_6563}), .b ({new_AGEMA_signal_1790, n2511}), .clk ( clk ), .r ({Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244]}), .c ({new_AGEMA_signal_1815, n2513}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2717 ( .a ({new_AGEMA_signal_6572, new_AGEMA_signal_6568}), .b ({new_AGEMA_signal_1792, n2590}), .clk ( clk ), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248]}), .c ({new_AGEMA_signal_1816, n2592}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2741 ( .a ({new_AGEMA_signal_1762, n2623}), .b ({new_AGEMA_signal_6576, new_AGEMA_signal_6574}), .clk ( clk ), .r ({Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_1793, n2637}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2767 ( .a ({new_AGEMA_signal_1794, n2667}), .b ({new_AGEMA_signal_6582, new_AGEMA_signal_6579}), .clk ( clk ), .r ({Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256]}), .c ({new_AGEMA_signal_1818, n2668}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2787 ( .a ({new_AGEMA_signal_6588, new_AGEMA_signal_6585}), .b ({new_AGEMA_signal_1795, n2703}), .clk ( clk ), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260]}), .c ({new_AGEMA_signal_1819, n2705}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2841 ( .a ({new_AGEMA_signal_6592, new_AGEMA_signal_6590}), .b ({new_AGEMA_signal_1767, n2803}), .clk ( clk ), .r ({Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_1796, n2805}) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C ( clk ), .D ( new_AGEMA_signal_6594 ), .Q ( new_AGEMA_signal_6595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C ( clk ), .D ( new_AGEMA_signal_6597 ), .Q ( new_AGEMA_signal_6598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C ( clk ), .D ( new_AGEMA_signal_6599 ), .Q ( new_AGEMA_signal_6600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C ( clk ), .D ( new_AGEMA_signal_6601 ), .Q ( new_AGEMA_signal_6602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C ( clk ), .D ( new_AGEMA_signal_6604 ), .Q ( new_AGEMA_signal_6605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C ( clk ), .D ( new_AGEMA_signal_6607 ), .Q ( new_AGEMA_signal_6608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C ( clk ), .D ( new_AGEMA_signal_6612 ), .Q ( new_AGEMA_signal_6613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C ( clk ), .D ( new_AGEMA_signal_6617 ), .Q ( new_AGEMA_signal_6618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C ( clk ), .D ( new_AGEMA_signal_6620 ), .Q ( new_AGEMA_signal_6621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C ( clk ), .D ( new_AGEMA_signal_6623 ), .Q ( new_AGEMA_signal_6624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C ( clk ), .D ( new_AGEMA_signal_6626 ), .Q ( new_AGEMA_signal_6627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C ( clk ), .D ( new_AGEMA_signal_6629 ), .Q ( new_AGEMA_signal_6630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C ( clk ), .D ( new_AGEMA_signal_6631 ), .Q ( new_AGEMA_signal_6632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C ( clk ), .D ( new_AGEMA_signal_6633 ), .Q ( new_AGEMA_signal_6634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C ( clk ), .D ( new_AGEMA_signal_6635 ), .Q ( new_AGEMA_signal_6636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C ( clk ), .D ( new_AGEMA_signal_6637 ), .Q ( new_AGEMA_signal_6638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C ( clk ), .D ( new_AGEMA_signal_6641 ), .Q ( new_AGEMA_signal_6642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C ( clk ), .D ( new_AGEMA_signal_6645 ), .Q ( new_AGEMA_signal_6646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C ( clk ), .D ( new_AGEMA_signal_6648 ), .Q ( new_AGEMA_signal_6649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C ( clk ), .D ( new_AGEMA_signal_6651 ), .Q ( new_AGEMA_signal_6652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C ( clk ), .D ( new_AGEMA_signal_6655 ), .Q ( new_AGEMA_signal_6656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C ( clk ), .D ( new_AGEMA_signal_6659 ), .Q ( new_AGEMA_signal_6660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C ( clk ), .D ( new_AGEMA_signal_6663 ), .Q ( new_AGEMA_signal_6664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C ( clk ), .D ( new_AGEMA_signal_6667 ), .Q ( new_AGEMA_signal_6668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C ( clk ), .D ( n2514 ), .Q ( new_AGEMA_signal_6669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C ( clk ), .D ( new_AGEMA_signal_1754 ), .Q ( new_AGEMA_signal_6670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C ( clk ), .D ( new_AGEMA_signal_6671 ), .Q ( new_AGEMA_signal_6672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C ( clk ), .D ( new_AGEMA_signal_6673 ), .Q ( new_AGEMA_signal_6674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C ( clk ), .D ( new_AGEMA_signal_6675 ), .Q ( new_AGEMA_signal_6676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C ( clk ), .D ( new_AGEMA_signal_6677 ), .Q ( new_AGEMA_signal_6678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C ( clk ), .D ( new_AGEMA_signal_6681 ), .Q ( new_AGEMA_signal_6682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C ( clk ), .D ( new_AGEMA_signal_6685 ), .Q ( new_AGEMA_signal_6686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C ( clk ), .D ( new_AGEMA_signal_6687 ), .Q ( new_AGEMA_signal_6688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C ( clk ), .D ( new_AGEMA_signal_6689 ), .Q ( new_AGEMA_signal_6690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C ( clk ), .D ( new_AGEMA_signal_6692 ), .Q ( new_AGEMA_signal_6693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C ( clk ), .D ( new_AGEMA_signal_6696 ), .Q ( new_AGEMA_signal_6697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C ( clk ), .D ( new_AGEMA_signal_6702 ), .Q ( new_AGEMA_signal_6703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C ( clk ), .D ( new_AGEMA_signal_6708 ), .Q ( new_AGEMA_signal_6709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C ( clk ), .D ( new_AGEMA_signal_6715 ), .Q ( new_AGEMA_signal_6716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C ( clk ), .D ( new_AGEMA_signal_6722 ), .Q ( new_AGEMA_signal_6723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C ( clk ), .D ( new_AGEMA_signal_6726 ), .Q ( new_AGEMA_signal_6727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C ( clk ), .D ( new_AGEMA_signal_6730 ), .Q ( new_AGEMA_signal_6731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C ( clk ), .D ( new_AGEMA_signal_6737 ), .Q ( new_AGEMA_signal_6738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C ( clk ), .D ( new_AGEMA_signal_6744 ), .Q ( new_AGEMA_signal_6745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C ( clk ), .D ( new_AGEMA_signal_6748 ), .Q ( new_AGEMA_signal_6749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C ( clk ), .D ( new_AGEMA_signal_6752 ), .Q ( new_AGEMA_signal_6753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C ( clk ), .D ( new_AGEMA_signal_6756 ), .Q ( new_AGEMA_signal_6757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C ( clk ), .D ( new_AGEMA_signal_6760 ), .Q ( new_AGEMA_signal_6761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C ( clk ), .D ( new_AGEMA_signal_6773 ), .Q ( new_AGEMA_signal_6774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C ( clk ), .D ( new_AGEMA_signal_6781 ), .Q ( new_AGEMA_signal_6782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C ( clk ), .D ( new_AGEMA_signal_6795 ), .Q ( new_AGEMA_signal_6796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C ( clk ), .D ( new_AGEMA_signal_6803 ), .Q ( new_AGEMA_signal_6804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C ( clk ), .D ( new_AGEMA_signal_6808 ), .Q ( new_AGEMA_signal_6809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C ( clk ), .D ( new_AGEMA_signal_6813 ), .Q ( new_AGEMA_signal_6814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C ( clk ), .D ( new_AGEMA_signal_6821 ), .Q ( new_AGEMA_signal_6822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C ( clk ), .D ( new_AGEMA_signal_6825 ), .Q ( new_AGEMA_signal_6826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C ( clk ), .D ( new_AGEMA_signal_6844 ), .Q ( new_AGEMA_signal_6845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C ( clk ), .D ( new_AGEMA_signal_6852 ), .Q ( new_AGEMA_signal_6853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C ( clk ), .D ( new_AGEMA_signal_6857 ), .Q ( new_AGEMA_signal_6858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C ( clk ), .D ( new_AGEMA_signal_6862 ), .Q ( new_AGEMA_signal_6863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C ( clk ), .D ( new_AGEMA_signal_6871 ), .Q ( new_AGEMA_signal_6872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C ( clk ), .D ( new_AGEMA_signal_6880 ), .Q ( new_AGEMA_signal_6881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C ( clk ), .D ( n2671 ), .Q ( new_AGEMA_signal_6889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C ( clk ), .D ( new_AGEMA_signal_1791 ), .Q ( new_AGEMA_signal_6893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C ( clk ), .D ( new_AGEMA_signal_6921 ), .Q ( new_AGEMA_signal_6922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C ( clk ), .D ( new_AGEMA_signal_6931 ), .Q ( new_AGEMA_signal_6932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C ( clk ), .D ( n2380 ), .Q ( new_AGEMA_signal_6945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C ( clk ), .D ( new_AGEMA_signal_1786 ), .Q ( new_AGEMA_signal_6951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C ( clk ), .D ( n2382 ), .Q ( new_AGEMA_signal_6957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C ( clk ), .D ( new_AGEMA_signal_1785 ), .Q ( new_AGEMA_signal_6964 ) ) ;

    /* cells in depth 10 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2117 ( .a ({new_AGEMA_signal_6598, new_AGEMA_signal_6595}), .b ({new_AGEMA_signal_1799, n1989}), .clk ( clk ), .r ({Fresh[3271], Fresh[3270], Fresh[3269], Fresh[3268]}), .c ({new_AGEMA_signal_1821, n2000}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2181 ( .a ({new_AGEMA_signal_1773, n2038}), .b ({new_AGEMA_signal_6602, new_AGEMA_signal_6600}), .clk ( clk ), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272]}), .c ({new_AGEMA_signal_1801, n2113}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2231 ( .a ({new_AGEMA_signal_1803, n2079}), .b ({new_AGEMA_signal_6608, new_AGEMA_signal_6605}), .clk ( clk ), .r ({Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_1822, n2109}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2264 ( .a ({new_AGEMA_signal_6618, new_AGEMA_signal_6613}), .b ({new_AGEMA_signal_1804, n2104}), .clk ( clk ), .r ({Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280]}), .c ({new_AGEMA_signal_1823, n2107}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2290 ( .a ({new_AGEMA_signal_6624, new_AGEMA_signal_6621}), .b ({new_AGEMA_signal_1805, n2127}), .clk ( clk ), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284]}), .c ({new_AGEMA_signal_1824, n2212}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2316 ( .a ({new_AGEMA_signal_6630, new_AGEMA_signal_6627}), .b ({new_AGEMA_signal_1806, n2147}), .clk ( clk ), .r ({Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_1825, n2149}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2366 ( .a ({new_AGEMA_signal_1808, n2199}), .b ({new_AGEMA_signal_6634, new_AGEMA_signal_6632}), .clk ( clk ), .r ({Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292]}), .c ({new_AGEMA_signal_1826, n2206}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2421 ( .a ({new_AGEMA_signal_6638, new_AGEMA_signal_6636}), .b ({new_AGEMA_signal_1809, n2257}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296]}), .c ({new_AGEMA_signal_1827, n2310}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2447 ( .a ({new_AGEMA_signal_1810, n2281}), .b ({new_AGEMA_signal_6646, new_AGEMA_signal_6642}), .clk ( clk ), .r ({Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_1828, n2308}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2476 ( .a ({new_AGEMA_signal_6652, new_AGEMA_signal_6649}), .b ({new_AGEMA_signal_1811, n2305}), .clk ( clk ), .r ({Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304]}), .c ({new_AGEMA_signal_1829, n2307}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2533 ( .a ({new_AGEMA_signal_6660, new_AGEMA_signal_6656}), .b ({new_AGEMA_signal_1812, n2368}), .clk ( clk ), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308]}), .c ({new_AGEMA_signal_1830, n2370}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2611 ( .a ({new_AGEMA_signal_1814, n2457}), .b ({new_AGEMA_signal_6668, new_AGEMA_signal_6664}), .clk ( clk ), .r ({Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_1831, n2530}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2660 ( .a ({new_AGEMA_signal_6670, new_AGEMA_signal_6669}), .b ({new_AGEMA_signal_1815, n2513}), .clk ( clk ), .r ({Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316]}), .c ({new_AGEMA_signal_1832, n2515}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2718 ( .a ({new_AGEMA_signal_6674, new_AGEMA_signal_6672}), .b ({new_AGEMA_signal_1816, n2592}), .clk ( clk ), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320]}), .c ({new_AGEMA_signal_1833, n2639}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2749 ( .a ({new_AGEMA_signal_1793, n2637}), .b ({new_AGEMA_signal_6678, new_AGEMA_signal_6676}), .clk ( clk ), .r ({Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_1817, n2638}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2788 ( .a ({new_AGEMA_signal_6686, new_AGEMA_signal_6682}), .b ({new_AGEMA_signal_1819, n2705}), .clk ( clk ), .r ({Fresh[3331], Fresh[3330], Fresh[3329], Fresh[3328]}), .c ({new_AGEMA_signal_1834, n2832}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2842 ( .a ({new_AGEMA_signal_6690, new_AGEMA_signal_6688}), .b ({new_AGEMA_signal_1796, n2805}), .clk ( clk ), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332]}), .c ({new_AGEMA_signal_1820, n2807}) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C ( clk ), .D ( new_AGEMA_signal_6693 ), .Q ( new_AGEMA_signal_6694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C ( clk ), .D ( new_AGEMA_signal_6697 ), .Q ( new_AGEMA_signal_6698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C ( clk ), .D ( new_AGEMA_signal_6703 ), .Q ( new_AGEMA_signal_6704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C ( clk ), .D ( new_AGEMA_signal_6709 ), .Q ( new_AGEMA_signal_6710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C ( clk ), .D ( new_AGEMA_signal_6716 ), .Q ( new_AGEMA_signal_6717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C ( clk ), .D ( new_AGEMA_signal_6723 ), .Q ( new_AGEMA_signal_6724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C ( clk ), .D ( new_AGEMA_signal_6727 ), .Q ( new_AGEMA_signal_6728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C ( clk ), .D ( new_AGEMA_signal_6731 ), .Q ( new_AGEMA_signal_6732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C ( clk ), .D ( new_AGEMA_signal_6738 ), .Q ( new_AGEMA_signal_6739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C ( clk ), .D ( new_AGEMA_signal_6745 ), .Q ( new_AGEMA_signal_6746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C ( clk ), .D ( new_AGEMA_signal_6749 ), .Q ( new_AGEMA_signal_6750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C ( clk ), .D ( new_AGEMA_signal_6753 ), .Q ( new_AGEMA_signal_6754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C ( clk ), .D ( new_AGEMA_signal_6757 ), .Q ( new_AGEMA_signal_6758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C ( clk ), .D ( new_AGEMA_signal_6761 ), .Q ( new_AGEMA_signal_6762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C ( clk ), .D ( n2002 ), .Q ( new_AGEMA_signal_6763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C ( clk ), .D ( new_AGEMA_signal_1798 ), .Q ( new_AGEMA_signal_6765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C ( clk ), .D ( new_AGEMA_signal_6774 ), .Q ( new_AGEMA_signal_6775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C ( clk ), .D ( new_AGEMA_signal_6782 ), .Q ( new_AGEMA_signal_6783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C ( clk ), .D ( n2208 ), .Q ( new_AGEMA_signal_6785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C ( clk ), .D ( new_AGEMA_signal_1807 ), .Q ( new_AGEMA_signal_6787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C ( clk ), .D ( new_AGEMA_signal_6796 ), .Q ( new_AGEMA_signal_6797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C ( clk ), .D ( new_AGEMA_signal_6804 ), .Q ( new_AGEMA_signal_6805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C ( clk ), .D ( new_AGEMA_signal_6809 ), .Q ( new_AGEMA_signal_6810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C ( clk ), .D ( new_AGEMA_signal_6814 ), .Q ( new_AGEMA_signal_6815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C ( clk ), .D ( n2668 ), .Q ( new_AGEMA_signal_6817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C ( clk ), .D ( new_AGEMA_signal_1818 ), .Q ( new_AGEMA_signal_6819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C ( clk ), .D ( new_AGEMA_signal_6822 ), .Q ( new_AGEMA_signal_6823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C ( clk ), .D ( new_AGEMA_signal_6826 ), .Q ( new_AGEMA_signal_6827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C ( clk ), .D ( n2016 ), .Q ( new_AGEMA_signal_6829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C ( clk ), .D ( new_AGEMA_signal_1800 ), .Q ( new_AGEMA_signal_6832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C ( clk ), .D ( n2111 ), .Q ( new_AGEMA_signal_6835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C ( clk ), .D ( new_AGEMA_signal_1802 ), .Q ( new_AGEMA_signal_6838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C ( clk ), .D ( new_AGEMA_signal_6845 ), .Q ( new_AGEMA_signal_6846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C ( clk ), .D ( new_AGEMA_signal_6853 ), .Q ( new_AGEMA_signal_6854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C ( clk ), .D ( new_AGEMA_signal_6858 ), .Q ( new_AGEMA_signal_6859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C ( clk ), .D ( new_AGEMA_signal_6863 ), .Q ( new_AGEMA_signal_6864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C ( clk ), .D ( new_AGEMA_signal_6872 ), .Q ( new_AGEMA_signal_6873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C ( clk ), .D ( new_AGEMA_signal_6881 ), .Q ( new_AGEMA_signal_6882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C ( clk ), .D ( new_AGEMA_signal_6889 ), .Q ( new_AGEMA_signal_6890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C ( clk ), .D ( new_AGEMA_signal_6893 ), .Q ( new_AGEMA_signal_6894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C ( clk ), .D ( n2019 ), .Q ( new_AGEMA_signal_6901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C ( clk ), .D ( new_AGEMA_signal_1797 ), .Q ( new_AGEMA_signal_6905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C ( clk ), .D ( new_AGEMA_signal_6922 ), .Q ( new_AGEMA_signal_6923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C ( clk ), .D ( new_AGEMA_signal_6932 ), .Q ( new_AGEMA_signal_6933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C ( clk ), .D ( new_AGEMA_signal_6945 ), .Q ( new_AGEMA_signal_6946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C ( clk ), .D ( new_AGEMA_signal_6951 ), .Q ( new_AGEMA_signal_6952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C ( clk ), .D ( new_AGEMA_signal_6957 ), .Q ( new_AGEMA_signal_6958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C ( clk ), .D ( new_AGEMA_signal_6964 ), .Q ( new_AGEMA_signal_6965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C ( clk ), .D ( n2426 ), .Q ( new_AGEMA_signal_6971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C ( clk ), .D ( new_AGEMA_signal_1813 ), .Q ( new_AGEMA_signal_6978 ) ) ;

    /* cells in depth 11 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2129 ( .a ({new_AGEMA_signal_1821, n2000}), .b ({new_AGEMA_signal_6698, new_AGEMA_signal_6694}), .clk ( clk ), .r ({Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_1836, n2001}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2267 ( .a ({new_AGEMA_signal_1823, n2107}), .b ({new_AGEMA_signal_6710, new_AGEMA_signal_6704}), .clk ( clk ), .r ({Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340]}), .c ({new_AGEMA_signal_1837, n2108}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2317 ( .a ({new_AGEMA_signal_6724, new_AGEMA_signal_6717}), .b ({new_AGEMA_signal_1825, n2149}), .clk ( clk ), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344]}), .c ({new_AGEMA_signal_1838, n2153}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2374 ( .a ({new_AGEMA_signal_1826, n2206}), .b ({new_AGEMA_signal_6732, new_AGEMA_signal_6728}), .clk ( clk ), .r ({Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_1839, n2207}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2477 ( .a ({new_AGEMA_signal_1828, n2308}), .b ({new_AGEMA_signal_1829, n2307}), .clk ( clk ), .r ({Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352]}), .c ({new_AGEMA_signal_1840, n2309}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2535 ( .a ({new_AGEMA_signal_1830, n2370}), .b ({new_AGEMA_signal_6746, new_AGEMA_signal_6739}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356]}), .c ({new_AGEMA_signal_1841, n2373}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2661 ( .a ({new_AGEMA_signal_6754, new_AGEMA_signal_6750}), .b ({new_AGEMA_signal_1832, n2515}), .clk ( clk ), .r ({Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({new_AGEMA_signal_1842, n2528}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2750 ( .a ({new_AGEMA_signal_1833, n2639}), .b ({new_AGEMA_signal_1817, n2638}), .clk ( clk ), .r ({Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364]}), .c ({new_AGEMA_signal_1843, n2669}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2843 ( .a ({new_AGEMA_signal_6762, new_AGEMA_signal_6758}), .b ({new_AGEMA_signal_1820, n2807}), .clk ( clk ), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368]}), .c ({new_AGEMA_signal_1835, n2830}) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C ( clk ), .D ( new_AGEMA_signal_6763 ), .Q ( new_AGEMA_signal_6764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C ( clk ), .D ( new_AGEMA_signal_6765 ), .Q ( new_AGEMA_signal_6766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C ( clk ), .D ( n2109 ), .Q ( new_AGEMA_signal_6767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_6768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C ( clk ), .D ( new_AGEMA_signal_6775 ), .Q ( new_AGEMA_signal_6776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C ( clk ), .D ( new_AGEMA_signal_6783 ), .Q ( new_AGEMA_signal_6784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C ( clk ), .D ( new_AGEMA_signal_6785 ), .Q ( new_AGEMA_signal_6786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C ( clk ), .D ( new_AGEMA_signal_6787 ), .Q ( new_AGEMA_signal_6788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C ( clk ), .D ( n2310 ), .Q ( new_AGEMA_signal_6789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C ( clk ), .D ( new_AGEMA_signal_1827 ), .Q ( new_AGEMA_signal_6790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C ( clk ), .D ( new_AGEMA_signal_6797 ), .Q ( new_AGEMA_signal_6798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C ( clk ), .D ( new_AGEMA_signal_6805 ), .Q ( new_AGEMA_signal_6806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C ( clk ), .D ( new_AGEMA_signal_6810 ), .Q ( new_AGEMA_signal_6811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C ( clk ), .D ( new_AGEMA_signal_6815 ), .Q ( new_AGEMA_signal_6816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C ( clk ), .D ( new_AGEMA_signal_6817 ), .Q ( new_AGEMA_signal_6818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C ( clk ), .D ( new_AGEMA_signal_6819 ), .Q ( new_AGEMA_signal_6820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C ( clk ), .D ( new_AGEMA_signal_6823 ), .Q ( new_AGEMA_signal_6824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C ( clk ), .D ( new_AGEMA_signal_6827 ), .Q ( new_AGEMA_signal_6828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C ( clk ), .D ( new_AGEMA_signal_6829 ), .Q ( new_AGEMA_signal_6830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C ( clk ), .D ( new_AGEMA_signal_6832 ), .Q ( new_AGEMA_signal_6833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C ( clk ), .D ( new_AGEMA_signal_6835 ), .Q ( new_AGEMA_signal_6836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C ( clk ), .D ( new_AGEMA_signal_6838 ), .Q ( new_AGEMA_signal_6839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C ( clk ), .D ( new_AGEMA_signal_6846 ), .Q ( new_AGEMA_signal_6847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C ( clk ), .D ( new_AGEMA_signal_6854 ), .Q ( new_AGEMA_signal_6855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C ( clk ), .D ( new_AGEMA_signal_6859 ), .Q ( new_AGEMA_signal_6860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C ( clk ), .D ( new_AGEMA_signal_6864 ), .Q ( new_AGEMA_signal_6865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C ( clk ), .D ( new_AGEMA_signal_6873 ), .Q ( new_AGEMA_signal_6874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C ( clk ), .D ( new_AGEMA_signal_6882 ), .Q ( new_AGEMA_signal_6883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C ( clk ), .D ( n2530 ), .Q ( new_AGEMA_signal_6885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C ( clk ), .D ( new_AGEMA_signal_1831 ), .Q ( new_AGEMA_signal_6887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C ( clk ), .D ( new_AGEMA_signal_6890 ), .Q ( new_AGEMA_signal_6891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C ( clk ), .D ( new_AGEMA_signal_6894 ), .Q ( new_AGEMA_signal_6895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C ( clk ), .D ( n2832 ), .Q ( new_AGEMA_signal_6897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C ( clk ), .D ( new_AGEMA_signal_1834 ), .Q ( new_AGEMA_signal_6899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C ( clk ), .D ( new_AGEMA_signal_6901 ), .Q ( new_AGEMA_signal_6902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C ( clk ), .D ( new_AGEMA_signal_6905 ), .Q ( new_AGEMA_signal_6906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C ( clk ), .D ( n2113 ), .Q ( new_AGEMA_signal_6909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C ( clk ), .D ( new_AGEMA_signal_1801 ), .Q ( new_AGEMA_signal_6912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C ( clk ), .D ( new_AGEMA_signal_6923 ), .Q ( new_AGEMA_signal_6924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C ( clk ), .D ( new_AGEMA_signal_6933 ), .Q ( new_AGEMA_signal_6934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C ( clk ), .D ( n2212 ), .Q ( new_AGEMA_signal_6937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C ( clk ), .D ( new_AGEMA_signal_1824 ), .Q ( new_AGEMA_signal_6941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C ( clk ), .D ( new_AGEMA_signal_6946 ), .Q ( new_AGEMA_signal_6947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C ( clk ), .D ( new_AGEMA_signal_6952 ), .Q ( new_AGEMA_signal_6953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C ( clk ), .D ( new_AGEMA_signal_6958 ), .Q ( new_AGEMA_signal_6959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C ( clk ), .D ( new_AGEMA_signal_6965 ), .Q ( new_AGEMA_signal_6966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C ( clk ), .D ( new_AGEMA_signal_6971 ), .Q ( new_AGEMA_signal_6972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C ( clk ), .D ( new_AGEMA_signal_6978 ), .Q ( new_AGEMA_signal_6979 ) ) ;

    /* cells in depth 12 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2130 ( .a ({new_AGEMA_signal_6766, new_AGEMA_signal_6764}), .b ({new_AGEMA_signal_1836, n2001}), .clk ( clk ), .r ({Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({new_AGEMA_signal_1845, n2017}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2268 ( .a ({new_AGEMA_signal_6768, new_AGEMA_signal_6767}), .b ({new_AGEMA_signal_1837, n2108}), .clk ( clk ), .r ({Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376]}), .c ({new_AGEMA_signal_1846, n2110}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2319 ( .a ({new_AGEMA_signal_1838, n2153}), .b ({new_AGEMA_signal_6784, new_AGEMA_signal_6776}), .clk ( clk ), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380]}), .c ({new_AGEMA_signal_1847, n2154}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2375 ( .a ({new_AGEMA_signal_6788, new_AGEMA_signal_6786}), .b ({new_AGEMA_signal_1839, n2207}), .clk ( clk ), .r ({Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({new_AGEMA_signal_1848, n2209}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2478 ( .a ({new_AGEMA_signal_6790, new_AGEMA_signal_6789}), .b ({new_AGEMA_signal_1840, n2309}), .clk ( clk ), .r ({Fresh[3391], Fresh[3390], Fresh[3389], Fresh[3388]}), .c ({new_AGEMA_signal_1849, n2311}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2537 ( .a ({new_AGEMA_signal_1841, n2373}), .b ({new_AGEMA_signal_6806, new_AGEMA_signal_6798}), .clk ( clk ), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392]}), .c ({new_AGEMA_signal_1850, n2374}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2672 ( .a ({new_AGEMA_signal_1842, n2528}), .b ({new_AGEMA_signal_6816, new_AGEMA_signal_6811}), .clk ( clk ), .r ({Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({new_AGEMA_signal_1851, n2529}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2768 ( .a ({new_AGEMA_signal_1843, n2669}), .b ({new_AGEMA_signal_6820, new_AGEMA_signal_6818}), .clk ( clk ), .r ({Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400]}), .c ({new_AGEMA_signal_1852, n2670}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2854 ( .a ({new_AGEMA_signal_1835, n2830}), .b ({new_AGEMA_signal_6828, new_AGEMA_signal_6824}), .clk ( clk ), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404]}), .c ({new_AGEMA_signal_1844, n2831}) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C ( clk ), .D ( new_AGEMA_signal_6830 ), .Q ( new_AGEMA_signal_6831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C ( clk ), .D ( new_AGEMA_signal_6833 ), .Q ( new_AGEMA_signal_6834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C ( clk ), .D ( new_AGEMA_signal_6836 ), .Q ( new_AGEMA_signal_6837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C ( clk ), .D ( new_AGEMA_signal_6839 ), .Q ( new_AGEMA_signal_6840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C ( clk ), .D ( new_AGEMA_signal_6847 ), .Q ( new_AGEMA_signal_6848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C ( clk ), .D ( new_AGEMA_signal_6855 ), .Q ( new_AGEMA_signal_6856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C ( clk ), .D ( new_AGEMA_signal_6860 ), .Q ( new_AGEMA_signal_6861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C ( clk ), .D ( new_AGEMA_signal_6865 ), .Q ( new_AGEMA_signal_6866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C ( clk ), .D ( new_AGEMA_signal_6874 ), .Q ( new_AGEMA_signal_6875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C ( clk ), .D ( new_AGEMA_signal_6883 ), .Q ( new_AGEMA_signal_6884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C ( clk ), .D ( new_AGEMA_signal_6885 ), .Q ( new_AGEMA_signal_6886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C ( clk ), .D ( new_AGEMA_signal_6887 ), .Q ( new_AGEMA_signal_6888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C ( clk ), .D ( new_AGEMA_signal_6891 ), .Q ( new_AGEMA_signal_6892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C ( clk ), .D ( new_AGEMA_signal_6895 ), .Q ( new_AGEMA_signal_6896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C ( clk ), .D ( new_AGEMA_signal_6897 ), .Q ( new_AGEMA_signal_6898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C ( clk ), .D ( new_AGEMA_signal_6899 ), .Q ( new_AGEMA_signal_6900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C ( clk ), .D ( new_AGEMA_signal_6902 ), .Q ( new_AGEMA_signal_6903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C ( clk ), .D ( new_AGEMA_signal_6906 ), .Q ( new_AGEMA_signal_6907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C ( clk ), .D ( new_AGEMA_signal_6909 ), .Q ( new_AGEMA_signal_6910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C ( clk ), .D ( new_AGEMA_signal_6912 ), .Q ( new_AGEMA_signal_6913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C ( clk ), .D ( new_AGEMA_signal_6924 ), .Q ( new_AGEMA_signal_6925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C ( clk ), .D ( new_AGEMA_signal_6934 ), .Q ( new_AGEMA_signal_6935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C ( clk ), .D ( new_AGEMA_signal_6937 ), .Q ( new_AGEMA_signal_6938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C ( clk ), .D ( new_AGEMA_signal_6941 ), .Q ( new_AGEMA_signal_6942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C ( clk ), .D ( new_AGEMA_signal_6947 ), .Q ( new_AGEMA_signal_6948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C ( clk ), .D ( new_AGEMA_signal_6953 ), .Q ( new_AGEMA_signal_6954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C ( clk ), .D ( new_AGEMA_signal_6959 ), .Q ( new_AGEMA_signal_6960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C ( clk ), .D ( new_AGEMA_signal_6966 ), .Q ( new_AGEMA_signal_6967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C ( clk ), .D ( new_AGEMA_signal_6972 ), .Q ( new_AGEMA_signal_6973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C ( clk ), .D ( new_AGEMA_signal_6979 ), .Q ( new_AGEMA_signal_6980 ) ) ;

    /* cells in depth 13 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2155 ( .a ({new_AGEMA_signal_1845, n2017}), .b ({new_AGEMA_signal_6834, new_AGEMA_signal_6831}), .clk ( clk ), .r ({Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({new_AGEMA_signal_1854, n2018}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2269 ( .a ({new_AGEMA_signal_6840, new_AGEMA_signal_6837}), .b ({new_AGEMA_signal_1846, n2110}), .clk ( clk ), .r ({Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412]}), .c ({new_AGEMA_signal_1855, n2112}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2320 ( .a ({new_AGEMA_signal_6856, new_AGEMA_signal_6848}), .b ({new_AGEMA_signal_1847, n2154}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416]}), .c ({new_AGEMA_signal_1856, n2210}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2479 ( .a ({new_AGEMA_signal_6866, new_AGEMA_signal_6861}), .b ({new_AGEMA_signal_1849, n2311}), .clk ( clk ), .r ({Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({new_AGEMA_signal_1857, N470}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2538 ( .a ({new_AGEMA_signal_6884, new_AGEMA_signal_6875}), .b ({new_AGEMA_signal_1850, n2374}), .clk ( clk ), .r ({Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424]}), .c ({new_AGEMA_signal_1858, n2378}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2673 ( .a ({new_AGEMA_signal_6888, new_AGEMA_signal_6886}), .b ({new_AGEMA_signal_1851, n2529}), .clk ( clk ), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428]}), .c ({new_AGEMA_signal_1859, N639}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2769 ( .a ({new_AGEMA_signal_6896, new_AGEMA_signal_6892}), .b ({new_AGEMA_signal_1852, n2670}), .clk ( clk ), .r ({Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({new_AGEMA_signal_1860, N723}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2855 ( .a ({new_AGEMA_signal_6900, new_AGEMA_signal_6898}), .b ({new_AGEMA_signal_1844, n2831}), .clk ( clk ), .r ({Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436]}), .c ({new_AGEMA_signal_1853, N789}) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C ( clk ), .D ( new_AGEMA_signal_6903 ), .Q ( new_AGEMA_signal_6904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C ( clk ), .D ( new_AGEMA_signal_6907 ), .Q ( new_AGEMA_signal_6908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C ( clk ), .D ( new_AGEMA_signal_6910 ), .Q ( new_AGEMA_signal_6911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C ( clk ), .D ( new_AGEMA_signal_6913 ), .Q ( new_AGEMA_signal_6914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C ( clk ), .D ( n2209 ), .Q ( new_AGEMA_signal_6915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C ( clk ), .D ( new_AGEMA_signal_1848 ), .Q ( new_AGEMA_signal_6916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C ( clk ), .D ( new_AGEMA_signal_6925 ), .Q ( new_AGEMA_signal_6926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C ( clk ), .D ( new_AGEMA_signal_6935 ), .Q ( new_AGEMA_signal_6936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C ( clk ), .D ( new_AGEMA_signal_6938 ), .Q ( new_AGEMA_signal_6939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C ( clk ), .D ( new_AGEMA_signal_6942 ), .Q ( new_AGEMA_signal_6943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C ( clk ), .D ( new_AGEMA_signal_6948 ), .Q ( new_AGEMA_signal_6949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C ( clk ), .D ( new_AGEMA_signal_6954 ), .Q ( new_AGEMA_signal_6955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C ( clk ), .D ( new_AGEMA_signal_6960 ), .Q ( new_AGEMA_signal_6961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C ( clk ), .D ( new_AGEMA_signal_6967 ), .Q ( new_AGEMA_signal_6968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C ( clk ), .D ( new_AGEMA_signal_6973 ), .Q ( new_AGEMA_signal_6974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C ( clk ), .D ( new_AGEMA_signal_6980 ), .Q ( new_AGEMA_signal_6981 ) ) ;

    /* cells in depth 14 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2156 ( .a ({new_AGEMA_signal_6908, new_AGEMA_signal_6904}), .b ({new_AGEMA_signal_1854, n2018}), .clk ( clk ), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440]}), .c ({new_AGEMA_signal_1861, N169}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2270 ( .a ({new_AGEMA_signal_6914, new_AGEMA_signal_6911}), .b ({new_AGEMA_signal_1855, n2112}), .clk ( clk ), .r ({Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({new_AGEMA_signal_1862, N277}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2376 ( .a ({new_AGEMA_signal_1856, n2210}), .b ({new_AGEMA_signal_6916, new_AGEMA_signal_6915}), .clk ( clk ), .r ({Fresh[3451], Fresh[3450], Fresh[3449], Fresh[3448]}), .c ({new_AGEMA_signal_1863, n2211}) ) ;
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2540 ( .a ({new_AGEMA_signal_1858, n2378}), .b ({new_AGEMA_signal_6936, new_AGEMA_signal_6926}), .clk ( clk ), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452]}), .c ({new_AGEMA_signal_1864, n2379}) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C ( clk ), .D ( new_AGEMA_signal_6939 ), .Q ( new_AGEMA_signal_6940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C ( clk ), .D ( new_AGEMA_signal_6943 ), .Q ( new_AGEMA_signal_6944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C ( clk ), .D ( new_AGEMA_signal_6949 ), .Q ( new_AGEMA_signal_6950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C ( clk ), .D ( new_AGEMA_signal_6955 ), .Q ( new_AGEMA_signal_6956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C ( clk ), .D ( new_AGEMA_signal_6961 ), .Q ( new_AGEMA_signal_6962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C ( clk ), .D ( new_AGEMA_signal_6968 ), .Q ( new_AGEMA_signal_6969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C ( clk ), .D ( new_AGEMA_signal_6974 ), .Q ( new_AGEMA_signal_6975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C ( clk ), .D ( new_AGEMA_signal_6981 ), .Q ( new_AGEMA_signal_6982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C ( clk ), .D ( N470 ), .Q ( new_AGEMA_signal_7001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C ( clk ), .D ( new_AGEMA_signal_1857 ), .Q ( new_AGEMA_signal_7005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C ( clk ), .D ( N639 ), .Q ( new_AGEMA_signal_7009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C ( clk ), .D ( new_AGEMA_signal_1859 ), .Q ( new_AGEMA_signal_7013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C ( clk ), .D ( N723 ), .Q ( new_AGEMA_signal_7017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C ( clk ), .D ( new_AGEMA_signal_1860 ), .Q ( new_AGEMA_signal_7021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C ( clk ), .D ( N789 ), .Q ( new_AGEMA_signal_7025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_7029 ) ) ;

    /* cells in depth 15 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2377 ( .a ({new_AGEMA_signal_6944, new_AGEMA_signal_6940}), .b ({new_AGEMA_signal_1863, n2211}), .clk ( clk ), .r ({Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({new_AGEMA_signal_1865, N379}) ) ;
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2541 ( .a ({new_AGEMA_signal_6956, new_AGEMA_signal_6950}), .b ({new_AGEMA_signal_1864, n2379}), .clk ( clk ), .r ({Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460]}), .c ({new_AGEMA_signal_1866, n2381}) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C ( clk ), .D ( new_AGEMA_signal_6962 ), .Q ( new_AGEMA_signal_6963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C ( clk ), .D ( new_AGEMA_signal_6969 ), .Q ( new_AGEMA_signal_6970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C ( clk ), .D ( new_AGEMA_signal_6975 ), .Q ( new_AGEMA_signal_6976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C ( clk ), .D ( new_AGEMA_signal_6982 ), .Q ( new_AGEMA_signal_6983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C ( clk ), .D ( N169 ), .Q ( new_AGEMA_signal_6985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C ( clk ), .D ( new_AGEMA_signal_1861 ), .Q ( new_AGEMA_signal_6988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C ( clk ), .D ( N277 ), .Q ( new_AGEMA_signal_6991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C ( clk ), .D ( new_AGEMA_signal_1862 ), .Q ( new_AGEMA_signal_6994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C ( clk ), .D ( new_AGEMA_signal_7001 ), .Q ( new_AGEMA_signal_7002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C ( clk ), .D ( new_AGEMA_signal_7005 ), .Q ( new_AGEMA_signal_7006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C ( clk ), .D ( new_AGEMA_signal_7009 ), .Q ( new_AGEMA_signal_7010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C ( clk ), .D ( new_AGEMA_signal_7013 ), .Q ( new_AGEMA_signal_7014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C ( clk ), .D ( new_AGEMA_signal_7017 ), .Q ( new_AGEMA_signal_7018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C ( clk ), .D ( new_AGEMA_signal_7021 ), .Q ( new_AGEMA_signal_7022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C ( clk ), .D ( new_AGEMA_signal_7025 ), .Q ( new_AGEMA_signal_7026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C ( clk ), .D ( new_AGEMA_signal_7029 ), .Q ( new_AGEMA_signal_7030 ) ) ;

    /* cells in depth 16 */
    nor_GHPC #(.low_latency(1), .pipeline(1)) U2542 ( .a ({new_AGEMA_signal_6970, new_AGEMA_signal_6963}), .b ({new_AGEMA_signal_1866, n2381}), .clk ( clk ), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464]}), .c ({new_AGEMA_signal_1867, n2427}) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C ( clk ), .D ( new_AGEMA_signal_6976 ), .Q ( new_AGEMA_signal_6977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C ( clk ), .D ( new_AGEMA_signal_6983 ), .Q ( new_AGEMA_signal_6984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C ( clk ), .D ( new_AGEMA_signal_6985 ), .Q ( new_AGEMA_signal_6986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C ( clk ), .D ( new_AGEMA_signal_6988 ), .Q ( new_AGEMA_signal_6989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C ( clk ), .D ( new_AGEMA_signal_6991 ), .Q ( new_AGEMA_signal_6992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C ( clk ), .D ( new_AGEMA_signal_6994 ), .Q ( new_AGEMA_signal_6995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C ( clk ), .D ( N379 ), .Q ( new_AGEMA_signal_6997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_6999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C ( clk ), .D ( new_AGEMA_signal_7002 ), .Q ( new_AGEMA_signal_7003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C ( clk ), .D ( new_AGEMA_signal_7006 ), .Q ( new_AGEMA_signal_7007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C ( clk ), .D ( new_AGEMA_signal_7010 ), .Q ( new_AGEMA_signal_7011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C ( clk ), .D ( new_AGEMA_signal_7014 ), .Q ( new_AGEMA_signal_7015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C ( clk ), .D ( new_AGEMA_signal_7018 ), .Q ( new_AGEMA_signal_7019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C ( clk ), .D ( new_AGEMA_signal_7022 ), .Q ( new_AGEMA_signal_7023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C ( clk ), .D ( new_AGEMA_signal_7026 ), .Q ( new_AGEMA_signal_7027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C ( clk ), .D ( new_AGEMA_signal_7030 ), .Q ( new_AGEMA_signal_7031 ) ) ;

    /* cells in depth 17 */
    nand_GHPC #(.low_latency(1), .pipeline(1)) U2584 ( .a ({new_AGEMA_signal_1867, n2427}), .b ({new_AGEMA_signal_6984, new_AGEMA_signal_6977}), .clk ( clk ), .r ({Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({new_AGEMA_signal_1868, N563}) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C ( clk ), .D ( new_AGEMA_signal_6986 ), .Q ( new_AGEMA_signal_6987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C ( clk ), .D ( new_AGEMA_signal_6989 ), .Q ( new_AGEMA_signal_6990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C ( clk ), .D ( new_AGEMA_signal_6992 ), .Q ( new_AGEMA_signal_6993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C ( clk ), .D ( new_AGEMA_signal_6995 ), .Q ( new_AGEMA_signal_6996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C ( clk ), .D ( new_AGEMA_signal_6997 ), .Q ( new_AGEMA_signal_6998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C ( clk ), .D ( new_AGEMA_signal_6999 ), .Q ( new_AGEMA_signal_7000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C ( clk ), .D ( new_AGEMA_signal_7003 ), .Q ( new_AGEMA_signal_7004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C ( clk ), .D ( new_AGEMA_signal_7007 ), .Q ( new_AGEMA_signal_7008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C ( clk ), .D ( new_AGEMA_signal_7011 ), .Q ( new_AGEMA_signal_7012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C ( clk ), .D ( new_AGEMA_signal_7015 ), .Q ( new_AGEMA_signal_7016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C ( clk ), .D ( new_AGEMA_signal_7019 ), .Q ( new_AGEMA_signal_7020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C ( clk ), .D ( new_AGEMA_signal_7023 ), .Q ( new_AGEMA_signal_7024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C ( clk ), .D ( new_AGEMA_signal_7027 ), .Q ( new_AGEMA_signal_7028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C ( clk ), .D ( new_AGEMA_signal_7031 ), .Q ( new_AGEMA_signal_7032 ) ) ;

    /* register cells */
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_6990, new_AGEMA_signal_6987}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_6996, new_AGEMA_signal_6993}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_7000, new_AGEMA_signal_6998}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_7008, new_AGEMA_signal_7004}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_1868, N563}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_7016, new_AGEMA_signal_7012}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_7024, new_AGEMA_signal_7020}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_7032, new_AGEMA_signal_7028}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
