/* modified netlist. Source: module AES in file /AES_round-based/AGEMA/AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_AIG_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] plaintext_s1 ;
    input [679:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_423 ;
    wire signal_425 ;
    wire signal_427 ;
    wire signal_429 ;
    wire signal_431 ;
    wire signal_433 ;
    wire signal_435 ;
    wire signal_437 ;
    wire signal_439 ;
    wire signal_441 ;
    wire signal_443 ;
    wire signal_445 ;
    wire signal_447 ;
    wire signal_449 ;
    wire signal_451 ;
    wire signal_453 ;
    wire signal_455 ;
    wire signal_457 ;
    wire signal_459 ;
    wire signal_461 ;
    wire signal_463 ;
    wire signal_465 ;
    wire signal_467 ;
    wire signal_469 ;
    wire signal_471 ;
    wire signal_473 ;
    wire signal_475 ;
    wire signal_477 ;
    wire signal_479 ;
    wire signal_481 ;
    wire signal_483 ;
    wire signal_485 ;
    wire signal_487 ;
    wire signal_489 ;
    wire signal_491 ;
    wire signal_493 ;
    wire signal_495 ;
    wire signal_497 ;
    wire signal_499 ;
    wire signal_501 ;
    wire signal_503 ;
    wire signal_505 ;
    wire signal_507 ;
    wire signal_509 ;
    wire signal_511 ;
    wire signal_513 ;
    wire signal_515 ;
    wire signal_517 ;
    wire signal_519 ;
    wire signal_521 ;
    wire signal_523 ;
    wire signal_525 ;
    wire signal_527 ;
    wire signal_529 ;
    wire signal_531 ;
    wire signal_533 ;
    wire signal_535 ;
    wire signal_537 ;
    wire signal_539 ;
    wire signal_541 ;
    wire signal_543 ;
    wire signal_545 ;
    wire signal_547 ;
    wire signal_549 ;
    wire signal_551 ;
    wire signal_553 ;
    wire signal_555 ;
    wire signal_557 ;
    wire signal_559 ;
    wire signal_561 ;
    wire signal_563 ;
    wire signal_565 ;
    wire signal_567 ;
    wire signal_569 ;
    wire signal_571 ;
    wire signal_573 ;
    wire signal_575 ;
    wire signal_577 ;
    wire signal_579 ;
    wire signal_581 ;
    wire signal_583 ;
    wire signal_585 ;
    wire signal_587 ;
    wire signal_589 ;
    wire signal_591 ;
    wire signal_593 ;
    wire signal_595 ;
    wire signal_597 ;
    wire signal_599 ;
    wire signal_601 ;
    wire signal_603 ;
    wire signal_605 ;
    wire signal_607 ;
    wire signal_609 ;
    wire signal_611 ;
    wire signal_613 ;
    wire signal_615 ;
    wire signal_617 ;
    wire signal_619 ;
    wire signal_621 ;
    wire signal_623 ;
    wire signal_625 ;
    wire signal_627 ;
    wire signal_629 ;
    wire signal_631 ;
    wire signal_633 ;
    wire signal_635 ;
    wire signal_637 ;
    wire signal_639 ;
    wire signal_641 ;
    wire signal_643 ;
    wire signal_645 ;
    wire signal_647 ;
    wire signal_649 ;
    wire signal_651 ;
    wire signal_653 ;
    wire signal_655 ;
    wire signal_657 ;
    wire signal_659 ;
    wire signal_661 ;
    wire signal_663 ;
    wire signal_665 ;
    wire signal_667 ;
    wire signal_669 ;
    wire signal_671 ;
    wire signal_673 ;
    wire signal_675 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3043 ;
    wire signal_3045 ;
    wire signal_3047 ;
    wire signal_3049 ;
    wire signal_3051 ;
    wire signal_3053 ;
    wire signal_3055 ;
    wire signal_3057 ;
    wire signal_3059 ;
    wire signal_3061 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3079 ;
    wire signal_3081 ;
    wire signal_3083 ;
    wire signal_3085 ;
    wire signal_3087 ;
    wire signal_3089 ;
    wire signal_3091 ;
    wire signal_3093 ;
    wire signal_3095 ;
    wire signal_3097 ;
    wire signal_3099 ;
    wire signal_3101 ;
    wire signal_3103 ;
    wire signal_3105 ;
    wire signal_3107 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3874 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3882 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3890 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3898 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3906 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3914 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3922 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3930 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3938 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3946 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3954 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3962 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3970 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3978 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3986 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4394 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4402 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4410 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4418 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4426 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4434 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4442 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4450 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4458 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4466 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4474 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4482 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4490 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4498 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4506 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4514 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;
    wire signal_7973 ;
    wire signal_7974 ;
    wire signal_7975 ;
    wire signal_7976 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_8256 ;
    wire signal_8257 ;
    wire signal_8258 ;
    wire signal_8259 ;
    wire signal_8260 ;
    wire signal_8261 ;
    wire signal_8262 ;
    wire signal_8263 ;
    wire signal_8264 ;
    wire signal_8265 ;
    wire signal_8266 ;
    wire signal_8267 ;
    wire signal_8268 ;
    wire signal_8269 ;
    wire signal_8270 ;
    wire signal_8271 ;
    wire signal_8272 ;
    wire signal_8273 ;
    wire signal_8274 ;
    wire signal_8275 ;
    wire signal_8276 ;
    wire signal_8277 ;
    wire signal_8278 ;
    wire signal_8279 ;
    wire signal_8280 ;
    wire signal_8281 ;
    wire signal_8282 ;
    wire signal_8283 ;
    wire signal_8284 ;
    wire signal_8285 ;
    wire signal_8286 ;
    wire signal_8287 ;
    wire signal_8288 ;
    wire signal_8289 ;
    wire signal_8290 ;
    wire signal_8291 ;
    wire signal_8292 ;
    wire signal_8293 ;
    wire signal_8294 ;
    wire signal_8295 ;
    wire signal_8296 ;
    wire signal_8297 ;
    wire signal_8298 ;
    wire signal_8299 ;
    wire signal_8300 ;
    wire signal_8301 ;
    wire signal_8302 ;
    wire signal_8303 ;
    wire signal_8304 ;
    wire signal_8305 ;
    wire signal_8306 ;
    wire signal_8307 ;
    wire signal_8308 ;
    wire signal_8309 ;
    wire signal_8310 ;
    wire signal_8311 ;
    wire signal_8312 ;
    wire signal_8313 ;
    wire signal_8314 ;
    wire signal_8315 ;
    wire signal_8316 ;
    wire signal_8317 ;
    wire signal_8318 ;
    wire signal_8319 ;
    wire signal_8320 ;
    wire signal_8321 ;
    wire signal_8322 ;
    wire signal_8323 ;
    wire signal_8324 ;
    wire signal_8325 ;
    wire signal_8326 ;
    wire signal_8327 ;
    wire signal_8328 ;
    wire signal_8329 ;
    wire signal_8330 ;
    wire signal_8331 ;
    wire signal_8332 ;
    wire signal_8333 ;
    wire signal_8334 ;
    wire signal_8335 ;
    wire signal_8336 ;
    wire signal_8337 ;
    wire signal_8338 ;
    wire signal_8339 ;
    wire signal_8340 ;
    wire signal_8341 ;
    wire signal_8342 ;
    wire signal_8343 ;
    wire signal_8344 ;
    wire signal_8345 ;
    wire signal_8346 ;
    wire signal_8347 ;
    wire signal_8348 ;
    wire signal_8349 ;
    wire signal_8350 ;
    wire signal_8351 ;
    wire signal_8352 ;
    wire signal_8353 ;
    wire signal_8354 ;
    wire signal_8355 ;
    wire signal_8356 ;
    wire signal_8357 ;
    wire signal_8358 ;
    wire signal_8359 ;
    wire signal_8360 ;
    wire signal_8361 ;
    wire signal_8362 ;
    wire signal_8363 ;
    wire signal_8364 ;
    wire signal_8365 ;
    wire signal_8366 ;
    wire signal_8367 ;
    wire signal_8368 ;
    wire signal_8369 ;
    wire signal_8370 ;
    wire signal_8371 ;
    wire signal_8372 ;
    wire signal_8373 ;
    wire signal_8374 ;
    wire signal_8375 ;
    wire signal_8376 ;
    wire signal_8377 ;
    wire signal_8378 ;
    wire signal_8379 ;
    wire signal_8380 ;
    wire signal_8381 ;
    wire signal_8382 ;
    wire signal_8383 ;
    wire signal_8384 ;
    wire signal_8385 ;
    wire signal_8386 ;
    wire signal_8387 ;
    wire signal_8388 ;
    wire signal_8389 ;
    wire signal_8390 ;
    wire signal_8391 ;
    wire signal_8392 ;
    wire signal_8393 ;
    wire signal_8394 ;
    wire signal_8395 ;
    wire signal_8396 ;
    wire signal_8397 ;
    wire signal_8398 ;
    wire signal_8399 ;
    wire signal_8400 ;
    wire signal_8401 ;
    wire signal_8402 ;
    wire signal_8403 ;
    wire signal_8404 ;
    wire signal_8405 ;
    wire signal_8406 ;
    wire signal_8407 ;
    wire signal_8408 ;
    wire signal_8409 ;
    wire signal_8410 ;
    wire signal_8411 ;
    wire signal_8412 ;
    wire signal_8413 ;
    wire signal_8414 ;
    wire signal_8415 ;
    wire signal_8416 ;
    wire signal_8417 ;
    wire signal_8418 ;
    wire signal_8419 ;
    wire signal_8420 ;
    wire signal_8421 ;
    wire signal_8422 ;
    wire signal_8423 ;
    wire signal_8424 ;
    wire signal_8425 ;
    wire signal_8426 ;
    wire signal_8427 ;
    wire signal_8428 ;
    wire signal_8429 ;
    wire signal_8430 ;
    wire signal_8431 ;
    wire signal_8432 ;
    wire signal_8433 ;
    wire signal_8434 ;
    wire signal_8435 ;
    wire signal_8436 ;
    wire signal_8437 ;
    wire signal_8438 ;
    wire signal_8439 ;
    wire signal_8440 ;
    wire signal_8441 ;
    wire signal_8442 ;
    wire signal_8443 ;
    wire signal_8444 ;
    wire signal_8445 ;
    wire signal_8446 ;
    wire signal_8447 ;
    wire signal_8448 ;
    wire signal_8449 ;
    wire signal_8450 ;
    wire signal_8451 ;
    wire signal_8452 ;
    wire signal_8453 ;
    wire signal_8454 ;
    wire signal_8455 ;
    wire signal_8456 ;
    wire signal_8457 ;
    wire signal_8458 ;
    wire signal_8459 ;
    wire signal_8460 ;
    wire signal_8461 ;
    wire signal_8462 ;
    wire signal_8463 ;
    wire signal_8464 ;
    wire signal_8465 ;
    wire signal_8466 ;
    wire signal_8467 ;
    wire signal_8468 ;
    wire signal_8469 ;
    wire signal_8470 ;
    wire signal_8471 ;
    wire signal_8472 ;
    wire signal_8473 ;
    wire signal_8474 ;
    wire signal_8475 ;
    wire signal_8476 ;
    wire signal_8477 ;
    wire signal_8478 ;
    wire signal_8479 ;
    wire signal_8480 ;
    wire signal_8481 ;
    wire signal_8482 ;
    wire signal_8483 ;
    wire signal_8484 ;
    wire signal_8485 ;
    wire signal_8486 ;
    wire signal_8487 ;
    wire signal_8488 ;
    wire signal_8489 ;
    wire signal_8490 ;
    wire signal_8491 ;
    wire signal_8492 ;
    wire signal_8493 ;
    wire signal_8494 ;
    wire signal_8495 ;
    wire signal_8496 ;
    wire signal_8497 ;
    wire signal_8498 ;
    wire signal_8499 ;
    wire signal_8500 ;
    wire signal_8501 ;
    wire signal_8502 ;
    wire signal_8503 ;
    wire signal_8504 ;
    wire signal_8505 ;
    wire signal_8506 ;
    wire signal_8507 ;
    wire signal_8508 ;
    wire signal_8509 ;
    wire signal_8510 ;
    wire signal_8511 ;
    wire signal_8512 ;
    wire signal_8513 ;
    wire signal_8514 ;
    wire signal_8515 ;
    wire signal_8516 ;
    wire signal_8517 ;
    wire signal_8518 ;
    wire signal_8519 ;
    wire signal_8520 ;
    wire signal_8521 ;
    wire signal_8522 ;
    wire signal_8523 ;
    wire signal_8524 ;
    wire signal_8525 ;
    wire signal_8526 ;
    wire signal_8527 ;
    wire signal_8528 ;
    wire signal_8529 ;
    wire signal_8530 ;
    wire signal_8531 ;
    wire signal_8532 ;
    wire signal_8533 ;
    wire signal_8534 ;
    wire signal_8535 ;
    wire signal_8536 ;
    wire signal_8537 ;
    wire signal_8538 ;
    wire signal_8539 ;
    wire signal_8540 ;
    wire signal_8541 ;
    wire signal_8542 ;
    wire signal_8543 ;
    wire signal_8544 ;
    wire signal_8545 ;
    wire signal_8546 ;
    wire signal_8547 ;
    wire signal_8548 ;
    wire signal_8549 ;
    wire signal_8550 ;
    wire signal_8551 ;
    wire signal_8552 ;
    wire signal_8553 ;
    wire signal_8554 ;
    wire signal_8555 ;
    wire signal_8556 ;
    wire signal_8557 ;
    wire signal_8558 ;
    wire signal_8559 ;
    wire signal_8560 ;
    wire signal_8561 ;
    wire signal_8562 ;
    wire signal_8563 ;
    wire signal_8564 ;
    wire signal_8565 ;
    wire signal_8566 ;
    wire signal_8567 ;
    wire signal_8568 ;
    wire signal_8569 ;
    wire signal_8570 ;
    wire signal_8571 ;
    wire signal_8572 ;
    wire signal_8573 ;
    wire signal_8574 ;
    wire signal_8575 ;
    wire signal_8576 ;
    wire signal_8577 ;
    wire signal_8578 ;
    wire signal_8579 ;
    wire signal_8580 ;
    wire signal_8581 ;
    wire signal_8582 ;
    wire signal_8583 ;
    wire signal_8584 ;
    wire signal_8585 ;
    wire signal_8586 ;
    wire signal_8587 ;
    wire signal_8588 ;
    wire signal_8589 ;
    wire signal_8590 ;
    wire signal_8591 ;
    wire signal_8592 ;
    wire signal_8593 ;
    wire signal_8594 ;
    wire signal_8595 ;
    wire signal_8596 ;
    wire signal_8597 ;
    wire signal_8598 ;
    wire signal_8599 ;
    wire signal_8600 ;
    wire signal_8601 ;
    wire signal_8602 ;
    wire signal_8603 ;
    wire signal_8604 ;
    wire signal_8605 ;
    wire signal_8606 ;
    wire signal_8607 ;
    wire signal_8608 ;
    wire signal_8609 ;
    wire signal_8610 ;
    wire signal_8611 ;
    wire signal_8612 ;
    wire signal_8613 ;
    wire signal_8614 ;
    wire signal_8615 ;
    wire signal_8616 ;
    wire signal_8617 ;
    wire signal_8618 ;
    wire signal_8619 ;
    wire signal_8620 ;
    wire signal_8621 ;
    wire signal_8622 ;
    wire signal_8623 ;
    wire signal_8624 ;
    wire signal_8625 ;
    wire signal_8626 ;
    wire signal_8627 ;
    wire signal_8628 ;
    wire signal_8629 ;
    wire signal_8630 ;
    wire signal_8631 ;
    wire signal_8632 ;
    wire signal_8633 ;
    wire signal_8634 ;
    wire signal_8635 ;
    wire signal_8636 ;
    wire signal_8637 ;
    wire signal_8638 ;
    wire signal_8639 ;
    wire signal_8640 ;
    wire signal_8641 ;
    wire signal_8642 ;
    wire signal_8643 ;
    wire signal_8644 ;
    wire signal_8645 ;
    wire signal_8646 ;
    wire signal_8647 ;
    wire signal_8648 ;
    wire signal_8649 ;
    wire signal_8650 ;
    wire signal_8651 ;
    wire signal_8652 ;
    wire signal_8653 ;
    wire signal_8654 ;
    wire signal_8655 ;
    wire signal_8656 ;
    wire signal_8657 ;
    wire signal_8658 ;
    wire signal_8659 ;
    wire signal_8660 ;
    wire signal_8661 ;
    wire signal_8662 ;
    wire signal_8663 ;
    wire signal_8664 ;
    wire signal_8665 ;
    wire signal_8666 ;
    wire signal_8667 ;
    wire signal_8668 ;
    wire signal_8669 ;
    wire signal_8670 ;
    wire signal_8671 ;
    wire signal_8672 ;
    wire signal_8673 ;
    wire signal_8674 ;
    wire signal_8675 ;
    wire signal_8676 ;
    wire signal_8677 ;
    wire signal_8678 ;
    wire signal_8679 ;
    wire signal_8680 ;
    wire signal_8681 ;
    wire signal_8682 ;
    wire signal_8683 ;
    wire signal_8684 ;
    wire signal_8685 ;
    wire signal_8686 ;
    wire signal_8687 ;
    wire signal_8688 ;
    wire signal_8689 ;
    wire signal_8690 ;
    wire signal_8691 ;
    wire signal_8692 ;
    wire signal_8693 ;
    wire signal_8694 ;
    wire signal_8695 ;
    wire signal_8696 ;
    wire signal_8697 ;
    wire signal_8698 ;
    wire signal_8699 ;
    wire signal_8700 ;
    wire signal_8701 ;
    wire signal_8702 ;
    wire signal_8703 ;
    wire signal_8704 ;
    wire signal_8705 ;
    wire signal_8706 ;
    wire signal_8707 ;
    wire signal_8708 ;
    wire signal_8709 ;
    wire signal_8710 ;
    wire signal_8711 ;
    wire signal_8712 ;
    wire signal_8713 ;
    wire signal_8714 ;
    wire signal_8715 ;
    wire signal_8716 ;
    wire signal_8717 ;
    wire signal_8718 ;
    wire signal_8719 ;
    wire signal_8720 ;
    wire signal_8721 ;
    wire signal_8722 ;
    wire signal_8723 ;
    wire signal_8724 ;
    wire signal_8725 ;
    wire signal_8726 ;
    wire signal_8727 ;
    wire signal_8728 ;
    wire signal_8729 ;
    wire signal_8730 ;
    wire signal_8731 ;
    wire signal_8732 ;
    wire signal_8733 ;
    wire signal_8734 ;
    wire signal_8735 ;
    wire signal_8736 ;
    wire signal_8737 ;
    wire signal_8738 ;
    wire signal_8739 ;
    wire signal_8740 ;
    wire signal_8741 ;
    wire signal_8742 ;
    wire signal_8743 ;
    wire signal_8744 ;
    wire signal_8745 ;
    wire signal_8746 ;
    wire signal_8747 ;
    wire signal_8748 ;
    wire signal_8749 ;
    wire signal_8750 ;
    wire signal_8751 ;
    wire signal_8752 ;
    wire signal_8753 ;
    wire signal_8754 ;
    wire signal_8755 ;
    wire signal_8756 ;
    wire signal_8757 ;
    wire signal_8758 ;
    wire signal_8759 ;
    wire signal_8760 ;
    wire signal_8761 ;
    wire signal_8762 ;
    wire signal_8763 ;
    wire signal_8764 ;
    wire signal_8765 ;
    wire signal_8766 ;
    wire signal_8767 ;
    wire signal_8768 ;
    wire signal_8769 ;
    wire signal_8770 ;
    wire signal_8771 ;
    wire signal_8772 ;
    wire signal_8773 ;
    wire signal_8774 ;
    wire signal_8775 ;
    wire signal_8776 ;
    wire signal_8777 ;
    wire signal_8778 ;
    wire signal_8779 ;
    wire signal_8780 ;
    wire signal_8781 ;
    wire signal_8782 ;
    wire signal_8783 ;
    wire signal_8784 ;
    wire signal_8785 ;
    wire signal_8786 ;
    wire signal_8787 ;
    wire signal_8788 ;
    wire signal_8789 ;
    wire signal_8790 ;
    wire signal_8791 ;
    wire signal_8792 ;
    wire signal_8793 ;
    wire signal_8794 ;
    wire signal_8795 ;
    wire signal_8796 ;
    wire signal_8797 ;
    wire signal_8798 ;
    wire signal_8799 ;
    wire signal_8800 ;
    wire signal_8801 ;
    wire signal_8802 ;
    wire signal_8803 ;
    wire signal_8804 ;
    wire signal_8805 ;
    wire signal_8806 ;
    wire signal_8807 ;
    wire signal_8808 ;
    wire signal_8809 ;
    wire signal_8810 ;
    wire signal_8811 ;
    wire signal_8812 ;
    wire signal_8813 ;
    wire signal_8814 ;
    wire signal_8815 ;
    wire signal_8816 ;
    wire signal_8817 ;
    wire signal_8818 ;
    wire signal_8819 ;
    wire signal_8820 ;
    wire signal_8821 ;
    wire signal_8822 ;
    wire signal_8823 ;
    wire signal_8824 ;
    wire signal_8825 ;
    wire signal_8826 ;
    wire signal_8827 ;
    wire signal_8828 ;
    wire signal_8829 ;
    wire signal_8830 ;
    wire signal_8831 ;
    wire signal_8832 ;
    wire signal_8833 ;
    wire signal_8834 ;
    wire signal_8835 ;
    wire signal_8836 ;
    wire signal_8837 ;
    wire signal_8838 ;
    wire signal_8839 ;
    wire signal_8840 ;
    wire signal_8841 ;
    wire signal_8842 ;
    wire signal_8843 ;
    wire signal_8844 ;
    wire signal_8845 ;
    wire signal_8846 ;
    wire signal_8847 ;
    wire signal_8848 ;
    wire signal_8849 ;
    wire signal_8850 ;
    wire signal_8851 ;
    wire signal_8852 ;
    wire signal_8853 ;
    wire signal_8854 ;
    wire signal_8855 ;
    wire signal_8856 ;
    wire signal_8857 ;
    wire signal_8858 ;
    wire signal_8859 ;
    wire signal_8860 ;
    wire signal_8861 ;
    wire signal_8862 ;
    wire signal_8863 ;
    wire signal_8864 ;
    wire signal_8865 ;
    wire signal_8866 ;
    wire signal_8867 ;
    wire signal_8868 ;
    wire signal_8869 ;
    wire signal_8870 ;
    wire signal_8871 ;
    wire signal_8872 ;
    wire signal_8873 ;
    wire signal_8874 ;
    wire signal_8875 ;
    wire signal_8876 ;
    wire signal_8877 ;
    wire signal_8878 ;
    wire signal_8879 ;
    wire signal_8880 ;
    wire signal_8881 ;
    wire signal_8882 ;
    wire signal_8883 ;
    wire signal_8884 ;
    wire signal_8885 ;
    wire signal_8886 ;
    wire signal_8887 ;
    wire signal_8888 ;
    wire signal_8889 ;
    wire signal_8890 ;
    wire signal_8891 ;
    wire signal_8892 ;
    wire signal_8893 ;
    wire signal_8894 ;
    wire signal_8895 ;
    wire signal_8896 ;
    wire signal_8897 ;
    wire signal_8898 ;
    wire signal_8899 ;
    wire signal_8900 ;
    wire signal_8901 ;
    wire signal_8902 ;
    wire signal_8903 ;
    wire signal_8904 ;
    wire signal_8905 ;
    wire signal_8906 ;
    wire signal_8907 ;
    wire signal_8908 ;
    wire signal_8909 ;
    wire signal_8910 ;
    wire signal_8911 ;
    wire signal_8912 ;
    wire signal_8913 ;
    wire signal_8914 ;
    wire signal_8915 ;
    wire signal_8916 ;
    wire signal_8917 ;
    wire signal_8918 ;
    wire signal_8919 ;
    wire signal_8920 ;
    wire signal_8921 ;
    wire signal_8922 ;
    wire signal_8923 ;
    wire signal_8924 ;
    wire signal_8925 ;
    wire signal_8926 ;
    wire signal_8927 ;
    wire signal_8928 ;
    wire signal_8929 ;
    wire signal_8930 ;
    wire signal_8931 ;
    wire signal_8932 ;
    wire signal_8933 ;
    wire signal_8934 ;
    wire signal_8935 ;
    wire signal_8936 ;
    wire signal_8937 ;
    wire signal_8938 ;
    wire signal_8939 ;
    wire signal_8940 ;
    wire signal_8941 ;
    wire signal_8942 ;
    wire signal_8943 ;
    wire signal_8944 ;
    wire signal_8945 ;
    wire signal_8946 ;
    wire signal_8947 ;
    wire signal_8948 ;
    wire signal_8949 ;
    wire signal_8950 ;
    wire signal_8951 ;
    wire signal_8952 ;
    wire signal_8953 ;
    wire signal_8954 ;
    wire signal_8955 ;
    wire signal_8956 ;
    wire signal_8957 ;
    wire signal_8958 ;
    wire signal_8959 ;
    wire signal_8960 ;
    wire signal_8961 ;
    wire signal_8962 ;
    wire signal_8963 ;
    wire signal_8964 ;
    wire signal_8965 ;
    wire signal_8966 ;
    wire signal_8967 ;
    wire signal_8968 ;
    wire signal_8969 ;
    wire signal_8970 ;
    wire signal_8971 ;
    wire signal_8972 ;
    wire signal_8973 ;
    wire signal_8974 ;
    wire signal_8975 ;
    wire signal_8976 ;
    wire signal_8977 ;
    wire signal_8978 ;
    wire signal_8979 ;
    wire signal_8980 ;
    wire signal_8981 ;
    wire signal_8982 ;
    wire signal_8983 ;
    wire signal_8984 ;
    wire signal_8985 ;
    wire signal_8986 ;
    wire signal_8987 ;
    wire signal_8988 ;
    wire signal_8989 ;
    wire signal_8990 ;
    wire signal_8991 ;
    wire signal_8992 ;
    wire signal_8993 ;
    wire signal_8994 ;
    wire signal_8995 ;
    wire signal_8996 ;
    wire signal_8997 ;
    wire signal_8998 ;
    wire signal_8999 ;
    wire signal_9000 ;
    wire signal_9001 ;
    wire signal_9002 ;
    wire signal_9003 ;
    wire signal_9004 ;
    wire signal_9005 ;
    wire signal_9006 ;
    wire signal_9007 ;
    wire signal_9008 ;
    wire signal_9009 ;
    wire signal_9010 ;
    wire signal_9011 ;
    wire signal_9012 ;
    wire signal_9013 ;
    wire signal_9014 ;
    wire signal_9015 ;
    wire signal_9016 ;
    wire signal_9017 ;
    wire signal_9018 ;
    wire signal_9019 ;
    wire signal_9020 ;
    wire signal_9021 ;
    wire signal_9022 ;
    wire signal_9023 ;
    wire signal_9024 ;
    wire signal_9025 ;
    wire signal_9026 ;
    wire signal_9027 ;
    wire signal_9028 ;
    wire signal_9029 ;
    wire signal_9030 ;
    wire signal_9031 ;
    wire signal_9032 ;
    wire signal_9033 ;
    wire signal_9034 ;
    wire signal_9035 ;
    wire signal_9036 ;
    wire signal_9037 ;
    wire signal_9038 ;
    wire signal_9039 ;
    wire signal_9040 ;
    wire signal_9041 ;
    wire signal_9042 ;
    wire signal_9043 ;
    wire signal_9044 ;
    wire signal_9045 ;
    wire signal_9046 ;
    wire signal_9047 ;
    wire signal_9048 ;
    wire signal_9049 ;
    wire signal_9050 ;
    wire signal_9051 ;
    wire signal_9052 ;
    wire signal_9053 ;
    wire signal_9054 ;
    wire signal_9055 ;
    wire signal_9056 ;
    wire signal_9057 ;
    wire signal_9058 ;
    wire signal_9059 ;
    wire signal_9060 ;
    wire signal_9061 ;
    wire signal_9062 ;
    wire signal_9063 ;
    wire signal_9064 ;
    wire signal_9065 ;
    wire signal_9066 ;
    wire signal_9067 ;
    wire signal_9068 ;
    wire signal_9069 ;
    wire signal_9070 ;
    wire signal_9071 ;
    wire signal_9072 ;
    wire signal_9073 ;
    wire signal_9074 ;
    wire signal_9075 ;
    wire signal_9076 ;
    wire signal_9077 ;
    wire signal_9078 ;
    wire signal_9079 ;
    wire signal_9080 ;
    wire signal_9081 ;
    wire signal_9082 ;
    wire signal_9083 ;
    wire signal_9084 ;
    wire signal_9085 ;
    wire signal_9086 ;
    wire signal_9087 ;
    wire signal_9088 ;
    wire signal_9089 ;
    wire signal_9090 ;
    wire signal_9091 ;
    wire signal_9092 ;
    wire signal_9093 ;
    wire signal_9094 ;
    wire signal_9095 ;
    wire signal_9096 ;
    wire signal_9097 ;
    wire signal_9098 ;
    wire signal_9099 ;
    wire signal_9100 ;
    wire signal_9101 ;
    wire signal_9102 ;
    wire signal_9103 ;
    wire signal_9104 ;
    wire signal_9105 ;
    wire signal_9106 ;
    wire signal_9107 ;
    wire signal_9108 ;
    wire signal_9109 ;
    wire signal_9110 ;
    wire signal_9111 ;
    wire signal_9112 ;
    wire signal_9113 ;
    wire signal_9114 ;
    wire signal_9115 ;
    wire signal_9116 ;
    wire signal_9117 ;
    wire signal_9118 ;
    wire signal_9119 ;
    wire signal_9120 ;
    wire signal_9121 ;
    wire signal_9122 ;
    wire signal_9123 ;
    wire signal_9124 ;
    wire signal_9125 ;
    wire signal_9126 ;
    wire signal_9127 ;
    wire signal_9128 ;
    wire signal_9129 ;
    wire signal_9130 ;
    wire signal_9131 ;
    wire signal_9132 ;
    wire signal_9133 ;
    wire signal_9134 ;
    wire signal_9135 ;
    wire signal_9136 ;
    wire signal_9137 ;
    wire signal_9138 ;
    wire signal_9139 ;
    wire signal_9140 ;
    wire signal_9141 ;
    wire signal_9142 ;
    wire signal_9143 ;
    wire signal_9144 ;
    wire signal_9145 ;
    wire signal_9146 ;
    wire signal_9147 ;
    wire signal_9148 ;
    wire signal_9149 ;
    wire signal_9150 ;
    wire signal_9151 ;
    wire signal_9152 ;
    wire signal_9153 ;
    wire signal_9154 ;
    wire signal_9155 ;
    wire signal_9156 ;
    wire signal_9157 ;
    wire signal_9158 ;
    wire signal_9159 ;
    wire signal_9160 ;
    wire signal_9161 ;
    wire signal_9162 ;
    wire signal_9163 ;
    wire signal_9164 ;
    wire signal_9165 ;
    wire signal_9166 ;
    wire signal_9167 ;
    wire signal_9168 ;
    wire signal_9169 ;
    wire signal_9170 ;
    wire signal_9171 ;
    wire signal_9172 ;
    wire signal_9173 ;
    wire signal_9174 ;
    wire signal_9175 ;
    wire signal_9176 ;
    wire signal_9177 ;
    wire signal_9178 ;
    wire signal_9179 ;
    wire signal_9180 ;
    wire signal_9181 ;
    wire signal_9182 ;
    wire signal_9183 ;
    wire signal_9184 ;
    wire signal_9185 ;
    wire signal_9186 ;
    wire signal_9187 ;
    wire signal_9188 ;
    wire signal_9189 ;
    wire signal_9190 ;
    wire signal_9191 ;
    wire signal_9192 ;
    wire signal_9193 ;
    wire signal_9194 ;
    wire signal_9195 ;
    wire signal_9196 ;
    wire signal_9197 ;
    wire signal_9198 ;
    wire signal_9199 ;
    wire signal_9200 ;
    wire signal_9201 ;
    wire signal_9202 ;
    wire signal_9203 ;
    wire signal_9204 ;
    wire signal_9205 ;
    wire signal_9206 ;
    wire signal_9207 ;
    wire signal_9208 ;
    wire signal_9209 ;
    wire signal_9210 ;
    wire signal_9211 ;
    wire signal_9212 ;
    wire signal_9213 ;
    wire signal_9214 ;
    wire signal_9215 ;
    wire signal_9216 ;
    wire signal_9217 ;
    wire signal_9218 ;
    wire signal_9219 ;
    wire signal_9220 ;
    wire signal_9221 ;
    wire signal_9222 ;
    wire signal_9223 ;
    wire signal_9224 ;
    wire signal_9225 ;
    wire signal_9226 ;
    wire signal_9227 ;
    wire signal_9228 ;
    wire signal_9229 ;
    wire signal_9230 ;
    wire signal_9231 ;
    wire signal_9232 ;
    wire signal_9233 ;
    wire signal_9234 ;
    wire signal_9235 ;
    wire signal_9236 ;
    wire signal_9237 ;
    wire signal_9238 ;
    wire signal_9239 ;
    wire signal_9240 ;
    wire signal_9241 ;
    wire signal_9242 ;
    wire signal_9243 ;
    wire signal_9244 ;
    wire signal_9245 ;
    wire signal_9246 ;
    wire signal_9247 ;
    wire signal_9248 ;
    wire signal_9249 ;
    wire signal_9250 ;
    wire signal_9251 ;
    wire signal_9252 ;
    wire signal_9253 ;
    wire signal_9254 ;
    wire signal_9255 ;
    wire signal_9256 ;
    wire signal_9257 ;
    wire signal_9258 ;
    wire signal_9259 ;
    wire signal_9260 ;
    wire signal_9261 ;
    wire signal_9262 ;
    wire signal_9263 ;
    wire signal_9264 ;
    wire signal_9265 ;
    wire signal_9266 ;
    wire signal_9267 ;
    wire signal_9268 ;
    wire signal_9269 ;
    wire signal_9270 ;
    wire signal_9271 ;
    wire signal_9272 ;
    wire signal_9273 ;
    wire signal_9274 ;
    wire signal_9275 ;
    wire signal_9276 ;
    wire signal_9277 ;
    wire signal_9278 ;
    wire signal_9279 ;
    wire signal_9280 ;
    wire signal_9281 ;
    wire signal_9282 ;
    wire signal_9283 ;
    wire signal_9284 ;
    wire signal_9285 ;
    wire signal_9286 ;
    wire signal_9287 ;
    wire signal_9288 ;
    wire signal_9289 ;
    wire signal_9290 ;
    wire signal_9291 ;
    wire signal_9292 ;
    wire signal_9293 ;
    wire signal_9294 ;
    wire signal_9295 ;
    wire signal_9296 ;
    wire signal_9297 ;
    wire signal_9298 ;
    wire signal_9299 ;
    wire signal_9300 ;
    wire signal_9301 ;
    wire signal_9302 ;
    wire signal_9303 ;
    wire signal_9304 ;
    wire signal_9305 ;
    wire signal_9306 ;
    wire signal_9307 ;
    wire signal_9308 ;
    wire signal_9309 ;
    wire signal_9310 ;
    wire signal_9311 ;
    wire signal_9312 ;
    wire signal_9313 ;
    wire signal_9314 ;
    wire signal_9315 ;
    wire signal_9316 ;
    wire signal_9317 ;
    wire signal_9318 ;
    wire signal_9319 ;
    wire signal_9320 ;
    wire signal_9321 ;
    wire signal_9322 ;
    wire signal_9323 ;
    wire signal_9324 ;
    wire signal_9325 ;
    wire signal_9326 ;
    wire signal_9327 ;
    wire signal_9328 ;
    wire signal_9329 ;
    wire signal_9330 ;
    wire signal_9331 ;
    wire signal_9332 ;
    wire signal_9333 ;
    wire signal_9334 ;
    wire signal_9335 ;
    wire signal_9336 ;
    wire signal_9337 ;
    wire signal_9338 ;
    wire signal_9339 ;
    wire signal_9340 ;
    wire signal_9341 ;
    wire signal_9342 ;
    wire signal_9343 ;
    wire signal_9344 ;
    wire signal_9345 ;
    wire signal_9346 ;
    wire signal_9347 ;
    wire signal_9348 ;
    wire signal_9349 ;
    wire signal_9350 ;
    wire signal_9351 ;
    wire signal_9352 ;
    wire signal_9353 ;
    wire signal_9354 ;
    wire signal_9355 ;
    wire signal_9356 ;
    wire signal_9357 ;
    wire signal_9358 ;
    wire signal_9359 ;
    wire signal_9360 ;
    wire signal_9361 ;
    wire signal_9362 ;
    wire signal_9363 ;
    wire signal_9364 ;
    wire signal_9365 ;
    wire signal_9366 ;
    wire signal_9367 ;
    wire signal_9368 ;
    wire signal_9369 ;
    wire signal_9370 ;
    wire signal_9371 ;
    wire signal_9372 ;
    wire signal_9373 ;
    wire signal_9374 ;
    wire signal_9375 ;
    wire signal_9376 ;
    wire signal_9377 ;
    wire signal_9378 ;
    wire signal_9379 ;
    wire signal_9380 ;
    wire signal_9381 ;
    wire signal_9382 ;
    wire signal_9383 ;
    wire signal_9384 ;
    wire signal_9385 ;
    wire signal_9386 ;
    wire signal_9387 ;
    wire signal_9388 ;
    wire signal_9389 ;
    wire signal_9390 ;
    wire signal_9391 ;
    wire signal_9392 ;
    wire signal_9393 ;
    wire signal_9394 ;
    wire signal_9395 ;
    wire signal_9396 ;
    wire signal_9397 ;
    wire signal_9398 ;
    wire signal_9399 ;
    wire signal_9400 ;
    wire signal_9401 ;
    wire signal_9402 ;
    wire signal_9403 ;
    wire signal_9404 ;
    wire signal_9405 ;
    wire signal_9406 ;
    wire signal_9407 ;
    wire signal_9408 ;
    wire signal_9409 ;
    wire signal_9410 ;
    wire signal_9411 ;
    wire signal_9412 ;
    wire signal_9413 ;
    wire signal_9414 ;
    wire signal_9415 ;
    wire signal_9416 ;
    wire signal_9417 ;
    wire signal_9418 ;
    wire signal_9419 ;
    wire signal_9420 ;
    wire signal_9421 ;
    wire signal_9422 ;
    wire signal_9423 ;
    wire signal_9424 ;
    wire signal_9425 ;
    wire signal_9426 ;
    wire signal_9427 ;
    wire signal_9428 ;
    wire signal_9429 ;
    wire signal_9430 ;
    wire signal_9431 ;
    wire signal_9432 ;
    wire signal_9433 ;
    wire signal_9434 ;
    wire signal_9435 ;
    wire signal_9436 ;
    wire signal_9437 ;
    wire signal_9438 ;
    wire signal_9439 ;
    wire signal_9440 ;
    wire signal_9441 ;
    wire signal_9442 ;
    wire signal_9443 ;
    wire signal_9444 ;
    wire signal_9445 ;
    wire signal_9446 ;
    wire signal_9447 ;
    wire signal_9448 ;
    wire signal_9449 ;
    wire signal_9450 ;
    wire signal_9451 ;
    wire signal_9452 ;
    wire signal_9453 ;
    wire signal_9454 ;
    wire signal_9455 ;
    wire signal_9456 ;
    wire signal_9457 ;
    wire signal_9458 ;
    wire signal_9459 ;
    wire signal_9460 ;
    wire signal_9461 ;
    wire signal_9462 ;
    wire signal_9463 ;
    wire signal_9464 ;
    wire signal_9465 ;
    wire signal_9466 ;
    wire signal_9467 ;
    wire signal_9468 ;
    wire signal_9469 ;
    wire signal_9470 ;
    wire signal_9471 ;
    wire signal_9472 ;
    wire signal_9473 ;
    wire signal_9474 ;
    wire signal_9475 ;
    wire signal_9476 ;
    wire signal_9477 ;
    wire signal_9478 ;
    wire signal_9479 ;
    wire signal_9480 ;
    wire signal_9481 ;
    wire signal_9482 ;
    wire signal_9483 ;
    wire signal_9484 ;
    wire signal_9485 ;
    wire signal_9486 ;
    wire signal_9487 ;
    wire signal_9488 ;
    wire signal_9489 ;
    wire signal_9490 ;
    wire signal_9491 ;
    wire signal_9492 ;
    wire signal_9493 ;
    wire signal_9494 ;
    wire signal_9495 ;
    wire signal_9496 ;
    wire signal_9497 ;
    wire signal_9498 ;
    wire signal_9499 ;
    wire signal_9500 ;
    wire signal_9501 ;
    wire signal_9502 ;
    wire signal_9503 ;
    wire signal_9504 ;
    wire signal_9505 ;
    wire signal_9506 ;
    wire signal_9507 ;
    wire signal_9508 ;
    wire signal_9509 ;
    wire signal_9510 ;
    wire signal_9511 ;
    wire signal_9512 ;
    wire signal_9513 ;
    wire signal_9514 ;
    wire signal_9515 ;
    wire signal_9516 ;
    wire signal_9517 ;
    wire signal_9518 ;
    wire signal_9519 ;
    wire signal_9520 ;
    wire signal_9521 ;
    wire signal_9522 ;
    wire signal_9523 ;
    wire signal_9524 ;
    wire signal_9525 ;
    wire signal_9526 ;
    wire signal_9527 ;
    wire signal_9528 ;
    wire signal_9529 ;
    wire signal_9530 ;
    wire signal_9531 ;
    wire signal_9532 ;
    wire signal_9533 ;
    wire signal_9534 ;
    wire signal_9535 ;
    wire signal_9536 ;
    wire signal_9537 ;
    wire signal_9538 ;
    wire signal_9539 ;
    wire signal_9540 ;
    wire signal_9541 ;
    wire signal_9542 ;
    wire signal_9543 ;
    wire signal_9544 ;
    wire signal_9545 ;
    wire signal_9546 ;
    wire signal_9547 ;
    wire signal_9548 ;
    wire signal_9549 ;
    wire signal_9550 ;
    wire signal_9551 ;
    wire signal_9552 ;
    wire signal_9553 ;
    wire signal_9554 ;
    wire signal_9555 ;
    wire signal_9556 ;
    wire signal_9557 ;
    wire signal_9558 ;
    wire signal_9559 ;
    wire signal_9560 ;
    wire signal_9561 ;
    wire signal_9562 ;
    wire signal_9563 ;
    wire signal_9564 ;
    wire signal_9565 ;
    wire signal_9566 ;
    wire signal_9567 ;
    wire signal_9568 ;
    wire signal_9569 ;
    wire signal_9570 ;
    wire signal_9571 ;
    wire signal_9572 ;
    wire signal_9573 ;
    wire signal_9574 ;
    wire signal_9575 ;
    wire signal_9576 ;
    wire signal_9577 ;
    wire signal_9578 ;
    wire signal_9579 ;
    wire signal_9580 ;
    wire signal_9581 ;
    wire signal_9582 ;
    wire signal_9583 ;
    wire signal_9584 ;
    wire signal_9585 ;
    wire signal_9586 ;
    wire signal_9587 ;
    wire signal_9588 ;
    wire signal_9589 ;
    wire signal_9590 ;
    wire signal_9591 ;
    wire signal_9592 ;
    wire signal_9593 ;
    wire signal_9594 ;
    wire signal_9595 ;
    wire signal_9596 ;
    wire signal_9597 ;
    wire signal_9598 ;
    wire signal_9599 ;
    wire signal_9600 ;
    wire signal_9601 ;
    wire signal_9602 ;
    wire signal_9603 ;
    wire signal_9604 ;
    wire signal_9605 ;
    wire signal_9606 ;
    wire signal_9607 ;
    wire signal_9608 ;
    wire signal_9609 ;
    wire signal_9610 ;
    wire signal_9611 ;
    wire signal_9612 ;
    wire signal_9613 ;
    wire signal_9614 ;
    wire signal_9615 ;
    wire signal_9616 ;
    wire signal_9617 ;
    wire signal_9618 ;
    wire signal_9619 ;
    wire signal_9620 ;
    wire signal_9621 ;
    wire signal_9622 ;
    wire signal_9623 ;
    wire signal_9624 ;
    wire signal_9625 ;
    wire signal_9626 ;
    wire signal_9627 ;
    wire signal_9628 ;
    wire signal_9629 ;
    wire signal_9630 ;
    wire signal_9631 ;
    wire signal_9632 ;
    wire signal_9633 ;
    wire signal_9634 ;
    wire signal_9635 ;
    wire signal_9636 ;
    wire signal_9637 ;
    wire signal_9638 ;
    wire signal_9639 ;
    wire signal_9640 ;
    wire signal_9641 ;
    wire signal_9642 ;
    wire signal_9643 ;
    wire signal_9644 ;
    wire signal_9645 ;
    wire signal_9646 ;
    wire signal_9647 ;
    wire signal_9648 ;
    wire signal_9649 ;
    wire signal_9650 ;
    wire signal_9651 ;
    wire signal_9652 ;
    wire signal_9653 ;
    wire signal_9654 ;
    wire signal_9655 ;
    wire signal_9656 ;
    wire signal_9657 ;
    wire signal_9658 ;
    wire signal_9659 ;
    wire signal_9660 ;
    wire signal_9661 ;
    wire signal_9662 ;
    wire signal_9663 ;
    wire signal_9664 ;
    wire signal_9665 ;
    wire signal_9666 ;
    wire signal_9667 ;
    wire signal_9668 ;
    wire signal_9669 ;
    wire signal_9670 ;
    wire signal_9671 ;
    wire signal_9672 ;
    wire signal_9673 ;
    wire signal_9674 ;
    wire signal_9675 ;
    wire signal_9676 ;
    wire signal_9677 ;
    wire signal_9678 ;
    wire signal_9679 ;
    wire signal_9680 ;
    wire signal_9681 ;
    wire signal_9682 ;
    wire signal_9683 ;
    wire signal_9684 ;
    wire signal_9685 ;
    wire signal_9686 ;
    wire signal_9687 ;
    wire signal_9688 ;
    wire signal_9689 ;
    wire signal_9690 ;
    wire signal_9691 ;
    wire signal_9692 ;
    wire signal_9693 ;
    wire signal_9694 ;
    wire signal_9695 ;
    wire signal_9696 ;
    wire signal_9697 ;
    wire signal_9698 ;
    wire signal_9699 ;
    wire signal_9700 ;
    wire signal_9701 ;
    wire signal_9702 ;
    wire signal_9703 ;
    wire signal_9704 ;
    wire signal_9705 ;
    wire signal_9706 ;
    wire signal_9707 ;
    wire signal_9708 ;
    wire signal_9709 ;
    wire signal_9710 ;
    wire signal_9711 ;
    wire signal_9712 ;
    wire signal_9713 ;
    wire signal_9714 ;
    wire signal_9715 ;
    wire signal_9716 ;
    wire signal_9717 ;
    wire signal_9718 ;
    wire signal_9719 ;
    wire signal_9720 ;
    wire signal_9721 ;
    wire signal_9722 ;
    wire signal_9723 ;
    wire signal_9724 ;
    wire signal_9725 ;
    wire signal_9726 ;
    wire signal_9727 ;
    wire signal_9728 ;
    wire signal_9729 ;
    wire signal_9730 ;
    wire signal_9731 ;
    wire signal_9732 ;
    wire signal_9733 ;
    wire signal_9734 ;
    wire signal_9735 ;
    wire signal_9736 ;
    wire signal_9737 ;
    wire signal_9738 ;
    wire signal_9739 ;
    wire signal_9740 ;
    wire signal_9741 ;
    wire signal_9742 ;
    wire signal_9743 ;
    wire signal_9744 ;
    wire signal_9745 ;
    wire signal_9746 ;
    wire signal_9747 ;
    wire signal_9748 ;
    wire signal_9749 ;
    wire signal_9750 ;
    wire signal_9751 ;
    wire signal_9752 ;
    wire signal_9753 ;
    wire signal_9754 ;
    wire signal_9755 ;
    wire signal_9756 ;
    wire signal_9757 ;
    wire signal_9758 ;
    wire signal_9759 ;
    wire signal_9760 ;
    wire signal_9761 ;
    wire signal_9762 ;
    wire signal_9763 ;
    wire signal_9764 ;
    wire signal_9765 ;
    wire signal_9766 ;
    wire signal_9767 ;
    wire signal_9768 ;
    wire signal_9769 ;
    wire signal_9770 ;
    wire signal_9771 ;
    wire signal_9772 ;
    wire signal_9773 ;
    wire signal_9774 ;
    wire signal_9775 ;
    wire signal_9776 ;
    wire signal_9777 ;
    wire signal_9778 ;
    wire signal_9779 ;
    wire signal_9780 ;
    wire signal_9781 ;
    wire signal_9782 ;
    wire signal_9783 ;
    wire signal_9784 ;
    wire signal_9785 ;
    wire signal_9786 ;
    wire signal_9787 ;
    wire signal_9788 ;
    wire signal_9789 ;
    wire signal_9790 ;
    wire signal_9791 ;
    wire signal_9792 ;
    wire signal_9793 ;
    wire signal_9794 ;
    wire signal_9795 ;
    wire signal_9796 ;
    wire signal_9797 ;
    wire signal_9798 ;
    wire signal_9799 ;
    wire signal_9800 ;
    wire signal_9801 ;
    wire signal_9802 ;
    wire signal_9803 ;
    wire signal_9804 ;
    wire signal_9805 ;
    wire signal_9806 ;
    wire signal_9807 ;
    wire signal_9808 ;
    wire signal_9809 ;
    wire signal_9810 ;
    wire signal_9811 ;
    wire signal_9812 ;
    wire signal_9813 ;
    wire signal_9814 ;
    wire signal_9815 ;
    wire signal_9816 ;
    wire signal_9817 ;
    wire signal_9818 ;
    wire signal_9819 ;
    wire signal_9820 ;
    wire signal_9821 ;
    wire signal_9822 ;
    wire signal_9823 ;
    wire signal_9824 ;
    wire signal_9825 ;
    wire signal_9826 ;
    wire signal_9827 ;
    wire signal_9828 ;
    wire signal_9829 ;
    wire signal_9830 ;
    wire signal_9831 ;
    wire signal_9832 ;
    wire signal_9833 ;
    wire signal_9834 ;
    wire signal_9835 ;
    wire signal_9836 ;
    wire signal_9837 ;
    wire signal_9838 ;
    wire signal_9839 ;
    wire signal_9840 ;
    wire signal_9841 ;
    wire signal_9842 ;
    wire signal_9843 ;
    wire signal_9844 ;
    wire signal_9845 ;
    wire signal_9846 ;
    wire signal_9847 ;
    wire signal_9848 ;
    wire signal_9849 ;
    wire signal_9850 ;
    wire signal_9851 ;
    wire signal_9852 ;
    wire signal_9853 ;
    wire signal_9854 ;
    wire signal_9855 ;
    wire signal_9856 ;
    wire signal_9857 ;
    wire signal_9858 ;
    wire signal_9859 ;
    wire signal_9860 ;
    wire signal_9861 ;
    wire signal_9862 ;
    wire signal_9863 ;
    wire signal_9864 ;
    wire signal_9865 ;
    wire signal_9866 ;
    wire signal_9867 ;
    wire signal_9868 ;
    wire signal_9869 ;
    wire signal_9870 ;
    wire signal_9871 ;
    wire signal_9872 ;
    wire signal_9873 ;
    wire signal_9874 ;
    wire signal_9875 ;
    wire signal_9876 ;
    wire signal_9877 ;
    wire signal_9878 ;
    wire signal_9879 ;
    wire signal_9880 ;
    wire signal_9881 ;
    wire signal_9882 ;
    wire signal_9883 ;
    wire signal_9884 ;
    wire signal_9885 ;
    wire signal_9886 ;
    wire signal_9887 ;
    wire signal_9888 ;
    wire signal_9889 ;
    wire signal_9890 ;
    wire signal_9891 ;
    wire signal_9892 ;
    wire signal_9893 ;
    wire signal_9894 ;
    wire signal_9895 ;
    wire signal_9896 ;
    wire signal_9897 ;
    wire signal_9898 ;
    wire signal_9899 ;
    wire signal_9900 ;
    wire signal_9901 ;
    wire signal_9902 ;
    wire signal_9903 ;
    wire signal_9904 ;
    wire signal_9905 ;
    wire signal_9906 ;
    wire signal_9907 ;
    wire signal_9908 ;
    wire signal_9909 ;
    wire signal_9910 ;
    wire signal_9911 ;
    wire signal_9912 ;
    wire signal_9913 ;
    wire signal_9914 ;
    wire signal_9915 ;
    wire signal_9916 ;
    wire signal_9917 ;
    wire signal_9918 ;
    wire signal_9919 ;
    wire signal_9920 ;
    wire signal_9921 ;
    wire signal_9922 ;
    wire signal_9923 ;
    wire signal_9924 ;
    wire signal_9925 ;
    wire signal_9926 ;
    wire signal_9927 ;
    wire signal_9928 ;
    wire signal_9929 ;
    wire signal_9930 ;
    wire signal_9931 ;
    wire signal_9932 ;
    wire signal_9933 ;
    wire signal_9934 ;
    wire signal_9935 ;
    wire signal_9936 ;
    wire signal_9937 ;
    wire signal_9938 ;
    wire signal_9939 ;
    wire signal_9940 ;
    wire signal_9941 ;
    wire signal_9942 ;
    wire signal_9943 ;
    wire signal_9944 ;
    wire signal_9945 ;
    wire signal_9946 ;
    wire signal_9947 ;
    wire signal_9948 ;
    wire signal_9949 ;
    wire signal_9950 ;
    wire signal_9951 ;
    wire signal_9952 ;
    wire signal_9953 ;
    wire signal_9954 ;
    wire signal_9955 ;
    wire signal_9956 ;
    wire signal_9957 ;
    wire signal_9958 ;
    wire signal_9959 ;
    wire signal_9960 ;
    wire signal_9961 ;
    wire signal_9962 ;
    wire signal_9963 ;
    wire signal_9964 ;
    wire signal_9965 ;
    wire signal_9966 ;
    wire signal_9967 ;
    wire signal_9968 ;
    wire signal_9969 ;
    wire signal_9970 ;
    wire signal_9971 ;
    wire signal_9972 ;
    wire signal_9973 ;
    wire signal_9974 ;
    wire signal_9975 ;
    wire signal_9976 ;
    wire signal_9977 ;
    wire signal_9978 ;
    wire signal_9979 ;
    wire signal_9980 ;
    wire signal_9981 ;
    wire signal_9982 ;
    wire signal_9983 ;
    wire signal_9984 ;
    wire signal_9985 ;
    wire signal_9986 ;
    wire signal_9987 ;
    wire signal_9988 ;
    wire signal_9989 ;
    wire signal_9990 ;
    wire signal_9991 ;
    wire signal_9992 ;
    wire signal_9993 ;
    wire signal_9994 ;
    wire signal_9995 ;
    wire signal_9996 ;
    wire signal_9997 ;
    wire signal_9998 ;
    wire signal_9999 ;
    wire signal_10000 ;
    wire signal_10001 ;
    wire signal_10002 ;
    wire signal_10003 ;
    wire signal_10004 ;
    wire signal_10005 ;
    wire signal_10006 ;
    wire signal_10007 ;
    wire signal_10008 ;
    wire signal_10009 ;
    wire signal_10010 ;
    wire signal_10011 ;
    wire signal_10012 ;
    wire signal_10013 ;
    wire signal_10014 ;
    wire signal_10015 ;
    wire signal_10016 ;
    wire signal_10017 ;
    wire signal_10018 ;
    wire signal_10019 ;
    wire signal_10020 ;
    wire signal_10021 ;
    wire signal_10022 ;
    wire signal_10023 ;
    wire signal_10024 ;
    wire signal_10025 ;
    wire signal_10026 ;
    wire signal_10027 ;
    wire signal_10028 ;
    wire signal_10029 ;
    wire signal_10030 ;
    wire signal_10031 ;
    wire signal_10032 ;
    wire signal_10033 ;
    wire signal_10034 ;
    wire signal_10035 ;
    wire signal_10036 ;
    wire signal_10037 ;
    wire signal_10038 ;
    wire signal_10039 ;
    wire signal_10040 ;
    wire signal_10041 ;
    wire signal_10042 ;
    wire signal_10043 ;
    wire signal_10044 ;
    wire signal_10045 ;
    wire signal_10046 ;
    wire signal_10047 ;
    wire signal_10048 ;
    wire signal_10049 ;
    wire signal_10050 ;
    wire signal_10051 ;
    wire signal_10052 ;
    wire signal_10053 ;
    wire signal_10054 ;
    wire signal_10055 ;
    wire signal_10056 ;
    wire signal_10057 ;
    wire signal_10058 ;
    wire signal_10059 ;
    wire signal_10060 ;
    wire signal_10061 ;
    wire signal_10062 ;
    wire signal_10063 ;
    wire signal_10064 ;
    wire signal_10065 ;
    wire signal_10066 ;
    wire signal_10067 ;
    wire signal_10068 ;
    wire signal_10069 ;
    wire signal_10070 ;
    wire signal_10071 ;
    wire signal_10072 ;
    wire signal_10073 ;
    wire signal_10074 ;
    wire signal_10075 ;
    wire signal_10076 ;
    wire signal_10077 ;
    wire signal_10078 ;
    wire signal_10079 ;
    wire signal_10080 ;
    wire signal_10081 ;
    wire signal_10082 ;
    wire signal_10083 ;
    wire signal_10084 ;
    wire signal_10085 ;
    wire signal_10086 ;
    wire signal_10087 ;
    wire signal_10088 ;
    wire signal_10089 ;
    wire signal_10090 ;
    wire signal_10091 ;
    wire signal_10092 ;
    wire signal_10093 ;
    wire signal_10094 ;
    wire signal_10095 ;
    wire signal_10096 ;
    wire signal_10097 ;
    wire signal_10098 ;
    wire signal_10099 ;
    wire signal_10100 ;
    wire signal_10101 ;
    wire signal_10102 ;
    wire signal_10103 ;
    wire signal_10104 ;
    wire signal_10105 ;
    wire signal_10106 ;
    wire signal_10107 ;
    wire signal_10108 ;
    wire signal_10109 ;
    wire signal_10110 ;
    wire signal_10111 ;
    wire signal_10112 ;
    wire signal_10113 ;
    wire signal_10114 ;
    wire signal_10115 ;
    wire signal_10116 ;
    wire signal_10117 ;
    wire signal_10118 ;
    wire signal_10119 ;
    wire signal_10120 ;
    wire signal_10121 ;
    wire signal_10122 ;
    wire signal_10123 ;
    wire signal_10124 ;
    wire signal_10125 ;
    wire signal_10126 ;
    wire signal_10127 ;
    wire signal_10128 ;
    wire signal_10129 ;
    wire signal_10130 ;
    wire signal_10131 ;
    wire signal_10132 ;
    wire signal_10133 ;
    wire signal_10134 ;
    wire signal_10135 ;
    wire signal_10136 ;
    wire signal_10137 ;
    wire signal_10138 ;
    wire signal_10139 ;
    wire signal_10140 ;
    wire signal_10141 ;
    wire signal_10142 ;
    wire signal_10143 ;
    wire signal_10144 ;
    wire signal_10145 ;
    wire signal_10146 ;
    wire signal_10147 ;
    wire signal_10148 ;
    wire signal_10149 ;
    wire signal_10150 ;
    wire signal_10151 ;
    wire signal_10152 ;
    wire signal_10153 ;
    wire signal_10154 ;
    wire signal_10155 ;
    wire signal_10156 ;
    wire signal_10157 ;
    wire signal_10158 ;
    wire signal_10159 ;
    wire signal_10160 ;
    wire signal_10161 ;
    wire signal_10162 ;
    wire signal_10163 ;
    wire signal_10164 ;
    wire signal_10165 ;
    wire signal_10166 ;
    wire signal_10167 ;
    wire signal_10168 ;
    wire signal_10169 ;
    wire signal_10170 ;
    wire signal_10171 ;
    wire signal_10172 ;
    wire signal_10173 ;
    wire signal_10174 ;
    wire signal_10175 ;
    wire signal_10176 ;
    wire signal_10177 ;
    wire signal_10178 ;
    wire signal_10179 ;
    wire signal_10180 ;
    wire signal_10181 ;
    wire signal_10182 ;
    wire signal_10183 ;
    wire signal_10184 ;
    wire signal_10185 ;
    wire signal_10186 ;
    wire signal_10187 ;
    wire signal_10188 ;
    wire signal_10189 ;
    wire signal_10190 ;
    wire signal_10191 ;
    wire signal_10192 ;
    wire signal_10193 ;
    wire signal_10194 ;
    wire signal_10195 ;
    wire signal_10196 ;
    wire signal_10197 ;
    wire signal_10198 ;
    wire signal_10199 ;
    wire signal_10200 ;
    wire signal_10201 ;
    wire signal_10202 ;
    wire signal_10203 ;
    wire signal_10204 ;
    wire signal_10205 ;
    wire signal_10206 ;
    wire signal_10207 ;
    wire signal_10208 ;
    wire signal_10209 ;
    wire signal_10210 ;
    wire signal_10211 ;
    wire signal_10212 ;
    wire signal_10213 ;
    wire signal_10214 ;
    wire signal_10215 ;
    wire signal_10216 ;
    wire signal_10217 ;
    wire signal_10218 ;
    wire signal_10219 ;
    wire signal_10220 ;
    wire signal_10221 ;
    wire signal_10222 ;
    wire signal_10223 ;
    wire signal_10224 ;
    wire signal_10225 ;
    wire signal_10226 ;
    wire signal_10227 ;
    wire signal_10228 ;
    wire signal_10229 ;
    wire signal_10230 ;
    wire signal_10231 ;
    wire signal_10232 ;
    wire signal_10233 ;
    wire signal_10234 ;
    wire signal_10235 ;
    wire signal_10236 ;
    wire signal_10237 ;
    wire signal_10238 ;
    wire signal_10239 ;
    wire signal_10240 ;
    wire signal_10241 ;
    wire signal_10242 ;
    wire signal_10243 ;
    wire signal_10244 ;
    wire signal_10245 ;
    wire signal_10246 ;
    wire signal_10247 ;
    wire signal_10248 ;
    wire signal_10249 ;
    wire signal_10250 ;
    wire signal_10251 ;
    wire signal_10252 ;
    wire signal_10253 ;
    wire signal_10254 ;
    wire signal_10255 ;
    wire signal_10256 ;
    wire signal_10257 ;
    wire signal_10258 ;
    wire signal_10259 ;
    wire signal_10260 ;
    wire signal_10261 ;
    wire signal_10262 ;
    wire signal_10263 ;
    wire signal_10264 ;
    wire signal_10265 ;
    wire signal_10266 ;
    wire signal_10267 ;
    wire signal_10268 ;
    wire signal_10269 ;
    wire signal_10270 ;
    wire signal_10271 ;
    wire signal_10272 ;
    wire signal_10273 ;
    wire signal_10274 ;
    wire signal_10275 ;
    wire signal_10276 ;
    wire signal_10277 ;
    wire signal_10278 ;
    wire signal_10279 ;
    wire signal_10280 ;
    wire signal_10281 ;
    wire signal_10282 ;
    wire signal_10283 ;
    wire signal_10284 ;
    wire signal_10285 ;
    wire signal_10286 ;
    wire signal_10287 ;
    wire signal_10288 ;
    wire signal_10289 ;
    wire signal_10290 ;
    wire signal_10291 ;
    wire signal_10292 ;
    wire signal_10293 ;
    wire signal_10294 ;
    wire signal_10295 ;
    wire signal_10296 ;
    wire signal_10297 ;
    wire signal_10298 ;
    wire signal_10299 ;
    wire signal_10300 ;
    wire signal_10301 ;
    wire signal_10302 ;
    wire signal_10303 ;
    wire signal_10304 ;
    wire signal_10305 ;
    wire signal_10306 ;
    wire signal_10307 ;
    wire signal_10308 ;
    wire signal_10309 ;
    wire signal_10310 ;
    wire signal_10311 ;
    wire signal_10312 ;
    wire signal_10313 ;
    wire signal_10314 ;
    wire signal_10315 ;
    wire signal_10316 ;
    wire signal_10317 ;
    wire signal_10318 ;
    wire signal_10319 ;
    wire signal_10320 ;
    wire signal_10321 ;
    wire signal_10322 ;
    wire signal_10323 ;
    wire signal_10324 ;
    wire signal_10325 ;
    wire signal_10326 ;
    wire signal_10327 ;
    wire signal_10328 ;
    wire signal_10329 ;
    wire signal_10330 ;
    wire signal_10331 ;
    wire signal_10332 ;
    wire signal_10333 ;
    wire signal_10334 ;
    wire signal_10335 ;
    wire signal_10336 ;
    wire signal_10337 ;
    wire signal_10338 ;
    wire signal_10339 ;
    wire signal_10340 ;
    wire signal_10341 ;
    wire signal_10342 ;
    wire signal_10343 ;
    wire signal_10344 ;
    wire signal_10345 ;
    wire signal_10346 ;
    wire signal_10347 ;
    wire signal_10348 ;
    wire signal_10349 ;
    wire signal_10350 ;
    wire signal_10351 ;
    wire signal_10352 ;
    wire signal_10353 ;
    wire signal_10354 ;
    wire signal_10355 ;
    wire signal_10356 ;
    wire signal_10357 ;
    wire signal_10358 ;
    wire signal_10359 ;
    wire signal_10360 ;
    wire signal_10361 ;
    wire signal_10362 ;
    wire signal_10363 ;
    wire signal_10364 ;
    wire signal_10365 ;
    wire signal_10366 ;
    wire signal_10367 ;
    wire signal_10368 ;
    wire signal_10369 ;
    wire signal_10370 ;
    wire signal_10371 ;
    wire signal_10372 ;
    wire signal_10373 ;
    wire signal_10374 ;
    wire signal_10375 ;
    wire signal_10376 ;
    wire signal_10377 ;
    wire signal_10378 ;
    wire signal_10379 ;
    wire signal_10380 ;
    wire signal_10381 ;
    wire signal_10382 ;
    wire signal_10383 ;
    wire signal_10384 ;
    wire signal_10385 ;
    wire signal_10386 ;
    wire signal_10387 ;
    wire signal_10388 ;
    wire signal_10389 ;
    wire signal_10390 ;
    wire signal_10391 ;
    wire signal_10392 ;
    wire signal_10393 ;
    wire signal_10394 ;
    wire signal_10395 ;
    wire signal_10396 ;
    wire signal_10397 ;
    wire signal_10398 ;
    wire signal_10399 ;
    wire signal_10400 ;
    wire signal_10401 ;
    wire signal_10402 ;
    wire signal_10403 ;
    wire signal_10404 ;
    wire signal_10405 ;
    wire signal_10406 ;
    wire signal_10407 ;
    wire signal_10408 ;
    wire signal_10409 ;
    wire signal_10410 ;
    wire signal_10411 ;
    wire signal_10412 ;
    wire signal_10413 ;
    wire signal_10414 ;
    wire signal_10415 ;
    wire signal_10416 ;
    wire signal_10417 ;
    wire signal_10418 ;
    wire signal_10419 ;
    wire signal_10420 ;
    wire signal_10421 ;
    wire signal_10422 ;
    wire signal_10423 ;
    wire signal_10424 ;
    wire signal_10425 ;
    wire signal_10426 ;
    wire signal_10427 ;
    wire signal_10428 ;
    wire signal_10429 ;
    wire signal_10430 ;
    wire signal_10431 ;
    wire signal_10432 ;
    wire signal_10433 ;
    wire signal_10434 ;
    wire signal_10435 ;
    wire signal_10436 ;
    wire signal_10437 ;
    wire signal_10438 ;
    wire signal_10439 ;
    wire signal_10440 ;
    wire signal_10441 ;
    wire signal_10442 ;
    wire signal_10443 ;
    wire signal_10444 ;
    wire signal_10445 ;
    wire signal_10446 ;
    wire signal_10447 ;
    wire signal_10448 ;
    wire signal_10449 ;
    wire signal_10450 ;
    wire signal_10451 ;
    wire signal_10452 ;
    wire signal_10453 ;
    wire signal_10454 ;
    wire signal_10455 ;
    wire signal_10457 ;
    wire signal_10459 ;
    wire signal_10461 ;
    wire signal_10463 ;
    wire signal_10465 ;
    wire signal_10467 ;
    wire signal_10469 ;
    wire signal_10471 ;
    wire signal_10473 ;
    wire signal_10475 ;
    wire signal_10477 ;
    wire signal_10479 ;
    wire signal_10481 ;
    wire signal_10483 ;
    wire signal_10485 ;
    wire signal_10486 ;
    wire signal_10487 ;
    wire signal_10488 ;
    wire signal_10489 ;
    wire signal_10490 ;
    wire signal_10491 ;
    wire signal_10492 ;
    wire signal_10493 ;
    wire signal_10494 ;
    wire signal_10495 ;
    wire signal_10496 ;
    wire signal_10497 ;
    wire signal_10498 ;
    wire signal_10499 ;
    wire signal_10500 ;
    wire signal_10501 ;
    wire signal_10502 ;
    wire signal_10503 ;
    wire signal_10504 ;
    wire signal_10505 ;
    wire signal_10506 ;
    wire signal_10507 ;
    wire signal_10508 ;
    wire signal_10509 ;
    wire signal_10510 ;
    wire signal_10511 ;
    wire signal_10512 ;
    wire signal_10513 ;
    wire signal_10514 ;
    wire signal_10515 ;
    wire signal_10516 ;
    wire signal_10517 ;
    wire signal_10518 ;
    wire signal_10519 ;
    wire signal_10520 ;
    wire signal_10521 ;
    wire signal_10522 ;
    wire signal_10523 ;
    wire signal_10524 ;
    wire signal_10525 ;
    wire signal_10526 ;
    wire signal_10527 ;
    wire signal_10528 ;
    wire signal_10529 ;
    wire signal_10530 ;
    wire signal_10531 ;
    wire signal_10532 ;
    wire signal_10533 ;
    wire signal_10534 ;
    wire signal_10535 ;
    wire signal_10536 ;
    wire signal_10537 ;
    wire signal_10538 ;
    wire signal_10539 ;
    wire signal_10540 ;
    wire signal_10541 ;
    wire signal_10542 ;
    wire signal_10543 ;
    wire signal_10544 ;
    wire signal_10545 ;
    wire signal_10546 ;
    wire signal_10547 ;
    wire signal_10548 ;
    wire signal_10549 ;
    wire signal_10550 ;
    wire signal_10551 ;
    wire signal_10552 ;
    wire signal_10553 ;
    wire signal_10554 ;
    wire signal_10555 ;
    wire signal_10556 ;
    wire signal_10557 ;
    wire signal_10558 ;
    wire signal_10559 ;
    wire signal_10560 ;
    wire signal_10561 ;
    wire signal_10562 ;
    wire signal_10563 ;
    wire signal_10564 ;
    wire signal_10565 ;
    wire signal_10566 ;
    wire signal_10567 ;
    wire signal_10568 ;
    wire signal_10569 ;
    wire signal_10570 ;
    wire signal_10571 ;
    wire signal_10572 ;
    wire signal_10573 ;
    wire signal_10574 ;
    wire signal_10575 ;
    wire signal_10576 ;
    wire signal_10577 ;
    wire signal_10578 ;
    wire signal_10579 ;
    wire signal_10580 ;
    wire signal_10581 ;
    wire signal_10582 ;
    wire signal_10583 ;
    wire signal_10584 ;
    wire signal_10585 ;
    wire signal_10586 ;
    wire signal_10587 ;
    wire signal_10588 ;
    wire signal_10589 ;
    wire signal_10590 ;
    wire signal_10591 ;
    wire signal_10592 ;
    wire signal_10593 ;
    wire signal_10594 ;
    wire signal_10595 ;
    wire signal_10596 ;
    wire signal_10597 ;
    wire signal_10598 ;
    wire signal_10599 ;
    wire signal_10600 ;
    wire signal_10601 ;
    wire signal_10602 ;
    wire signal_10603 ;
    wire signal_10604 ;
    wire signal_10605 ;
    wire signal_10606 ;
    wire signal_10607 ;
    wire signal_10608 ;
    wire signal_10609 ;
    wire signal_10610 ;
    wire signal_10611 ;
    wire signal_10612 ;
    wire signal_10613 ;
    wire signal_10614 ;
    wire signal_10615 ;
    wire signal_10616 ;
    wire signal_10617 ;
    wire signal_10618 ;
    wire signal_10619 ;
    wire signal_10620 ;
    wire signal_10621 ;
    wire signal_10622 ;
    wire signal_10623 ;
    wire signal_10624 ;
    wire signal_10625 ;
    wire signal_10626 ;
    wire signal_10627 ;
    wire signal_10628 ;
    wire signal_10629 ;
    wire signal_10630 ;
    wire signal_10631 ;
    wire signal_10632 ;
    wire signal_10633 ;
    wire signal_10634 ;
    wire signal_10635 ;
    wire signal_10636 ;
    wire signal_10637 ;
    wire signal_10638 ;
    wire signal_10639 ;
    wire signal_10640 ;
    wire signal_10641 ;
    wire signal_10642 ;
    wire signal_10643 ;
    wire signal_10644 ;
    wire signal_10645 ;
    wire signal_10646 ;
    wire signal_10647 ;
    wire signal_10648 ;
    wire signal_10649 ;
    wire signal_10650 ;
    wire signal_10651 ;
    wire signal_10652 ;
    wire signal_10653 ;
    wire signal_10654 ;
    wire signal_10655 ;
    wire signal_10656 ;
    wire signal_10657 ;
    wire signal_10658 ;
    wire signal_10659 ;
    wire signal_10660 ;
    wire signal_10661 ;
    wire signal_10662 ;
    wire signal_10663 ;
    wire signal_10664 ;
    wire signal_10665 ;
    wire signal_10666 ;
    wire signal_10667 ;
    wire signal_10668 ;
    wire signal_10669 ;
    wire signal_10670 ;
    wire signal_10671 ;
    wire signal_10672 ;
    wire signal_10673 ;
    wire signal_10674 ;
    wire signal_10675 ;
    wire signal_10676 ;
    wire signal_10677 ;
    wire signal_10678 ;
    wire signal_10679 ;
    wire signal_10680 ;
    wire signal_10681 ;
    wire signal_10682 ;
    wire signal_10683 ;
    wire signal_10684 ;
    wire signal_10685 ;
    wire signal_10686 ;
    wire signal_10687 ;
    wire signal_10688 ;
    wire signal_10689 ;
    wire signal_10690 ;
    wire signal_10691 ;
    wire signal_10692 ;
    wire signal_10693 ;
    wire signal_10694 ;
    wire signal_10695 ;
    wire signal_10696 ;
    wire signal_10697 ;
    wire signal_10698 ;
    wire signal_10699 ;
    wire signal_10700 ;
    wire signal_10701 ;
    wire signal_10702 ;
    wire signal_10703 ;
    wire signal_10704 ;
    wire signal_10705 ;
    wire signal_10707 ;
    wire signal_10709 ;
    wire signal_10711 ;
    wire signal_10713 ;
    wire signal_10715 ;
    wire signal_10717 ;
    wire signal_10719 ;
    wire signal_10721 ;
    wire signal_10723 ;
    wire signal_10725 ;
    wire signal_10727 ;
    wire signal_10729 ;
    wire signal_10731 ;
    wire signal_10733 ;
    wire signal_10735 ;
    wire signal_10737 ;
    wire signal_10739 ;
    wire signal_10741 ;
    wire signal_10743 ;
    wire signal_10745 ;
    wire signal_10747 ;
    wire signal_10749 ;
    wire signal_10751 ;
    wire signal_10753 ;
    wire signal_10755 ;
    wire signal_10757 ;
    wire signal_10759 ;
    wire signal_10761 ;
    wire signal_10763 ;
    wire signal_10764 ;
    wire signal_10765 ;
    wire signal_10766 ;
    wire signal_10767 ;
    wire signal_10768 ;
    wire signal_10769 ;
    wire signal_10770 ;
    wire signal_10771 ;
    wire signal_10772 ;
    wire signal_10773 ;
    wire signal_10774 ;
    wire signal_10775 ;
    wire signal_10776 ;
    wire signal_10777 ;
    wire signal_10778 ;
    wire signal_10779 ;
    wire signal_10780 ;
    wire signal_10781 ;
    wire signal_10782 ;
    wire signal_10783 ;
    wire signal_10784 ;
    wire signal_10785 ;
    wire signal_10786 ;
    wire signal_10787 ;
    wire signal_10788 ;
    wire signal_10789 ;
    wire signal_10790 ;
    wire signal_10791 ;
    wire signal_10792 ;
    wire signal_10793 ;
    wire signal_10794 ;
    wire signal_10795 ;
    wire signal_10796 ;
    wire signal_10797 ;
    wire signal_10798 ;
    wire signal_10799 ;
    wire signal_10800 ;
    wire signal_10801 ;
    wire signal_10802 ;
    wire signal_10803 ;
    wire signal_10804 ;
    wire signal_10805 ;
    wire signal_10806 ;
    wire signal_10807 ;
    wire signal_10808 ;
    wire signal_10809 ;
    wire signal_10810 ;
    wire signal_10811 ;
    wire signal_10812 ;
    wire signal_10813 ;
    wire signal_10814 ;
    wire signal_10815 ;
    wire signal_10816 ;
    wire signal_10817 ;
    wire signal_10818 ;
    wire signal_10819 ;
    wire signal_10820 ;
    wire signal_10821 ;
    wire signal_10822 ;
    wire signal_10823 ;
    wire signal_10824 ;
    wire signal_10825 ;
    wire signal_10826 ;
    wire signal_10827 ;
    wire signal_10828 ;
    wire signal_10829 ;
    wire signal_10830 ;
    wire signal_10831 ;
    wire signal_10832 ;
    wire signal_10833 ;
    wire signal_10834 ;
    wire signal_10835 ;
    wire signal_10836 ;
    wire signal_10837 ;
    wire signal_10838 ;
    wire signal_10839 ;
    wire signal_10840 ;
    wire signal_10841 ;
    wire signal_10842 ;
    wire signal_10843 ;
    wire signal_10844 ;
    wire signal_10845 ;
    wire signal_10846 ;
    wire signal_10847 ;
    wire signal_10848 ;
    wire signal_10849 ;
    wire signal_10850 ;
    wire signal_10851 ;
    wire signal_10852 ;
    wire signal_10853 ;
    wire signal_10854 ;
    wire signal_10855 ;
    wire signal_10856 ;
    wire signal_10857 ;
    wire signal_10858 ;
    wire signal_10859 ;
    wire signal_10860 ;
    wire signal_10861 ;
    wire signal_10862 ;
    wire signal_10863 ;
    wire signal_10864 ;
    wire signal_10865 ;
    wire signal_10866 ;
    wire signal_10867 ;
    wire signal_10868 ;
    wire signal_10869 ;
    wire signal_10870 ;
    wire signal_10871 ;
    wire signal_10872 ;
    wire signal_10873 ;
    wire signal_10874 ;
    wire signal_10875 ;
    wire signal_10876 ;
    wire signal_10877 ;
    wire signal_10878 ;
    wire signal_10879 ;
    wire signal_10880 ;
    wire signal_10881 ;
    wire signal_10882 ;
    wire signal_10883 ;
    wire signal_10884 ;
    wire signal_10885 ;
    wire signal_10886 ;
    wire signal_10887 ;
    wire signal_10888 ;
    wire signal_10889 ;
    wire signal_10890 ;
    wire signal_10891 ;
    wire signal_10892 ;
    wire signal_10893 ;
    wire signal_10894 ;
    wire signal_10895 ;
    wire signal_10896 ;
    wire signal_10897 ;
    wire signal_10898 ;
    wire signal_10899 ;
    wire signal_10900 ;
    wire signal_10901 ;
    wire signal_10902 ;
    wire signal_10903 ;
    wire signal_10904 ;
    wire signal_10905 ;
    wire signal_10906 ;
    wire signal_10907 ;
    wire signal_10908 ;
    wire signal_10909 ;
    wire signal_10910 ;
    wire signal_10911 ;
    wire signal_10912 ;
    wire signal_10913 ;
    wire signal_10914 ;
    wire signal_10915 ;
    wire signal_10916 ;
    wire signal_10917 ;
    wire signal_10918 ;
    wire signal_10919 ;
    wire signal_10920 ;
    wire signal_10921 ;
    wire signal_10922 ;
    wire signal_10923 ;
    wire signal_10924 ;
    wire signal_10925 ;
    wire signal_10926 ;
    wire signal_10927 ;
    wire signal_10928 ;
    wire signal_10929 ;
    wire signal_10930 ;
    wire signal_10931 ;
    wire signal_10932 ;
    wire signal_10933 ;
    wire signal_10934 ;
    wire signal_10935 ;
    wire signal_10937 ;
    wire signal_10939 ;
    wire signal_10941 ;
    wire signal_10943 ;
    wire signal_10945 ;
    wire signal_10947 ;
    wire signal_10949 ;
    wire signal_10951 ;
    wire signal_10953 ;
    wire signal_10955 ;
    wire signal_10957 ;
    wire signal_10959 ;
    wire signal_10961 ;
    wire signal_10963 ;
    wire signal_10965 ;
    wire signal_10967 ;
    wire signal_10969 ;
    wire signal_10971 ;
    wire signal_10973 ;
    wire signal_10975 ;
    wire signal_10977 ;
    wire signal_10979 ;
    wire signal_10981 ;
    wire signal_10983 ;
    wire signal_10985 ;
    wire signal_10987 ;
    wire signal_10989 ;
    wire signal_10991 ;
    wire signal_10993 ;
    wire signal_10995 ;
    wire signal_10997 ;
    wire signal_10999 ;
    wire signal_11000 ;
    wire signal_11001 ;
    wire signal_11002 ;
    wire signal_11003 ;
    wire signal_11004 ;
    wire signal_11005 ;
    wire signal_11006 ;
    wire signal_11007 ;
    wire signal_11008 ;
    wire signal_11009 ;
    wire signal_11010 ;
    wire signal_11011 ;
    wire signal_11012 ;
    wire signal_11013 ;
    wire signal_11014 ;
    wire signal_11015 ;
    wire signal_11016 ;
    wire signal_11017 ;
    wire signal_11018 ;
    wire signal_11019 ;
    wire signal_11020 ;
    wire signal_11021 ;
    wire signal_11022 ;
    wire signal_11023 ;
    wire signal_11024 ;
    wire signal_11025 ;
    wire signal_11026 ;
    wire signal_11027 ;
    wire signal_11028 ;
    wire signal_11029 ;
    wire signal_11030 ;
    wire signal_11031 ;
    wire signal_11032 ;
    wire signal_11033 ;
    wire signal_11034 ;
    wire signal_11035 ;
    wire signal_11036 ;
    wire signal_11037 ;
    wire signal_11038 ;
    wire signal_11039 ;
    wire signal_11040 ;
    wire signal_11041 ;
    wire signal_11042 ;
    wire signal_11043 ;
    wire signal_11044 ;
    wire signal_11045 ;
    wire signal_11046 ;
    wire signal_11047 ;
    wire signal_11048 ;
    wire signal_11049 ;
    wire signal_11050 ;
    wire signal_11051 ;
    wire signal_11052 ;
    wire signal_11053 ;
    wire signal_11054 ;
    wire signal_11055 ;
    wire signal_11056 ;
    wire signal_11057 ;
    wire signal_11058 ;
    wire signal_11059 ;
    wire signal_11060 ;
    wire signal_11061 ;
    wire signal_11062 ;
    wire signal_11063 ;
    wire signal_11064 ;
    wire signal_11065 ;
    wire signal_11066 ;
    wire signal_11067 ;
    wire signal_11068 ;
    wire signal_11069 ;
    wire signal_11070 ;
    wire signal_11071 ;
    wire signal_11072 ;
    wire signal_11073 ;
    wire signal_11074 ;
    wire signal_11075 ;
    wire signal_11076 ;
    wire signal_11077 ;
    wire signal_11078 ;
    wire signal_11079 ;
    wire signal_11080 ;
    wire signal_11081 ;
    wire signal_11082 ;
    wire signal_11083 ;
    wire signal_11084 ;
    wire signal_11085 ;
    wire signal_11086 ;
    wire signal_11087 ;
    wire signal_11088 ;
    wire signal_11089 ;
    wire signal_11090 ;
    wire signal_11091 ;
    wire signal_11092 ;
    wire signal_11093 ;
    wire signal_11094 ;
    wire signal_11095 ;
    wire signal_11096 ;
    wire signal_11097 ;
    wire signal_11098 ;
    wire signal_11099 ;
    wire signal_11100 ;
    wire signal_11101 ;
    wire signal_11102 ;
    wire signal_11103 ;
    wire signal_11104 ;
    wire signal_11105 ;
    wire signal_11106 ;
    wire signal_11107 ;
    wire signal_11108 ;
    wire signal_11109 ;
    wire signal_11110 ;
    wire signal_11111 ;
    wire signal_11112 ;
    wire signal_11113 ;
    wire signal_11114 ;
    wire signal_11115 ;
    wire signal_11116 ;
    wire signal_11117 ;
    wire signal_11118 ;
    wire signal_11119 ;
    wire signal_11120 ;
    wire signal_11121 ;
    wire signal_11122 ;
    wire signal_11123 ;
    wire signal_11124 ;
    wire signal_11125 ;
    wire signal_11126 ;
    wire signal_11127 ;
    wire signal_11128 ;
    wire signal_11129 ;
    wire signal_11130 ;
    wire signal_11131 ;
    wire signal_11132 ;
    wire signal_11133 ;
    wire signal_11134 ;
    wire signal_11135 ;
    wire signal_11136 ;
    wire signal_11137 ;
    wire signal_11138 ;
    wire signal_11139 ;
    wire signal_11140 ;
    wire signal_11141 ;
    wire signal_11142 ;
    wire signal_11143 ;
    wire signal_11144 ;
    wire signal_11145 ;
    wire signal_11146 ;
    wire signal_11147 ;
    wire signal_11148 ;
    wire signal_11149 ;
    wire signal_11150 ;
    wire signal_11151 ;
    wire signal_11152 ;
    wire signal_11153 ;
    wire signal_11154 ;
    wire signal_11155 ;
    wire signal_11156 ;
    wire signal_11157 ;
    wire signal_11158 ;
    wire signal_11159 ;
    wire signal_11160 ;
    wire signal_11161 ;
    wire signal_11162 ;
    wire signal_11163 ;
    wire signal_11164 ;
    wire signal_11165 ;
    wire signal_11166 ;
    wire signal_11167 ;
    wire signal_11168 ;
    wire signal_11169 ;
    wire signal_11170 ;
    wire signal_11171 ;
    wire signal_11172 ;
    wire signal_11173 ;
    wire signal_11174 ;
    wire signal_11175 ;
    wire signal_11176 ;
    wire signal_11177 ;
    wire signal_11178 ;
    wire signal_11179 ;
    wire signal_11180 ;
    wire signal_11181 ;
    wire signal_11182 ;
    wire signal_11183 ;
    wire signal_11184 ;
    wire signal_11185 ;
    wire signal_11186 ;
    wire signal_11187 ;
    wire signal_11188 ;
    wire signal_11189 ;
    wire signal_11190 ;
    wire signal_11191 ;
    wire signal_11192 ;
    wire signal_11193 ;
    wire signal_11194 ;
    wire signal_11195 ;
    wire signal_11196 ;
    wire signal_11197 ;
    wire signal_11198 ;
    wire signal_11199 ;
    wire signal_11200 ;
    wire signal_11202 ;
    wire signal_11204 ;
    wire signal_11206 ;
    wire signal_11208 ;
    wire signal_11210 ;
    wire signal_11212 ;
    wire signal_11214 ;
    wire signal_11216 ;
    wire signal_11218 ;
    wire signal_11220 ;
    wire signal_11222 ;
    wire signal_11224 ;
    wire signal_11226 ;
    wire signal_11228 ;
    wire signal_11230 ;
    wire signal_11232 ;
    wire signal_11234 ;
    wire signal_11236 ;
    wire signal_11238 ;
    wire signal_11240 ;
    wire signal_11242 ;
    wire signal_11244 ;
    wire signal_11246 ;
    wire signal_11248 ;
    wire signal_11250 ;
    wire signal_11252 ;
    wire signal_11254 ;
    wire signal_11256 ;
    wire signal_11258 ;
    wire signal_11260 ;
    wire signal_11262 ;
    wire signal_11264 ;
    wire signal_11265 ;
    wire signal_11266 ;
    wire signal_11267 ;
    wire signal_11268 ;
    wire signal_11269 ;
    wire signal_11270 ;
    wire signal_11271 ;
    wire signal_11272 ;
    wire signal_11273 ;
    wire signal_11274 ;
    wire signal_11275 ;
    wire signal_11276 ;
    wire signal_11277 ;
    wire signal_11278 ;
    wire signal_11279 ;
    wire signal_11280 ;
    wire signal_11281 ;
    wire signal_11282 ;
    wire signal_11283 ;
    wire signal_11284 ;
    wire signal_11285 ;
    wire signal_11286 ;
    wire signal_11287 ;
    wire signal_11288 ;
    wire signal_11289 ;
    wire signal_11290 ;
    wire signal_11291 ;
    wire signal_11292 ;
    wire signal_11293 ;
    wire signal_11294 ;
    wire signal_11295 ;
    wire signal_11296 ;
    wire signal_11297 ;
    wire signal_11298 ;
    wire signal_11299 ;
    wire signal_11300 ;
    wire signal_11301 ;
    wire signal_11302 ;
    wire signal_11303 ;
    wire signal_11304 ;
    wire signal_11305 ;
    wire signal_11306 ;
    wire signal_11307 ;
    wire signal_11308 ;
    wire signal_11309 ;
    wire signal_11310 ;
    wire signal_11311 ;
    wire signal_11312 ;
    wire signal_11313 ;
    wire signal_11314 ;
    wire signal_11315 ;
    wire signal_11316 ;
    wire signal_11317 ;
    wire signal_11318 ;
    wire signal_11319 ;
    wire signal_11320 ;
    wire signal_11321 ;
    wire signal_11322 ;
    wire signal_11323 ;
    wire signal_11324 ;
    wire signal_11325 ;
    wire signal_11326 ;
    wire signal_11327 ;
    wire signal_11328 ;
    wire signal_11329 ;
    wire signal_11330 ;
    wire signal_11331 ;
    wire signal_11332 ;
    wire signal_11333 ;
    wire signal_11334 ;
    wire signal_11335 ;
    wire signal_11336 ;
    wire signal_11337 ;
    wire signal_11338 ;
    wire signal_11339 ;
    wire signal_11340 ;
    wire signal_11341 ;
    wire signal_11342 ;
    wire signal_11343 ;
    wire signal_11344 ;
    wire signal_11345 ;
    wire signal_11346 ;
    wire signal_11347 ;
    wire signal_11348 ;
    wire signal_11349 ;
    wire signal_11350 ;
    wire signal_11351 ;
    wire signal_11352 ;
    wire signal_11353 ;
    wire signal_11354 ;
    wire signal_11355 ;
    wire signal_11356 ;
    wire signal_11357 ;
    wire signal_11358 ;
    wire signal_11359 ;
    wire signal_11360 ;
    wire signal_11361 ;
    wire signal_11362 ;
    wire signal_11363 ;
    wire signal_11364 ;
    wire signal_11365 ;
    wire signal_11366 ;
    wire signal_11367 ;
    wire signal_11368 ;
    wire signal_11369 ;
    wire signal_11370 ;
    wire signal_11371 ;
    wire signal_11372 ;
    wire signal_11373 ;
    wire signal_11374 ;
    wire signal_11375 ;
    wire signal_11376 ;
    wire signal_11377 ;
    wire signal_11378 ;
    wire signal_11379 ;
    wire signal_11380 ;
    wire signal_11381 ;
    wire signal_11382 ;
    wire signal_11383 ;
    wire signal_11384 ;
    wire signal_11385 ;
    wire signal_11386 ;
    wire signal_11387 ;
    wire signal_11388 ;
    wire signal_11389 ;
    wire signal_11390 ;
    wire signal_11391 ;
    wire signal_11392 ;
    wire signal_11393 ;
    wire signal_11394 ;
    wire signal_11395 ;
    wire signal_11396 ;
    wire signal_11397 ;
    wire signal_11398 ;
    wire signal_11399 ;
    wire signal_11400 ;
    wire signal_11401 ;
    wire signal_11402 ;
    wire signal_11403 ;
    wire signal_11404 ;
    wire signal_11405 ;
    wire signal_11406 ;
    wire signal_11407 ;
    wire signal_11408 ;
    wire signal_11409 ;
    wire signal_11410 ;
    wire signal_11411 ;
    wire signal_11412 ;
    wire signal_11413 ;
    wire signal_11414 ;
    wire signal_11415 ;
    wire signal_11416 ;
    wire signal_11417 ;
    wire signal_11418 ;
    wire signal_11419 ;
    wire signal_11420 ;
    wire signal_11421 ;
    wire signal_11422 ;
    wire signal_11423 ;
    wire signal_11424 ;
    wire signal_11425 ;
    wire signal_11426 ;
    wire signal_11427 ;
    wire signal_11428 ;
    wire signal_11429 ;
    wire signal_11430 ;
    wire signal_11431 ;
    wire signal_11432 ;
    wire signal_11433 ;
    wire signal_11434 ;
    wire signal_11435 ;
    wire signal_11436 ;
    wire signal_11437 ;
    wire signal_11438 ;
    wire signal_11439 ;
    wire signal_11440 ;
    wire signal_11441 ;
    wire signal_11442 ;
    wire signal_11443 ;
    wire signal_11444 ;
    wire signal_11445 ;
    wire signal_11446 ;
    wire signal_11447 ;
    wire signal_11448 ;
    wire signal_11449 ;
    wire signal_11450 ;
    wire signal_11451 ;
    wire signal_11452 ;
    wire signal_11453 ;
    wire signal_11454 ;
    wire signal_11455 ;
    wire signal_11456 ;
    wire signal_11457 ;
    wire signal_11459 ;
    wire signal_11461 ;
    wire signal_11463 ;
    wire signal_11465 ;
    wire signal_11467 ;
    wire signal_11469 ;
    wire signal_11471 ;
    wire signal_11473 ;
    wire signal_11475 ;
    wire signal_11477 ;
    wire signal_11479 ;
    wire signal_11481 ;
    wire signal_11483 ;
    wire signal_11485 ;
    wire signal_11487 ;
    wire signal_11489 ;
    wire signal_11491 ;
    wire signal_11493 ;
    wire signal_11495 ;
    wire signal_11497 ;
    wire signal_11499 ;
    wire signal_11501 ;
    wire signal_11503 ;
    wire signal_11505 ;
    wire signal_11507 ;
    wire signal_11509 ;
    wire signal_11511 ;
    wire signal_11513 ;
    wire signal_11515 ;
    wire signal_11517 ;
    wire signal_11519 ;
    wire signal_11521 ;
    wire signal_11523 ;
    wire signal_11525 ;
    wire signal_11527 ;
    wire signal_11529 ;
    wire signal_11531 ;
    wire signal_11533 ;
    wire signal_11535 ;
    wire signal_11537 ;
    wire signal_11539 ;
    wire signal_11541 ;
    wire signal_11543 ;
    wire signal_11545 ;
    wire signal_11547 ;
    wire signal_11549 ;
    wire signal_11551 ;
    wire signal_11553 ;
    wire signal_11555 ;
    wire signal_11556 ;
    wire signal_11557 ;
    wire signal_11558 ;
    wire signal_11559 ;
    wire signal_11560 ;
    wire signal_11561 ;
    wire signal_11562 ;
    wire signal_11563 ;
    wire signal_11564 ;
    wire signal_11565 ;
    wire signal_11566 ;
    wire signal_11567 ;
    wire signal_11568 ;
    wire signal_11569 ;
    wire signal_11570 ;
    wire signal_11571 ;
    wire signal_11572 ;
    wire signal_11573 ;
    wire signal_11574 ;
    wire signal_11575 ;
    wire signal_11576 ;
    wire signal_11577 ;
    wire signal_11578 ;
    wire signal_11579 ;
    wire signal_11580 ;
    wire signal_11581 ;
    wire signal_11582 ;
    wire signal_11583 ;
    wire signal_11584 ;
    wire signal_11585 ;
    wire signal_11586 ;
    wire signal_11587 ;
    wire signal_11588 ;
    wire signal_11589 ;
    wire signal_11590 ;
    wire signal_11592 ;
    wire signal_11594 ;
    wire signal_11596 ;
    wire signal_11598 ;
    wire signal_11600 ;
    wire signal_11602 ;
    wire signal_11604 ;
    wire signal_11606 ;
    wire signal_11608 ;
    wire signal_11610 ;
    wire signal_11612 ;
    wire signal_11614 ;
    wire signal_11616 ;
    wire signal_11618 ;
    wire signal_11620 ;
    wire signal_11622 ;
    wire signal_11624 ;
    wire signal_11626 ;
    wire signal_11628 ;
    wire signal_11630 ;
    wire signal_11632 ;
    wire signal_11634 ;
    wire signal_11636 ;
    wire signal_11638 ;
    wire signal_11640 ;
    wire signal_11642 ;
    wire signal_11644 ;
    wire signal_11646 ;
    wire signal_11648 ;
    wire signal_11650 ;
    wire signal_11652 ;
    wire signal_11654 ;
    wire signal_11656 ;
    wire signal_11658 ;
    wire signal_11660 ;
    wire signal_11662 ;
    wire signal_11664 ;
    wire signal_11666 ;
    wire signal_11668 ;
    wire signal_11670 ;
    wire signal_11672 ;
    wire signal_11674 ;
    wire signal_11676 ;
    wire signal_11678 ;
    wire signal_11680 ;
    wire signal_11682 ;
    wire signal_11684 ;
    wire signal_11686 ;
    wire signal_11688 ;
    wire signal_11690 ;
    wire signal_11692 ;
    wire signal_11694 ;
    wire signal_11696 ;
    wire signal_11698 ;
    wire signal_11700 ;
    wire signal_11702 ;
    wire signal_11704 ;
    wire signal_11706 ;
    wire signal_11708 ;
    wire signal_11710 ;
    wire signal_11712 ;
    wire signal_11714 ;
    wire signal_11716 ;
    wire signal_11718 ;
    wire signal_11720 ;
    wire signal_11722 ;
    wire signal_11724 ;
    wire signal_11726 ;
    wire signal_11728 ;
    wire signal_11730 ;
    wire signal_11732 ;
    wire signal_11734 ;
    wire signal_11736 ;
    wire signal_11738 ;
    wire signal_11740 ;
    wire signal_11742 ;
    wire signal_11744 ;
    wire signal_11746 ;
    wire signal_11748 ;
    wire signal_11750 ;
    wire signal_11752 ;
    wire signal_11754 ;
    wire signal_11756 ;
    wire signal_11758 ;
    wire signal_11760 ;
    wire signal_11762 ;
    wire signal_11764 ;
    wire signal_11766 ;
    wire signal_11768 ;
    wire signal_11770 ;
    wire signal_11772 ;
    wire signal_11774 ;
    wire signal_11776 ;
    wire signal_11778 ;
    wire signal_11780 ;
    wire signal_11782 ;
    wire signal_11784 ;
    wire signal_11786 ;
    wire signal_11788 ;
    wire signal_12469 ;

    /* cells in depth 0 */
    INV_X1 cell_0 ( .A (signal_395), .ZN (signal_400) ) ;
    INV_X1 cell_1 ( .A (signal_395), .ZN (signal_401) ) ;
    INV_X1 cell_2 ( .A (signal_395), .ZN (signal_398) ) ;
    INV_X1 cell_3 ( .A (signal_395), .ZN (signal_396) ) ;
    INV_X1 cell_4 ( .A (signal_395), .ZN (signal_397) ) ;
    INV_X1 cell_5 ( .A (signal_395), .ZN (signal_399) ) ;
    NOR2_X1 cell_6 ( .A1 (signal_406), .A2 (signal_411), .ZN (signal_395) ) ;
    INV_X1 cell_7 ( .A (signal_4388), .ZN (signal_406) ) ;
    INV_X1 cell_8 ( .A (signal_395), .ZN (signal_402) ) ;
    NOR2_X1 cell_9 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_404) ) ;
    INV_X1 cell_10 ( .A (signal_404), .ZN (signal_403) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_4388), .A2 (signal_403), .ZN (signal_4384) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_4388), .A2 (signal_4385), .ZN (signal_418) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_418), .A2 (signal_403), .ZN (signal_4383) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_4385), .A2 (signal_404), .ZN (signal_411) ) ;
    INV_X1 cell_15 ( .A (signal_4386), .ZN (signal_409) ) ;
    AND2_X1 cell_16 ( .A1 (signal_409), .A2 (signal_4387), .ZN (signal_414) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_418), .A2 (signal_414), .ZN (signal_405) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_402), .A2 (signal_405), .ZN (signal_4382) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_4385), .A2 (signal_406), .ZN (signal_416) ) ;
    NAND2_X1 cell_20 ( .A1 (signal_414), .A2 (signal_416), .ZN (signal_408) ) ;
    NAND2_X1 cell_21 ( .A1 (signal_4385), .A2 (signal_4384), .ZN (signal_407) ) ;
    NAND2_X1 cell_22 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_4381) ) ;
    NOR2_X1 cell_23 ( .A1 (signal_4387), .A2 (signal_409), .ZN (signal_412) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_418), .A2 (signal_412), .ZN (signal_410) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_411), .A2 (signal_410), .ZN (signal_4380) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_416), .A2 (signal_412), .ZN (signal_413) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_402), .A2 (signal_413), .ZN (signal_4379) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_179 ( .a ({signal_7457, signal_3750}), .b ({signal_7458, signal_4258}), .c ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_180 ( .a ({signal_7460, signal_3749}), .b ({signal_7461, signal_4257}), .c ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_181 ( .a ({signal_7463, signal_3748}), .b ({signal_7464, signal_4256}), .c ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_182 ( .a ({signal_7466, signal_3747}), .b ({signal_7467, signal_4255}), .c ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_183 ( .a ({signal_7469, signal_3746}), .b ({signal_7470, signal_4254}), .c ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_184 ( .a ({signal_7472, signal_3745}), .b ({signal_7473, signal_4253}), .c ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_185 ( .a ({signal_7475, signal_3744}), .b ({signal_7476, signal_4252}), .c ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_186 ( .a ({signal_7478, signal_3743}), .b ({signal_7479, signal_4251}), .c ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_235 ( .a ({signal_7481, signal_3814}), .b ({signal_7482, signal_4322}), .c ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_236 ( .a ({signal_7484, signal_3813}), .b ({signal_7485, signal_4321}), .c ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_237 ( .a ({signal_7487, signal_3812}), .b ({signal_7488, signal_4320}), .c ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_238 ( .a ({signal_7490, signal_3811}), .b ({signal_7491, signal_4319}), .c ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_240 ( .a ({signal_7493, signal_3810}), .b ({signal_7494, signal_4318}), .c ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_241 ( .a ({signal_7496, signal_3809}), .b ({signal_7497, signal_4317}), .c ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_242 ( .a ({signal_7499, signal_3808}), .b ({signal_7500, signal_4316}), .c ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_243 ( .a ({signal_7502, signal_3807}), .b ({signal_7503, signal_4315}), .c ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_270 ( .a ({signal_7505, signal_3782}), .b ({signal_7506, signal_4290}), .c ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_271 ( .a ({signal_7508, signal_3781}), .b ({signal_7509, signal_4289}), .c ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_273 ( .a ({signal_7511, signal_3780}), .b ({signal_7512, signal_4288}), .c ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_274 ( .a ({signal_7514, signal_3779}), .b ({signal_7515, signal_4287}), .c ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_275 ( .a ({signal_7517, signal_3778}), .b ({signal_7518, signal_4286}), .c ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_276 ( .a ({signal_7520, signal_3777}), .b ({signal_7521, signal_4285}), .c ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_277 ( .a ({signal_7523, signal_3776}), .b ({signal_7524, signal_4284}), .c ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_278 ( .a ({signal_7526, signal_3775}), .b ({signal_7527, signal_4283}), .c ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    NAND2_X1 cell_284 ( .A1 (signal_4385), .A2 (signal_414), .ZN (signal_415) ) ;
    NOR2_X1 cell_285 ( .A1 (signal_4388), .A2 (signal_415), .ZN (done) ) ;
    INV_X1 cell_286 ( .A (signal_416), .ZN (signal_417) ) ;
    NAND2_X1 cell_287 ( .A1 (signal_4386), .A2 (signal_4387), .ZN (signal_419) ) ;
    NOR2_X1 cell_288 ( .A1 (signal_417), .A2 (signal_419), .ZN (signal_393) ) ;
    INV_X1 cell_289 ( .A (signal_418), .ZN (signal_420) ) ;
    NOR2_X1 cell_290 ( .A1 (signal_420), .A2 (signal_419), .ZN (signal_394) ) ;
    INV_X1 cell_4187 ( .A (signal_3597), .ZN (signal_3607) ) ;
    MUX2_X1 cell_4188 ( .S (signal_3609), .A (signal_3598), .B (signal_3599), .Z (signal_3597) ) ;
    NOR2_X1 cell_4189 ( .A1 (reset), .A2 (signal_3600), .ZN (signal_3610) ) ;
    XNOR2_X1 cell_4190 ( .A (signal_4388), .B (signal_4387), .ZN (signal_3600) ) ;
    MUX2_X1 cell_4191 ( .S (signal_4385), .A (signal_3601), .B (signal_3602), .Z (signal_3608) ) ;
    NAND2_X1 cell_4192 ( .A1 (signal_3598), .A2 (signal_3603), .ZN (signal_3602) ) ;
    NAND2_X1 cell_4193 ( .A1 (signal_3609), .A2 (signal_3606), .ZN (signal_3603) ) ;
    NOR2_X1 cell_4194 ( .A1 (signal_3604), .A2 (signal_3612), .ZN (signal_3598) ) ;
    NOR2_X1 cell_4195 ( .A1 (signal_4387), .A2 (reset), .ZN (signal_3604) ) ;
    NOR2_X1 cell_4196 ( .A1 (signal_3609), .A2 (signal_3599), .ZN (signal_3601) ) ;
    NAND2_X1 cell_4197 ( .A1 (signal_4387), .A2 (signal_3605), .ZN (signal_3599) ) ;
    NOR2_X1 cell_4198 ( .A1 (reset), .A2 (signal_3611), .ZN (signal_3605) ) ;
    NOR2_X1 cell_4199 ( .A1 (reset), .A2 (signal_4388), .ZN (signal_3612) ) ;
    INV_X1 cell_4200 ( .A (reset), .ZN (signal_3606) ) ;
    INV_X1 cell_4201 ( .A (signal_4388), .ZN (signal_3611) ) ;
    INV_X1 cell_4205 ( .A (signal_4386), .ZN (signal_3609) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4209 ( .a ({signal_7529, signal_4378}), .b ({signal_7530, signal_3870}), .c ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4210 ( .a ({signal_7532, signal_4278}), .b ({signal_7533, signal_3770}), .c ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4211 ( .a ({signal_7535, signal_4277}), .b ({signal_7536, signal_3769}), .c ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4212 ( .a ({signal_7538, signal_4276}), .b ({signal_7539, signal_3768}), .c ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4213 ( .a ({signal_7541, signal_4275}), .b ({signal_7542, signal_3767}), .c ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4214 ( .a ({signal_7544, signal_4274}), .b ({signal_7545, signal_3766}), .c ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4215 ( .a ({signal_7547, signal_4273}), .b ({signal_7548, signal_3765}), .c ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4216 ( .a ({signal_7550, signal_4272}), .b ({signal_7551, signal_3764}), .c ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4217 ( .a ({signal_7553, signal_4271}), .b ({signal_7554, signal_3763}), .c ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4218 ( .a ({signal_7556, signal_4270}), .b ({signal_7557, signal_3762}), .c ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4219 ( .a ({signal_7559, signal_4269}), .b ({signal_7560, signal_3761}), .c ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4220 ( .a ({signal_7562, signal_4368}), .b ({signal_7563, signal_3860}), .c ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4221 ( .a ({signal_7565, signal_4268}), .b ({signal_7566, signal_3760}), .c ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4222 ( .a ({signal_7568, signal_4267}), .b ({signal_7569, signal_3759}), .c ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4223 ( .a ({signal_7571, signal_4266}), .b ({signal_7572, signal_3758}), .c ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4224 ( .a ({signal_7574, signal_4265}), .b ({signal_7575, signal_3757}), .c ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4225 ( .a ({signal_7577, signal_4264}), .b ({signal_7578, signal_3756}), .c ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4226 ( .a ({signal_7580, signal_4263}), .b ({signal_7581, signal_3755}), .c ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4227 ( .a ({signal_7583, signal_4262}), .b ({signal_7584, signal_3754}), .c ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4228 ( .a ({signal_7586, signal_4261}), .b ({signal_7587, signal_3753}), .c ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4229 ( .a ({signal_7589, signal_4260}), .b ({signal_7590, signal_3752}), .c ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4230 ( .a ({signal_7592, signal_4259}), .b ({signal_7593, signal_3751}), .c ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4231 ( .a ({signal_7595, signal_4367}), .b ({signal_7596, signal_3859}), .c ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4232 ( .a ({signal_7598, signal_4366}), .b ({signal_7599, signal_3858}), .c ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4233 ( .a ({signal_7601, signal_4365}), .b ({signal_7602, signal_3857}), .c ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4234 ( .a ({signal_7604, signal_4364}), .b ({signal_7605, signal_3856}), .c ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4235 ( .a ({signal_7607, signal_4363}), .b ({signal_7608, signal_3855}), .c ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4236 ( .a ({signal_7610, signal_4362}), .b ({signal_7611, signal_3854}), .c ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4237 ( .a ({signal_7613, signal_4361}), .b ({signal_7614, signal_3853}), .c ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4238 ( .a ({signal_7616, signal_4360}), .b ({signal_7617, signal_3852}), .c ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4239 ( .a ({signal_7619, signal_4359}), .b ({signal_7620, signal_3851}), .c ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4240 ( .a ({signal_7622, signal_4377}), .b ({signal_7623, signal_3869}), .c ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4241 ( .a ({signal_7625, signal_4358}), .b ({signal_7626, signal_3850}), .c ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4242 ( .a ({signal_7628, signal_4357}), .b ({signal_7629, signal_3849}), .c ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4243 ( .a ({signal_7631, signal_4356}), .b ({signal_7632, signal_3848}), .c ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4244 ( .a ({signal_7634, signal_4355}), .b ({signal_7635, signal_3847}), .c ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4245 ( .a ({signal_7637, signal_4354}), .b ({signal_7638, signal_3846}), .c ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4246 ( .a ({signal_7640, signal_4353}), .b ({signal_7641, signal_3845}), .c ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4247 ( .a ({signal_7643, signal_4352}), .b ({signal_7644, signal_3844}), .c ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4248 ( .a ({signal_7646, signal_4351}), .b ({signal_7647, signal_3843}), .c ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4249 ( .a ({signal_7649, signal_4350}), .b ({signal_7650, signal_3842}), .c ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4250 ( .a ({signal_7652, signal_4349}), .b ({signal_7653, signal_3841}), .c ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4251 ( .a ({signal_7655, signal_4376}), .b ({signal_7656, signal_3868}), .c ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4252 ( .a ({signal_7658, signal_4348}), .b ({signal_7659, signal_3840}), .c ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4253 ( .a ({signal_7661, signal_4347}), .b ({signal_7662, signal_3839}), .c ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4254 ( .a ({signal_7664, signal_4346}), .b ({signal_7665, signal_3838}), .c ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4255 ( .a ({signal_7667, signal_4345}), .b ({signal_7668, signal_3837}), .c ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4256 ( .a ({signal_7670, signal_4344}), .b ({signal_7671, signal_3836}), .c ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4257 ( .a ({signal_7673, signal_4343}), .b ({signal_7674, signal_3835}), .c ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4258 ( .a ({signal_7676, signal_4342}), .b ({signal_7677, signal_3834}), .c ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4259 ( .a ({signal_7679, signal_4341}), .b ({signal_7680, signal_3833}), .c ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4260 ( .a ({signal_7682, signal_4340}), .b ({signal_7683, signal_3832}), .c ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4261 ( .a ({signal_7685, signal_4339}), .b ({signal_7686, signal_3831}), .c ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4262 ( .a ({signal_7688, signal_4375}), .b ({signal_7689, signal_3867}), .c ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4263 ( .a ({signal_7691, signal_4338}), .b ({signal_7692, signal_3830}), .c ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4264 ( .a ({signal_7694, signal_4337}), .b ({signal_7695, signal_3829}), .c ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4265 ( .a ({signal_7697, signal_4336}), .b ({signal_7698, signal_3828}), .c ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4266 ( .a ({signal_7700, signal_4335}), .b ({signal_7701, signal_3827}), .c ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4267 ( .a ({signal_7703, signal_4334}), .b ({signal_7704, signal_3826}), .c ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4268 ( .a ({signal_7706, signal_4333}), .b ({signal_7707, signal_3825}), .c ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4269 ( .a ({signal_7709, signal_4332}), .b ({signal_7710, signal_3824}), .c ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4270 ( .a ({signal_7712, signal_4331}), .b ({signal_7713, signal_3823}), .c ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4271 ( .a ({signal_7715, signal_4330}), .b ({signal_7716, signal_3822}), .c ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4272 ( .a ({signal_7718, signal_4329}), .b ({signal_7719, signal_3821}), .c ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4273 ( .a ({signal_7721, signal_4374}), .b ({signal_7722, signal_3866}), .c ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4274 ( .a ({signal_7724, signal_4328}), .b ({signal_7725, signal_3820}), .c ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4275 ( .a ({signal_7727, signal_4327}), .b ({signal_7728, signal_3819}), .c ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4276 ( .a ({signal_7730, signal_4326}), .b ({signal_7731, signal_3818}), .c ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4277 ( .a ({signal_7733, signal_4325}), .b ({signal_7734, signal_3817}), .c ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4278 ( .a ({signal_7736, signal_4324}), .b ({signal_7737, signal_3816}), .c ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4279 ( .a ({signal_7739, signal_4323}), .b ({signal_7740, signal_3815}), .c ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4280 ( .a ({signal_7742, signal_4373}), .b ({signal_7743, signal_3865}), .c ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4281 ( .a ({signal_7745, signal_4314}), .b ({signal_7746, signal_3806}), .c ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4282 ( .a ({signal_7748, signal_4313}), .b ({signal_7749, signal_3805}), .c ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4283 ( .a ({signal_7751, signal_4312}), .b ({signal_7752, signal_3804}), .c ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4284 ( .a ({signal_7754, signal_4311}), .b ({signal_7755, signal_3803}), .c ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4285 ( .a ({signal_7757, signal_4310}), .b ({signal_7758, signal_3802}), .c ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4286 ( .a ({signal_7760, signal_4309}), .b ({signal_7761, signal_3801}), .c ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4287 ( .a ({signal_7763, signal_4372}), .b ({signal_7764, signal_3864}), .c ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4288 ( .a ({signal_7766, signal_4308}), .b ({signal_7767, signal_3800}), .c ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4289 ( .a ({signal_7769, signal_4307}), .b ({signal_7770, signal_3799}), .c ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4290 ( .a ({signal_7772, signal_4306}), .b ({signal_7773, signal_3798}), .c ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4291 ( .a ({signal_7775, signal_4305}), .b ({signal_7776, signal_3797}), .c ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4292 ( .a ({signal_7778, signal_4304}), .b ({signal_7779, signal_3796}), .c ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4293 ( .a ({signal_7781, signal_4303}), .b ({signal_7782, signal_3795}), .c ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4294 ( .a ({signal_7784, signal_4302}), .b ({signal_7785, signal_3794}), .c ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4295 ( .a ({signal_7787, signal_4301}), .b ({signal_7788, signal_3793}), .c ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4296 ( .a ({signal_7790, signal_4300}), .b ({signal_7791, signal_3792}), .c ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4297 ( .a ({signal_7793, signal_4299}), .b ({signal_7794, signal_3791}), .c ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4298 ( .a ({signal_7796, signal_4371}), .b ({signal_7797, signal_3863}), .c ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4299 ( .a ({signal_7799, signal_4298}), .b ({signal_7800, signal_3790}), .c ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4300 ( .a ({signal_7802, signal_4297}), .b ({signal_7803, signal_3789}), .c ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4301 ( .a ({signal_7805, signal_4296}), .b ({signal_7806, signal_3788}), .c ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4302 ( .a ({signal_7808, signal_4295}), .b ({signal_7809, signal_3787}), .c ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4303 ( .a ({signal_7811, signal_4294}), .b ({signal_7812, signal_3786}), .c ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4304 ( .a ({signal_7814, signal_4293}), .b ({signal_7815, signal_3785}), .c ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4305 ( .a ({signal_7817, signal_4292}), .b ({signal_7818, signal_3784}), .c ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4306 ( .a ({signal_7820, signal_4291}), .b ({signal_7821, signal_3783}), .c ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4307 ( .a ({signal_7823, signal_4370}), .b ({signal_7824, signal_3862}), .c ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4308 ( .a ({signal_7826, signal_4282}), .b ({signal_7827, signal_3774}), .c ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4309 ( .a ({signal_7829, signal_4281}), .b ({signal_7830, signal_3773}), .c ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4310 ( .a ({signal_7832, signal_4280}), .b ({signal_7833, signal_3772}), .c ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4311 ( .a ({signal_7835, signal_4279}), .b ({signal_7836, signal_3771}), .c ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4312 ( .a ({signal_7838, signal_4369}), .b ({signal_7839, signal_3861}), .c ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4313 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_7881, signal_4549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4314 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_7882, signal_4550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4315 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .c ({signal_7883, signal_4551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4316 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_7884, signal_4552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4317 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .c ({signal_7885, signal_4553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4318 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_7886, signal_4554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4319 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .c ({signal_7887, signal_4555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4320 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .c ({signal_7888, signal_4556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4321 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .c ({signal_7889, signal_4557}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4322 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .c ({signal_7890, signal_4558}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4323 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_7891, signal_4559}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4324 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_7892, signal_4560}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4325 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .c ({signal_7893, signal_4561}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4326 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_7894, signal_4562}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4327 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .c ({signal_7895, signal_4563}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4328 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_7896, signal_4564}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4329 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .c ({signal_7897, signal_4565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4330 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .c ({signal_7898, signal_4566}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4331 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .c ({signal_7899, signal_4567}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4332 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .c ({signal_7900, signal_4568}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4333 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_7901, signal_4569}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4334 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_7902, signal_4570}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4335 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .c ({signal_7903, signal_4571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4336 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_7904, signal_4572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4337 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .c ({signal_7905, signal_4573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4338 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_7906, signal_4574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4339 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .c ({signal_7907, signal_4575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4340 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .c ({signal_7908, signal_4576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4341 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .c ({signal_7909, signal_4577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4342 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .c ({signal_7910, signal_4578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4343 ( .a ({signal_7634, signal_4355}), .b ({signal_7625, signal_4358}), .c ({signal_7841, signal_4579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4344 ( .a ({signal_7634, signal_4355}), .b ({signal_7616, signal_4360}), .c ({signal_7842, signal_4580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4345 ( .a ({signal_7634, signal_4355}), .b ({signal_7613, signal_4361}), .c ({signal_7843, signal_4581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4346 ( .a ({signal_7625, signal_4358}), .b ({signal_7616, signal_4360}), .c ({signal_7844, signal_4582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4347 ( .a ({signal_7619, signal_4359}), .b ({signal_7613, signal_4361}), .c ({signal_7845, signal_4583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4348 ( .a ({signal_7631, signal_4356}), .b ({signal_7628, signal_4357}), .c ({signal_7846, signal_4584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4349 ( .a ({signal_7631, signal_4356}), .b ({signal_7616, signal_4360}), .c ({signal_7847, signal_4585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4350 ( .a ({signal_7628, signal_4357}), .b ({signal_7616, signal_4360}), .c ({signal_7848, signal_4586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4351 ( .a ({signal_7625, signal_4358}), .b ({signal_7610, signal_4362}), .c ({signal_7849, signal_4587}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4352 ( .a ({signal_7613, signal_4361}), .b ({signal_7610, signal_4362}), .c ({signal_7850, signal_4588}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4353 ( .a ({signal_7607, signal_4363}), .b ({signal_7598, signal_4366}), .c ({signal_7851, signal_4589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4354 ( .a ({signal_7607, signal_4363}), .b ({signal_7562, signal_4368}), .c ({signal_7852, signal_4590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4355 ( .a ({signal_7607, signal_4363}), .b ({signal_7838, signal_4369}), .c ({signal_7853, signal_4591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4356 ( .a ({signal_7598, signal_4366}), .b ({signal_7562, signal_4368}), .c ({signal_7854, signal_4592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4357 ( .a ({signal_7595, signal_4367}), .b ({signal_7838, signal_4369}), .c ({signal_7855, signal_4593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4358 ( .a ({signal_7604, signal_4364}), .b ({signal_7601, signal_4365}), .c ({signal_7856, signal_4594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4359 ( .a ({signal_7604, signal_4364}), .b ({signal_7562, signal_4368}), .c ({signal_7857, signal_4595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4360 ( .a ({signal_7601, signal_4365}), .b ({signal_7562, signal_4368}), .c ({signal_7858, signal_4596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4361 ( .a ({signal_7598, signal_4366}), .b ({signal_7823, signal_4370}), .c ({signal_7859, signal_4597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4362 ( .a ({signal_7838, signal_4369}), .b ({signal_7823, signal_4370}), .c ({signal_7860, signal_4598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4363 ( .a ({signal_7796, signal_4371}), .b ({signal_7721, signal_4374}), .c ({signal_7861, signal_4599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4364 ( .a ({signal_7796, signal_4371}), .b ({signal_7655, signal_4376}), .c ({signal_7862, signal_4600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4365 ( .a ({signal_7796, signal_4371}), .b ({signal_7622, signal_4377}), .c ({signal_7863, signal_4601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4366 ( .a ({signal_7721, signal_4374}), .b ({signal_7655, signal_4376}), .c ({signal_7864, signal_4602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4367 ( .a ({signal_7688, signal_4375}), .b ({signal_7622, signal_4377}), .c ({signal_7865, signal_4603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4368 ( .a ({signal_7763, signal_4372}), .b ({signal_7742, signal_4373}), .c ({signal_7866, signal_4604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4369 ( .a ({signal_7763, signal_4372}), .b ({signal_7655, signal_4376}), .c ({signal_7867, signal_4605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4370 ( .a ({signal_7742, signal_4373}), .b ({signal_7655, signal_4376}), .c ({signal_7868, signal_4606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4371 ( .a ({signal_7721, signal_4374}), .b ({signal_7529, signal_4378}), .c ({signal_7869, signal_4607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4372 ( .a ({signal_7622, signal_4377}), .b ({signal_7529, signal_4378}), .c ({signal_7870, signal_4608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4373 ( .a ({signal_7661, signal_4347}), .b ({signal_7649, signal_4350}), .c ({signal_7871, signal_4609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4374 ( .a ({signal_7661, signal_4347}), .b ({signal_7643, signal_4352}), .c ({signal_7872, signal_4610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4375 ( .a ({signal_7661, signal_4347}), .b ({signal_7640, signal_4353}), .c ({signal_7873, signal_4611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4376 ( .a ({signal_7649, signal_4350}), .b ({signal_7643, signal_4352}), .c ({signal_7874, signal_4612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4377 ( .a ({signal_7646, signal_4351}), .b ({signal_7640, signal_4353}), .c ({signal_7875, signal_4613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4378 ( .a ({signal_7658, signal_4348}), .b ({signal_7652, signal_4349}), .c ({signal_7876, signal_4614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4379 ( .a ({signal_7658, signal_4348}), .b ({signal_7643, signal_4352}), .c ({signal_7877, signal_4615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4380 ( .a ({signal_7652, signal_4349}), .b ({signal_7643, signal_4352}), .c ({signal_7878, signal_4616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4381 ( .a ({signal_7649, signal_4350}), .b ({signal_7637, signal_4354}), .c ({signal_7879, signal_4617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4382 ( .a ({signal_7640, signal_4353}), .b ({signal_7637, signal_4354}), .c ({signal_7880, signal_4618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4383 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_7911, signal_4619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4384 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_7912, signal_4620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4385 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .c ({signal_7913, signal_4621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4386 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_7914, signal_4622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4387 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .c ({signal_7915, signal_4623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4388 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_7916, signal_4624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4389 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .c ({signal_7917, signal_4625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4390 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .c ({signal_7918, signal_4626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4391 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .c ({signal_7919, signal_4627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4392 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .c ({signal_7920, signal_4628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4393 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_7921, signal_4629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4394 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .c ({signal_7922, signal_4630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4395 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_7923, signal_4631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4396 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .c ({signal_7924, signal_4632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4397 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_7925, signal_4633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4398 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_7926, signal_4634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4399 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .c ({signal_7927, signal_4635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4400 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .c ({signal_7928, signal_4636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4401 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .c ({signal_7929, signal_4637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4402 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .c ({signal_7930, signal_4638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4403 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_7931, signal_4639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4404 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_7932, signal_4640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4405 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .c ({signal_7933, signal_4641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4406 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_7934, signal_4642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4407 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .c ({signal_7935, signal_4643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4408 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_7936, signal_4644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4409 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .c ({signal_7937, signal_4645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4410 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .c ({signal_7938, signal_4646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4411 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .c ({signal_7939, signal_4647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4412 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .c ({signal_7940, signal_4648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4413 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_7941, signal_4649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4414 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_7942, signal_4650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4415 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .c ({signal_7943, signal_4651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4416 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_7944, signal_4652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4417 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .c ({signal_7945, signal_4653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4418 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_7946, signal_4654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4419 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .c ({signal_7947, signal_4655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4420 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .c ({signal_7948, signal_4656}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4421 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .c ({signal_7949, signal_4657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4422 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .c ({signal_7950, signal_4658}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4423 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_7951, signal_4659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4424 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_7952, signal_4660}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4425 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .c ({signal_7953, signal_4661}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4426 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_7954, signal_4662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4427 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .c ({signal_7955, signal_4663}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4428 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_7956, signal_4664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4429 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .c ({signal_7957, signal_4665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4430 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .c ({signal_7958, signal_4666}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4431 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .c ({signal_7959, signal_4667}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4432 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .c ({signal_7960, signal_4668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4433 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_7961, signal_4669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4434 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_7962, signal_4670}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4435 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .c ({signal_7963, signal_4671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4436 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_7964, signal_4672}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4437 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .c ({signal_7965, signal_4673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4438 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_7966, signal_4674}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4439 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .c ({signal_7967, signal_4675}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4440 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .c ({signal_7968, signal_4676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4441 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .c ({signal_7969, signal_4677}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4442 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .c ({signal_7970, signal_4678}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4443 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_7971, signal_4679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4444 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_7972, signal_4680}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4445 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .c ({signal_7973, signal_4681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4446 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_7974, signal_4682}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4447 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .c ({signal_7975, signal_4683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4448 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_7976, signal_4684}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4449 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .c ({signal_7977, signal_4685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4450 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .c ({signal_7978, signal_4686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4451 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .c ({signal_7979, signal_4687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4452 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .c ({signal_7980, signal_4688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4453 ( .a ({signal_7881, signal_4549}), .b ({signal_7885, signal_4553}), .c ({signal_8073, signal_4689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4454 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_7886, signal_4554}), .c ({signal_8074, signal_4690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4455 ( .a ({signal_7883, signal_4551}), .b ({signal_7884, signal_4552}), .c ({signal_8075, signal_4691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4456 ( .a ({signal_7885, signal_4553}), .b ({signal_7887, signal_4555}), .c ({signal_8076, signal_4692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4457 ( .a ({signal_7885, signal_4553}), .b ({signal_7888, signal_4556}), .c ({signal_8077, signal_4693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4458 ( .a ({signal_7886, signal_4554}), .b ({signal_7889, signal_4557}), .c ({signal_8078, signal_4694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4459 ( .a ({signal_7886, signal_4554}), .b ({signal_7890, signal_4558}), .c ({signal_8079, signal_4695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4460 ( .a ({signal_7881, signal_4549}), .b ({signal_7888, signal_4556}), .c ({signal_8080, signal_4696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4461 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_7981, signal_4697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4462 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_7982, signal_4698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4463 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .c ({signal_7983, signal_4699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4464 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_7984, signal_4700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4465 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .c ({signal_7985, signal_4701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4466 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_7986, signal_4702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4467 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .c ({signal_7987, signal_4703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4468 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .c ({signal_7988, signal_4704}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4469 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .c ({signal_7989, signal_4705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4470 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .c ({signal_7990, signal_4706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4471 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_7991, signal_4707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4472 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_7992, signal_4708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4473 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .c ({signal_7993, signal_4709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4474 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_7994, signal_4710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4475 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .c ({signal_7995, signal_4711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4476 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_7996, signal_4712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4477 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .c ({signal_7997, signal_4713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4478 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .c ({signal_7998, signal_4714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4479 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .c ({signal_7999, signal_4715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4480 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .c ({signal_8000, signal_4716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4481 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_8001, signal_4717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4482 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_8002, signal_4718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4483 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .c ({signal_8003, signal_4719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4484 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_8004, signal_4720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4485 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .c ({signal_8005, signal_4721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4486 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_8006, signal_4722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4487 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .c ({signal_8007, signal_4723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4488 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .c ({signal_8008, signal_4724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4489 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .c ({signal_8009, signal_4725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4490 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .c ({signal_8010, signal_4726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4491 ( .a ({signal_7891, signal_4559}), .b ({signal_7895, signal_4563}), .c ({signal_8081, signal_4727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4492 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_7896, signal_4564}), .c ({signal_8082, signal_4728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4493 ( .a ({signal_7893, signal_4561}), .b ({signal_7894, signal_4562}), .c ({signal_8083, signal_4729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4494 ( .a ({signal_7895, signal_4563}), .b ({signal_7897, signal_4565}), .c ({signal_8084, signal_4730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4495 ( .a ({signal_7895, signal_4563}), .b ({signal_7898, signal_4566}), .c ({signal_8085, signal_4731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4496 ( .a ({signal_7896, signal_4564}), .b ({signal_7899, signal_4567}), .c ({signal_8086, signal_4732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4497 ( .a ({signal_7896, signal_4564}), .b ({signal_7900, signal_4568}), .c ({signal_8087, signal_4733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4498 ( .a ({signal_7891, signal_4559}), .b ({signal_7898, signal_4566}), .c ({signal_8088, signal_4734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4499 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .c ({signal_8011, signal_4735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4500 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8012, signal_4736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4501 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_8013, signal_4737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4502 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8014, signal_4738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4503 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .c ({signal_8015, signal_4739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4504 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .c ({signal_8016, signal_4740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4505 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8017, signal_4741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4506 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .c ({signal_8018, signal_4742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4507 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .c ({signal_8019, signal_4743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4508 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .c ({signal_8020, signal_4744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4509 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_8021, signal_4745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4510 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_8022, signal_4746}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4511 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .c ({signal_8023, signal_4747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4512 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_8024, signal_4748}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4513 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .c ({signal_8025, signal_4749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4514 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_8026, signal_4750}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4515 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .c ({signal_8027, signal_4751}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4516 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .c ({signal_8028, signal_4752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4517 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .c ({signal_8029, signal_4753}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4518 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .c ({signal_8030, signal_4754}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4519 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_8031, signal_4755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4520 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_8032, signal_4756}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4521 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .c ({signal_8033, signal_4757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4522 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_8034, signal_4758}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4523 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .c ({signal_8035, signal_4759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4524 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_8036, signal_4760}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4525 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .c ({signal_8037, signal_4761}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4526 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .c ({signal_8038, signal_4762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4527 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .c ({signal_8039, signal_4763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4528 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .c ({signal_8040, signal_4764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4529 ( .a ({signal_7901, signal_4569}), .b ({signal_7905, signal_4573}), .c ({signal_8089, signal_4765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4530 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_7906, signal_4574}), .c ({signal_8090, signal_4766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4531 ( .a ({signal_7903, signal_4571}), .b ({signal_7904, signal_4572}), .c ({signal_8091, signal_4767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4532 ( .a ({signal_7905, signal_4573}), .b ({signal_7907, signal_4575}), .c ({signal_8092, signal_4768}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4533 ( .a ({signal_7905, signal_4573}), .b ({signal_7908, signal_4576}), .c ({signal_8093, signal_4769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4534 ( .a ({signal_7906, signal_4574}), .b ({signal_7909, signal_4577}), .c ({signal_8094, signal_4770}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4535 ( .a ({signal_7906, signal_4574}), .b ({signal_7910, signal_4578}), .c ({signal_8095, signal_4771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4536 ( .a ({signal_7901, signal_4569}), .b ({signal_7908, signal_4576}), .c ({signal_8096, signal_4772}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4537 ( .a ({signal_7841, signal_4579}), .b ({signal_7845, signal_4583}), .c ({signal_8041, signal_4773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4538 ( .a ({signal_7610, signal_4362}), .b ({signal_7846, signal_4584}), .c ({signal_8042, signal_4774}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4539 ( .a ({signal_7843, signal_4581}), .b ({signal_7844, signal_4582}), .c ({signal_8043, signal_4775}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4540 ( .a ({signal_7845, signal_4583}), .b ({signal_7847, signal_4585}), .c ({signal_8044, signal_4776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4541 ( .a ({signal_7845, signal_4583}), .b ({signal_7848, signal_4586}), .c ({signal_8045, signal_4777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4542 ( .a ({signal_7846, signal_4584}), .b ({signal_7849, signal_4587}), .c ({signal_8046, signal_4778}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4543 ( .a ({signal_7846, signal_4584}), .b ({signal_7850, signal_4588}), .c ({signal_8047, signal_4779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4544 ( .a ({signal_7841, signal_4579}), .b ({signal_7848, signal_4586}), .c ({signal_8048, signal_4780}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4545 ( .a ({signal_7851, signal_4589}), .b ({signal_7855, signal_4593}), .c ({signal_8049, signal_4781}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4546 ( .a ({signal_7823, signal_4370}), .b ({signal_7856, signal_4594}), .c ({signal_8050, signal_4782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4547 ( .a ({signal_7853, signal_4591}), .b ({signal_7854, signal_4592}), .c ({signal_8051, signal_4783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4548 ( .a ({signal_7855, signal_4593}), .b ({signal_7857, signal_4595}), .c ({signal_8052, signal_4784}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4549 ( .a ({signal_7855, signal_4593}), .b ({signal_7858, signal_4596}), .c ({signal_8053, signal_4785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4550 ( .a ({signal_7856, signal_4594}), .b ({signal_7859, signal_4597}), .c ({signal_8054, signal_4786}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4551 ( .a ({signal_7856, signal_4594}), .b ({signal_7860, signal_4598}), .c ({signal_8055, signal_4787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4552 ( .a ({signal_7851, signal_4589}), .b ({signal_7858, signal_4596}), .c ({signal_8056, signal_4788}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4553 ( .a ({signal_7861, signal_4599}), .b ({signal_7865, signal_4603}), .c ({signal_8057, signal_4789}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4554 ( .a ({signal_7529, signal_4378}), .b ({signal_7866, signal_4604}), .c ({signal_8058, signal_4790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4555 ( .a ({signal_7863, signal_4601}), .b ({signal_7864, signal_4602}), .c ({signal_8059, signal_4791}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4556 ( .a ({signal_7865, signal_4603}), .b ({signal_7867, signal_4605}), .c ({signal_8060, signal_4792}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4557 ( .a ({signal_7865, signal_4603}), .b ({signal_7868, signal_4606}), .c ({signal_8061, signal_4793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4558 ( .a ({signal_7866, signal_4604}), .b ({signal_7869, signal_4607}), .c ({signal_8062, signal_4794}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4559 ( .a ({signal_7866, signal_4604}), .b ({signal_7870, signal_4608}), .c ({signal_8063, signal_4795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4560 ( .a ({signal_7861, signal_4599}), .b ({signal_7868, signal_4606}), .c ({signal_8064, signal_4796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4561 ( .a ({signal_7871, signal_4609}), .b ({signal_7875, signal_4613}), .c ({signal_8065, signal_4797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4562 ( .a ({signal_7637, signal_4354}), .b ({signal_7876, signal_4614}), .c ({signal_8066, signal_4798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4563 ( .a ({signal_7873, signal_4611}), .b ({signal_7874, signal_4612}), .c ({signal_8067, signal_4799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4564 ( .a ({signal_7875, signal_4613}), .b ({signal_7877, signal_4615}), .c ({signal_8068, signal_4800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4565 ( .a ({signal_7875, signal_4613}), .b ({signal_7878, signal_4616}), .c ({signal_8069, signal_4801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4566 ( .a ({signal_7876, signal_4614}), .b ({signal_7879, signal_4617}), .c ({signal_8070, signal_4802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4567 ( .a ({signal_7876, signal_4614}), .b ({signal_7880, signal_4618}), .c ({signal_8071, signal_4803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4568 ( .a ({signal_7871, signal_4609}), .b ({signal_7878, signal_4616}), .c ({signal_8072, signal_4804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4611 ( .a ({signal_7911, signal_4619}), .b ({signal_7915, signal_4623}), .c ({signal_8121, signal_4847}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4612 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_7916, signal_4624}), .c ({signal_8122, signal_4848}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4613 ( .a ({signal_7913, signal_4621}), .b ({signal_7914, signal_4622}), .c ({signal_8123, signal_4849}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4614 ( .a ({signal_7915, signal_4623}), .b ({signal_7917, signal_4625}), .c ({signal_8124, signal_4850}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4615 ( .a ({signal_7915, signal_4623}), .b ({signal_7918, signal_4626}), .c ({signal_8125, signal_4851}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4616 ( .a ({signal_7916, signal_4624}), .b ({signal_7919, signal_4627}), .c ({signal_8126, signal_4852}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4617 ( .a ({signal_7916, signal_4624}), .b ({signal_7920, signal_4628}), .c ({signal_8127, signal_4853}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4618 ( .a ({signal_7911, signal_4619}), .b ({signal_7918, signal_4626}), .c ({signal_8128, signal_4854}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4619 ( .a ({signal_7921, signal_4629}), .b ({signal_7925, signal_4633}), .c ({signal_8129, signal_4855}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4620 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_7926, signal_4634}), .c ({signal_8130, signal_4856}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4621 ( .a ({signal_7923, signal_4631}), .b ({signal_7924, signal_4632}), .c ({signal_8131, signal_4857}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4622 ( .a ({signal_7925, signal_4633}), .b ({signal_7927, signal_4635}), .c ({signal_8132, signal_4858}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4623 ( .a ({signal_7925, signal_4633}), .b ({signal_7928, signal_4636}), .c ({signal_8133, signal_4859}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4624 ( .a ({signal_7926, signal_4634}), .b ({signal_7929, signal_4637}), .c ({signal_8134, signal_4860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4625 ( .a ({signal_7926, signal_4634}), .b ({signal_7930, signal_4638}), .c ({signal_8135, signal_4861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4626 ( .a ({signal_7921, signal_4629}), .b ({signal_7928, signal_4636}), .c ({signal_8136, signal_4862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4627 ( .a ({signal_7931, signal_4639}), .b ({signal_7935, signal_4643}), .c ({signal_8137, signal_4863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4628 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_7936, signal_4644}), .c ({signal_8138, signal_4864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4629 ( .a ({signal_7933, signal_4641}), .b ({signal_7934, signal_4642}), .c ({signal_8139, signal_4865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4630 ( .a ({signal_7935, signal_4643}), .b ({signal_7937, signal_4645}), .c ({signal_8140, signal_4866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4631 ( .a ({signal_7935, signal_4643}), .b ({signal_7938, signal_4646}), .c ({signal_8141, signal_4867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4632 ( .a ({signal_7936, signal_4644}), .b ({signal_7939, signal_4647}), .c ({signal_8142, signal_4868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4633 ( .a ({signal_7936, signal_4644}), .b ({signal_7940, signal_4648}), .c ({signal_8143, signal_4869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4634 ( .a ({signal_7931, signal_4639}), .b ({signal_7938, signal_4646}), .c ({signal_8144, signal_4870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4635 ( .a ({signal_7941, signal_4649}), .b ({signal_7945, signal_4653}), .c ({signal_8145, signal_4871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4636 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_7946, signal_4654}), .c ({signal_8146, signal_4872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4637 ( .a ({signal_7943, signal_4651}), .b ({signal_7944, signal_4652}), .c ({signal_8147, signal_4873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4638 ( .a ({signal_7945, signal_4653}), .b ({signal_7947, signal_4655}), .c ({signal_8148, signal_4874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4639 ( .a ({signal_7945, signal_4653}), .b ({signal_7948, signal_4656}), .c ({signal_8149, signal_4875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4640 ( .a ({signal_7946, signal_4654}), .b ({signal_7949, signal_4657}), .c ({signal_8150, signal_4876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4641 ( .a ({signal_7946, signal_4654}), .b ({signal_7950, signal_4658}), .c ({signal_8151, signal_4877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4642 ( .a ({signal_7941, signal_4649}), .b ({signal_7948, signal_4656}), .c ({signal_8152, signal_4878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4643 ( .a ({signal_7951, signal_4659}), .b ({signal_7955, signal_4663}), .c ({signal_8153, signal_4879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4644 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_7956, signal_4664}), .c ({signal_8154, signal_4880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4645 ( .a ({signal_7953, signal_4661}), .b ({signal_7954, signal_4662}), .c ({signal_8155, signal_4881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4646 ( .a ({signal_7955, signal_4663}), .b ({signal_7957, signal_4665}), .c ({signal_8156, signal_4882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4647 ( .a ({signal_7955, signal_4663}), .b ({signal_7958, signal_4666}), .c ({signal_8157, signal_4883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4648 ( .a ({signal_7956, signal_4664}), .b ({signal_7959, signal_4667}), .c ({signal_8158, signal_4884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4649 ( .a ({signal_7956, signal_4664}), .b ({signal_7960, signal_4668}), .c ({signal_8159, signal_4885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4650 ( .a ({signal_7951, signal_4659}), .b ({signal_7958, signal_4666}), .c ({signal_8160, signal_4886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4651 ( .a ({signal_7961, signal_4669}), .b ({signal_7965, signal_4673}), .c ({signal_8161, signal_4887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4652 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_7966, signal_4674}), .c ({signal_8162, signal_4888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4653 ( .a ({signal_7963, signal_4671}), .b ({signal_7964, signal_4672}), .c ({signal_8163, signal_4889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4654 ( .a ({signal_7965, signal_4673}), .b ({signal_7967, signal_4675}), .c ({signal_8164, signal_4890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4655 ( .a ({signal_7965, signal_4673}), .b ({signal_7968, signal_4676}), .c ({signal_8165, signal_4891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4656 ( .a ({signal_7966, signal_4674}), .b ({signal_7969, signal_4677}), .c ({signal_8166, signal_4892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4657 ( .a ({signal_7966, signal_4674}), .b ({signal_7970, signal_4678}), .c ({signal_8167, signal_4893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4658 ( .a ({signal_7961, signal_4669}), .b ({signal_7968, signal_4676}), .c ({signal_8168, signal_4894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4659 ( .a ({signal_7971, signal_4679}), .b ({signal_7975, signal_4683}), .c ({signal_8169, signal_4895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4660 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_7976, signal_4684}), .c ({signal_8170, signal_4896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4661 ( .a ({signal_7973, signal_4681}), .b ({signal_7974, signal_4682}), .c ({signal_8171, signal_4897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4662 ( .a ({signal_7975, signal_4683}), .b ({signal_7977, signal_4685}), .c ({signal_8172, signal_4898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4663 ( .a ({signal_7975, signal_4683}), .b ({signal_7978, signal_4686}), .c ({signal_8173, signal_4899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4664 ( .a ({signal_7976, signal_4684}), .b ({signal_7979, signal_4687}), .c ({signal_8174, signal_4900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4665 ( .a ({signal_7976, signal_4684}), .b ({signal_7980, signal_4688}), .c ({signal_8175, signal_4901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4666 ( .a ({signal_7971, signal_4679}), .b ({signal_7978, signal_4686}), .c ({signal_8176, signal_4902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4667 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_8073, signal_4689}), .c ({signal_8271, signal_4903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4668 ( .a ({signal_7886, signal_4554}), .b ({signal_8073, signal_4689}), .c ({signal_8272, signal_4904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4669 ( .a ({signal_7887, signal_4555}), .b ({signal_8073, signal_4689}), .c ({signal_8273, signal_4905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4670 ( .a ({signal_8074, signal_4690}), .b ({signal_8077, signal_4693}), .c ({signal_8274, signal_4906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4671 ( .a ({signal_7881, signal_4549}), .b ({signal_8078, signal_4694}), .c ({signal_8275, signal_4907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4672 ( .a ({signal_7882, signal_4550}), .b ({signal_8079, signal_4695}), .c ({signal_8276, signal_4908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4673 ( .a ({signal_7883, signal_4551}), .b ({signal_8077, signal_4693}), .c ({signal_8277, signal_4909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4674 ( .a ({signal_7981, signal_4697}), .b ({signal_7985, signal_4701}), .c ({signal_8177, signal_4910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4675 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_7986, signal_4702}), .c ({signal_8178, signal_4911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4676 ( .a ({signal_7983, signal_4699}), .b ({signal_7984, signal_4700}), .c ({signal_8179, signal_4912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4677 ( .a ({signal_7985, signal_4701}), .b ({signal_7987, signal_4703}), .c ({signal_8180, signal_4913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4678 ( .a ({signal_7985, signal_4701}), .b ({signal_7988, signal_4704}), .c ({signal_8181, signal_4914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4679 ( .a ({signal_7986, signal_4702}), .b ({signal_7989, signal_4705}), .c ({signal_8182, signal_4915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4680 ( .a ({signal_7986, signal_4702}), .b ({signal_7990, signal_4706}), .c ({signal_8183, signal_4916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4681 ( .a ({signal_7981, signal_4697}), .b ({signal_7988, signal_4704}), .c ({signal_8184, signal_4917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4682 ( .a ({signal_7991, signal_4707}), .b ({signal_7995, signal_4711}), .c ({signal_8185, signal_4918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4683 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_7996, signal_4712}), .c ({signal_8186, signal_4919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4684 ( .a ({signal_7993, signal_4709}), .b ({signal_7994, signal_4710}), .c ({signal_8187, signal_4920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4685 ( .a ({signal_7995, signal_4711}), .b ({signal_7997, signal_4713}), .c ({signal_8188, signal_4921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4686 ( .a ({signal_7995, signal_4711}), .b ({signal_7998, signal_4714}), .c ({signal_8189, signal_4922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4687 ( .a ({signal_7996, signal_4712}), .b ({signal_7999, signal_4715}), .c ({signal_8190, signal_4923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4688 ( .a ({signal_7996, signal_4712}), .b ({signal_8000, signal_4716}), .c ({signal_8191, signal_4924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4689 ( .a ({signal_7991, signal_4707}), .b ({signal_7998, signal_4714}), .c ({signal_8192, signal_4925}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4690 ( .a ({signal_8001, signal_4717}), .b ({signal_8005, signal_4721}), .c ({signal_8193, signal_4926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4691 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_8006, signal_4722}), .c ({signal_8194, signal_4927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4692 ( .a ({signal_8003, signal_4719}), .b ({signal_8004, signal_4720}), .c ({signal_8195, signal_4928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4693 ( .a ({signal_8005, signal_4721}), .b ({signal_8007, signal_4723}), .c ({signal_8196, signal_4929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4694 ( .a ({signal_8005, signal_4721}), .b ({signal_8008, signal_4724}), .c ({signal_8197, signal_4930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4695 ( .a ({signal_8006, signal_4722}), .b ({signal_8009, signal_4725}), .c ({signal_8198, signal_4931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4696 ( .a ({signal_8006, signal_4722}), .b ({signal_8010, signal_4726}), .c ({signal_8199, signal_4932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4697 ( .a ({signal_8001, signal_4717}), .b ({signal_8008, signal_4724}), .c ({signal_8200, signal_4933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4698 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_8081, signal_4727}), .c ({signal_8278, signal_4934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4699 ( .a ({signal_7896, signal_4564}), .b ({signal_8081, signal_4727}), .c ({signal_8279, signal_4935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4700 ( .a ({signal_7897, signal_4565}), .b ({signal_8081, signal_4727}), .c ({signal_8280, signal_4936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4701 ( .a ({signal_8082, signal_4728}), .b ({signal_8085, signal_4731}), .c ({signal_8281, signal_4937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4702 ( .a ({signal_7891, signal_4559}), .b ({signal_8086, signal_4732}), .c ({signal_8282, signal_4938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4703 ( .a ({signal_7892, signal_4560}), .b ({signal_8087, signal_4733}), .c ({signal_8283, signal_4939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4704 ( .a ({signal_7893, signal_4561}), .b ({signal_8085, signal_4731}), .c ({signal_8284, signal_4940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4705 ( .a ({signal_8011, signal_4735}), .b ({signal_8015, signal_4739}), .c ({signal_8201, signal_4941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4706 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_8016, signal_4740}), .c ({signal_8202, signal_4942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4707 ( .a ({signal_8013, signal_4737}), .b ({signal_8014, signal_4738}), .c ({signal_8203, signal_4943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4708 ( .a ({signal_8015, signal_4739}), .b ({signal_8017, signal_4741}), .c ({signal_8204, signal_4944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4709 ( .a ({signal_8015, signal_4739}), .b ({signal_8018, signal_4742}), .c ({signal_8205, signal_4945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4710 ( .a ({signal_8016, signal_4740}), .b ({signal_8019, signal_4743}), .c ({signal_8206, signal_4946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4711 ( .a ({signal_8016, signal_4740}), .b ({signal_8020, signal_4744}), .c ({signal_8207, signal_4947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4712 ( .a ({signal_8011, signal_4735}), .b ({signal_8018, signal_4742}), .c ({signal_8208, signal_4948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4713 ( .a ({signal_8021, signal_4745}), .b ({signal_8025, signal_4749}), .c ({signal_8209, signal_4949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4714 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_8026, signal_4750}), .c ({signal_8210, signal_4950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4715 ( .a ({signal_8023, signal_4747}), .b ({signal_8024, signal_4748}), .c ({signal_8211, signal_4951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4716 ( .a ({signal_8025, signal_4749}), .b ({signal_8027, signal_4751}), .c ({signal_8212, signal_4952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4717 ( .a ({signal_8025, signal_4749}), .b ({signal_8028, signal_4752}), .c ({signal_8213, signal_4953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4718 ( .a ({signal_8026, signal_4750}), .b ({signal_8029, signal_4753}), .c ({signal_8214, signal_4954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4719 ( .a ({signal_8026, signal_4750}), .b ({signal_8030, signal_4754}), .c ({signal_8215, signal_4955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4720 ( .a ({signal_8021, signal_4745}), .b ({signal_8028, signal_4752}), .c ({signal_8216, signal_4956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4721 ( .a ({signal_8031, signal_4755}), .b ({signal_8035, signal_4759}), .c ({signal_8217, signal_4957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4722 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_8036, signal_4760}), .c ({signal_8218, signal_4958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4723 ( .a ({signal_8033, signal_4757}), .b ({signal_8034, signal_4758}), .c ({signal_8219, signal_4959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4724 ( .a ({signal_8035, signal_4759}), .b ({signal_8037, signal_4761}), .c ({signal_8220, signal_4960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4725 ( .a ({signal_8035, signal_4759}), .b ({signal_8038, signal_4762}), .c ({signal_8221, signal_4961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4726 ( .a ({signal_8036, signal_4760}), .b ({signal_8039, signal_4763}), .c ({signal_8222, signal_4962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4727 ( .a ({signal_8036, signal_4760}), .b ({signal_8040, signal_4764}), .c ({signal_8223, signal_4963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4728 ( .a ({signal_8031, signal_4755}), .b ({signal_8038, signal_4762}), .c ({signal_8224, signal_4964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4729 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_8089, signal_4765}), .c ({signal_8285, signal_4965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4730 ( .a ({signal_7906, signal_4574}), .b ({signal_8089, signal_4765}), .c ({signal_8286, signal_4966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4731 ( .a ({signal_7907, signal_4575}), .b ({signal_8089, signal_4765}), .c ({signal_8287, signal_4967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4732 ( .a ({signal_8090, signal_4766}), .b ({signal_8093, signal_4769}), .c ({signal_8288, signal_4968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4733 ( .a ({signal_7901, signal_4569}), .b ({signal_8094, signal_4770}), .c ({signal_8289, signal_4969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4734 ( .a ({signal_7902, signal_4570}), .b ({signal_8095, signal_4771}), .c ({signal_8290, signal_4970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4735 ( .a ({signal_7903, signal_4571}), .b ({signal_8093, signal_4769}), .c ({signal_8291, signal_4971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4736 ( .a ({signal_7610, signal_4362}), .b ({signal_8041, signal_4773}), .c ({signal_8225, signal_4972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4737 ( .a ({signal_7846, signal_4584}), .b ({signal_8041, signal_4773}), .c ({signal_8226, signal_4973}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4738 ( .a ({signal_7847, signal_4585}), .b ({signal_8041, signal_4773}), .c ({signal_8227, signal_4974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4739 ( .a ({signal_8042, signal_4774}), .b ({signal_8045, signal_4777}), .c ({signal_8228, signal_4975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4740 ( .a ({signal_7841, signal_4579}), .b ({signal_8046, signal_4778}), .c ({signal_8229, signal_4976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4741 ( .a ({signal_7842, signal_4580}), .b ({signal_8047, signal_4779}), .c ({signal_8230, signal_4977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4742 ( .a ({signal_7843, signal_4581}), .b ({signal_8045, signal_4777}), .c ({signal_8231, signal_4978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4743 ( .a ({signal_7823, signal_4370}), .b ({signal_8049, signal_4781}), .c ({signal_8232, signal_4979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4744 ( .a ({signal_7856, signal_4594}), .b ({signal_8049, signal_4781}), .c ({signal_8233, signal_4980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4745 ( .a ({signal_7857, signal_4595}), .b ({signal_8049, signal_4781}), .c ({signal_8234, signal_4981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4746 ( .a ({signal_8050, signal_4782}), .b ({signal_8053, signal_4785}), .c ({signal_8235, signal_4982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4747 ( .a ({signal_7851, signal_4589}), .b ({signal_8054, signal_4786}), .c ({signal_8236, signal_4983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4748 ( .a ({signal_7852, signal_4590}), .b ({signal_8055, signal_4787}), .c ({signal_8237, signal_4984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4749 ( .a ({signal_7853, signal_4591}), .b ({signal_8053, signal_4785}), .c ({signal_8238, signal_4985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4750 ( .a ({signal_7529, signal_4378}), .b ({signal_8057, signal_4789}), .c ({signal_8239, signal_4986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4751 ( .a ({signal_7866, signal_4604}), .b ({signal_8057, signal_4789}), .c ({signal_8240, signal_4987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4752 ( .a ({signal_7867, signal_4605}), .b ({signal_8057, signal_4789}), .c ({signal_8241, signal_4988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4753 ( .a ({signal_8058, signal_4790}), .b ({signal_8061, signal_4793}), .c ({signal_8242, signal_4989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4754 ( .a ({signal_7861, signal_4599}), .b ({signal_8062, signal_4794}), .c ({signal_8243, signal_4990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4755 ( .a ({signal_7862, signal_4600}), .b ({signal_8063, signal_4795}), .c ({signal_8244, signal_4991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4756 ( .a ({signal_7863, signal_4601}), .b ({signal_8061, signal_4793}), .c ({signal_8245, signal_4992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4757 ( .a ({signal_7637, signal_4354}), .b ({signal_8065, signal_4797}), .c ({signal_8246, signal_4993}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4758 ( .a ({signal_7876, signal_4614}), .b ({signal_8065, signal_4797}), .c ({signal_8247, signal_4994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4759 ( .a ({signal_7877, signal_4615}), .b ({signal_8065, signal_4797}), .c ({signal_8248, signal_4995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4760 ( .a ({signal_8066, signal_4798}), .b ({signal_8069, signal_4801}), .c ({signal_8249, signal_4996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4761 ( .a ({signal_7871, signal_4609}), .b ({signal_8070, signal_4802}), .c ({signal_8250, signal_4997}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4762 ( .a ({signal_7872, signal_4610}), .b ({signal_8071, signal_4803}), .c ({signal_8251, signal_4998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4763 ( .a ({signal_7873, signal_4611}), .b ({signal_8069, signal_4801}), .c ({signal_8252, signal_4999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4863 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_8121, signal_4847}), .c ({signal_8382, signal_5099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4864 ( .a ({signal_7916, signal_4624}), .b ({signal_8121, signal_4847}), .c ({signal_8383, signal_5100}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4865 ( .a ({signal_7917, signal_4625}), .b ({signal_8121, signal_4847}), .c ({signal_8384, signal_5101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4866 ( .a ({signal_8122, signal_4848}), .b ({signal_8125, signal_4851}), .c ({signal_8385, signal_5102}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4867 ( .a ({signal_7911, signal_4619}), .b ({signal_8126, signal_4852}), .c ({signal_8386, signal_5103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4868 ( .a ({signal_7912, signal_4620}), .b ({signal_8127, signal_4853}), .c ({signal_8387, signal_5104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4869 ( .a ({signal_7913, signal_4621}), .b ({signal_8125, signal_4851}), .c ({signal_8388, signal_5105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4870 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_8129, signal_4855}), .c ({signal_8389, signal_5106}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4871 ( .a ({signal_7926, signal_4634}), .b ({signal_8129, signal_4855}), .c ({signal_8390, signal_5107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4872 ( .a ({signal_7927, signal_4635}), .b ({signal_8129, signal_4855}), .c ({signal_8391, signal_5108}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4873 ( .a ({signal_8130, signal_4856}), .b ({signal_8133, signal_4859}), .c ({signal_8392, signal_5109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4874 ( .a ({signal_7921, signal_4629}), .b ({signal_8134, signal_4860}), .c ({signal_8393, signal_5110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4875 ( .a ({signal_7922, signal_4630}), .b ({signal_8135, signal_4861}), .c ({signal_8394, signal_5111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4876 ( .a ({signal_7923, signal_4631}), .b ({signal_8133, signal_4859}), .c ({signal_8395, signal_5112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4877 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_8137, signal_4863}), .c ({signal_8396, signal_5113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4878 ( .a ({signal_7936, signal_4644}), .b ({signal_8137, signal_4863}), .c ({signal_8397, signal_5114}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4879 ( .a ({signal_7937, signal_4645}), .b ({signal_8137, signal_4863}), .c ({signal_8398, signal_5115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4880 ( .a ({signal_8138, signal_4864}), .b ({signal_8141, signal_4867}), .c ({signal_8399, signal_5116}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4881 ( .a ({signal_7931, signal_4639}), .b ({signal_8142, signal_4868}), .c ({signal_8400, signal_5117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4882 ( .a ({signal_7932, signal_4640}), .b ({signal_8143, signal_4869}), .c ({signal_8401, signal_5118}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4883 ( .a ({signal_7933, signal_4641}), .b ({signal_8141, signal_4867}), .c ({signal_8402, signal_5119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4884 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_8145, signal_4871}), .c ({signal_8403, signal_5120}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4885 ( .a ({signal_7946, signal_4654}), .b ({signal_8145, signal_4871}), .c ({signal_8404, signal_5121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4886 ( .a ({signal_7947, signal_4655}), .b ({signal_8145, signal_4871}), .c ({signal_8405, signal_5122}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4887 ( .a ({signal_8146, signal_4872}), .b ({signal_8149, signal_4875}), .c ({signal_8406, signal_5123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4888 ( .a ({signal_7941, signal_4649}), .b ({signal_8150, signal_4876}), .c ({signal_8407, signal_5124}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4889 ( .a ({signal_7942, signal_4650}), .b ({signal_8151, signal_4877}), .c ({signal_8408, signal_5125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4890 ( .a ({signal_7943, signal_4651}), .b ({signal_8149, signal_4875}), .c ({signal_8409, signal_5126}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4891 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_8153, signal_4879}), .c ({signal_8410, signal_5127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4892 ( .a ({signal_7956, signal_4664}), .b ({signal_8153, signal_4879}), .c ({signal_8411, signal_5128}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4893 ( .a ({signal_7957, signal_4665}), .b ({signal_8153, signal_4879}), .c ({signal_8412, signal_5129}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4894 ( .a ({signal_8154, signal_4880}), .b ({signal_8157, signal_4883}), .c ({signal_8413, signal_5130}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4895 ( .a ({signal_7951, signal_4659}), .b ({signal_8158, signal_4884}), .c ({signal_8414, signal_5131}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4896 ( .a ({signal_7952, signal_4660}), .b ({signal_8159, signal_4885}), .c ({signal_8415, signal_5132}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4897 ( .a ({signal_7953, signal_4661}), .b ({signal_8157, signal_4883}), .c ({signal_8416, signal_5133}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4898 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_8161, signal_4887}), .c ({signal_8417, signal_5134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4899 ( .a ({signal_7966, signal_4674}), .b ({signal_8161, signal_4887}), .c ({signal_8418, signal_5135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4900 ( .a ({signal_7967, signal_4675}), .b ({signal_8161, signal_4887}), .c ({signal_8419, signal_5136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4901 ( .a ({signal_8162, signal_4888}), .b ({signal_8165, signal_4891}), .c ({signal_8420, signal_5137}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4902 ( .a ({signal_7961, signal_4669}), .b ({signal_8166, signal_4892}), .c ({signal_8421, signal_5138}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4903 ( .a ({signal_7962, signal_4670}), .b ({signal_8167, signal_4893}), .c ({signal_8422, signal_5139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4904 ( .a ({signal_7963, signal_4671}), .b ({signal_8165, signal_4891}), .c ({signal_8423, signal_5140}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4905 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_8169, signal_4895}), .c ({signal_8424, signal_5141}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4906 ( .a ({signal_7976, signal_4684}), .b ({signal_8169, signal_4895}), .c ({signal_8425, signal_5142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4907 ( .a ({signal_7977, signal_4685}), .b ({signal_8169, signal_4895}), .c ({signal_8426, signal_5143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4908 ( .a ({signal_8170, signal_4896}), .b ({signal_8173, signal_4899}), .c ({signal_8427, signal_5144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4909 ( .a ({signal_7971, signal_4679}), .b ({signal_8174, signal_4900}), .c ({signal_8428, signal_5145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4910 ( .a ({signal_7972, signal_4680}), .b ({signal_8175, signal_4901}), .c ({signal_8429, signal_5146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4911 ( .a ({signal_7973, signal_4681}), .b ({signal_8173, signal_4899}), .c ({signal_8430, signal_5147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4912 ( .a ({signal_7882, signal_4550}), .b ({signal_8272, signal_4904}), .c ({signal_8506, signal_5148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4913 ( .a ({signal_8274, signal_4906}), .b ({signal_8275, signal_4907}), .c ({signal_8507, signal_5149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4918 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_8177, signal_4910}), .c ({signal_8431, signal_5154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4919 ( .a ({signal_7986, signal_4702}), .b ({signal_8177, signal_4910}), .c ({signal_8432, signal_5155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4920 ( .a ({signal_7987, signal_4703}), .b ({signal_8177, signal_4910}), .c ({signal_8433, signal_5156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4921 ( .a ({signal_8178, signal_4911}), .b ({signal_8181, signal_4914}), .c ({signal_8434, signal_5157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4922 ( .a ({signal_7981, signal_4697}), .b ({signal_8182, signal_4915}), .c ({signal_8435, signal_5158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4923 ( .a ({signal_7982, signal_4698}), .b ({signal_8183, signal_4916}), .c ({signal_8436, signal_5159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4924 ( .a ({signal_7983, signal_4699}), .b ({signal_8181, signal_4914}), .c ({signal_8437, signal_5160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4925 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_8185, signal_4918}), .c ({signal_8438, signal_5161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4926 ( .a ({signal_7996, signal_4712}), .b ({signal_8185, signal_4918}), .c ({signal_8439, signal_5162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4927 ( .a ({signal_7997, signal_4713}), .b ({signal_8185, signal_4918}), .c ({signal_8440, signal_5163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4928 ( .a ({signal_8186, signal_4919}), .b ({signal_8189, signal_4922}), .c ({signal_8441, signal_5164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4929 ( .a ({signal_7991, signal_4707}), .b ({signal_8190, signal_4923}), .c ({signal_8442, signal_5165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4930 ( .a ({signal_7992, signal_4708}), .b ({signal_8191, signal_4924}), .c ({signal_8443, signal_5166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4931 ( .a ({signal_7993, signal_4709}), .b ({signal_8189, signal_4922}), .c ({signal_8444, signal_5167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4932 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_8193, signal_4926}), .c ({signal_8445, signal_5168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4933 ( .a ({signal_8006, signal_4722}), .b ({signal_8193, signal_4926}), .c ({signal_8446, signal_5169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4934 ( .a ({signal_8007, signal_4723}), .b ({signal_8193, signal_4926}), .c ({signal_8447, signal_5170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4935 ( .a ({signal_8194, signal_4927}), .b ({signal_8197, signal_4930}), .c ({signal_8448, signal_5171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4936 ( .a ({signal_8001, signal_4717}), .b ({signal_8198, signal_4931}), .c ({signal_8449, signal_5172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4937 ( .a ({signal_8002, signal_4718}), .b ({signal_8199, signal_4932}), .c ({signal_8450, signal_5173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4938 ( .a ({signal_8003, signal_4719}), .b ({signal_8197, signal_4930}), .c ({signal_8451, signal_5174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4939 ( .a ({signal_7892, signal_4560}), .b ({signal_8279, signal_4935}), .c ({signal_8512, signal_5175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4940 ( .a ({signal_8281, signal_4937}), .b ({signal_8282, signal_4938}), .c ({signal_8513, signal_5176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4945 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_8201, signal_4941}), .c ({signal_8452, signal_5181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4946 ( .a ({signal_8016, signal_4740}), .b ({signal_8201, signal_4941}), .c ({signal_8453, signal_5182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4947 ( .a ({signal_8017, signal_4741}), .b ({signal_8201, signal_4941}), .c ({signal_8454, signal_5183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4948 ( .a ({signal_8202, signal_4942}), .b ({signal_8205, signal_4945}), .c ({signal_8455, signal_5184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4949 ( .a ({signal_8011, signal_4735}), .b ({signal_8206, signal_4946}), .c ({signal_8456, signal_5185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4950 ( .a ({signal_8012, signal_4736}), .b ({signal_8207, signal_4947}), .c ({signal_8457, signal_5186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4951 ( .a ({signal_8013, signal_4737}), .b ({signal_8205, signal_4945}), .c ({signal_8458, signal_5187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4952 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_8209, signal_4949}), .c ({signal_8459, signal_5188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4953 ( .a ({signal_8026, signal_4750}), .b ({signal_8209, signal_4949}), .c ({signal_8460, signal_5189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4954 ( .a ({signal_8027, signal_4751}), .b ({signal_8209, signal_4949}), .c ({signal_8461, signal_5190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4955 ( .a ({signal_8210, signal_4950}), .b ({signal_8213, signal_4953}), .c ({signal_8462, signal_5191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4956 ( .a ({signal_8021, signal_4745}), .b ({signal_8214, signal_4954}), .c ({signal_8463, signal_5192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4957 ( .a ({signal_8022, signal_4746}), .b ({signal_8215, signal_4955}), .c ({signal_8464, signal_5193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4958 ( .a ({signal_8023, signal_4747}), .b ({signal_8213, signal_4953}), .c ({signal_8465, signal_5194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4959 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_8217, signal_4957}), .c ({signal_8466, signal_5195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4960 ( .a ({signal_8036, signal_4760}), .b ({signal_8217, signal_4957}), .c ({signal_8467, signal_5196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4961 ( .a ({signal_8037, signal_4761}), .b ({signal_8217, signal_4957}), .c ({signal_8468, signal_5197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4962 ( .a ({signal_8218, signal_4958}), .b ({signal_8221, signal_4961}), .c ({signal_8469, signal_5198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4963 ( .a ({signal_8031, signal_4755}), .b ({signal_8222, signal_4962}), .c ({signal_8470, signal_5199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4964 ( .a ({signal_8032, signal_4756}), .b ({signal_8223, signal_4963}), .c ({signal_8471, signal_5200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4965 ( .a ({signal_8033, signal_4757}), .b ({signal_8221, signal_4961}), .c ({signal_8472, signal_5201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4966 ( .a ({signal_7902, signal_4570}), .b ({signal_8286, signal_4966}), .c ({signal_8518, signal_5202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4967 ( .a ({signal_8288, signal_4968}), .b ({signal_8289, signal_4969}), .c ({signal_8519, signal_5203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4972 ( .a ({signal_7842, signal_4580}), .b ({signal_8226, signal_4973}), .c ({signal_8473, signal_5208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4973 ( .a ({signal_8228, signal_4975}), .b ({signal_8229, signal_4976}), .c ({signal_8474, signal_5209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4978 ( .a ({signal_7852, signal_4590}), .b ({signal_8233, signal_4980}), .c ({signal_8479, signal_5214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4979 ( .a ({signal_8235, signal_4982}), .b ({signal_8236, signal_4983}), .c ({signal_8480, signal_5215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4984 ( .a ({signal_7862, signal_4600}), .b ({signal_8240, signal_4987}), .c ({signal_8485, signal_5220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4985 ( .a ({signal_8242, signal_4989}), .b ({signal_8243, signal_4990}), .c ({signal_8486, signal_5221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4990 ( .a ({signal_7872, signal_4610}), .b ({signal_8247, signal_4994}), .c ({signal_8491, signal_5226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4991 ( .a ({signal_8249, signal_4996}), .b ({signal_8250, signal_4997}), .c ({signal_8492, signal_5227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5035 ( .a ({signal_7912, signal_4620}), .b ({signal_8383, signal_5100}), .c ({signal_8563, signal_5271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5036 ( .a ({signal_8385, signal_5102}), .b ({signal_8386, signal_5103}), .c ({signal_8564, signal_5272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5041 ( .a ({signal_7922, signal_4630}), .b ({signal_8390, signal_5107}), .c ({signal_8569, signal_5277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5042 ( .a ({signal_8392, signal_5109}), .b ({signal_8393, signal_5110}), .c ({signal_8570, signal_5278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5047 ( .a ({signal_7932, signal_4640}), .b ({signal_8397, signal_5114}), .c ({signal_8575, signal_5283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5048 ( .a ({signal_8399, signal_5116}), .b ({signal_8400, signal_5117}), .c ({signal_8576, signal_5284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5053 ( .a ({signal_7942, signal_4650}), .b ({signal_8404, signal_5121}), .c ({signal_8581, signal_5289}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5054 ( .a ({signal_8406, signal_5123}), .b ({signal_8407, signal_5124}), .c ({signal_8582, signal_5290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5059 ( .a ({signal_7952, signal_4660}), .b ({signal_8411, signal_5128}), .c ({signal_8587, signal_5295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5060 ( .a ({signal_8413, signal_5130}), .b ({signal_8414, signal_5131}), .c ({signal_8588, signal_5296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5065 ( .a ({signal_7962, signal_4670}), .b ({signal_8418, signal_5135}), .c ({signal_8593, signal_5301}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5066 ( .a ({signal_8420, signal_5137}), .b ({signal_8421, signal_5138}), .c ({signal_8594, signal_5302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5071 ( .a ({signal_7972, signal_4680}), .b ({signal_8425, signal_5142}), .c ({signal_8599, signal_5307}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5072 ( .a ({signal_8427, signal_5144}), .b ({signal_8428, signal_5145}), .c ({signal_8600, signal_5308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5082 ( .a ({signal_7982, signal_4698}), .b ({signal_8432, signal_5155}), .c ({signal_8605, signal_5318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5083 ( .a ({signal_8434, signal_5157}), .b ({signal_8435, signal_5158}), .c ({signal_8606, signal_5319}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5088 ( .a ({signal_7992, signal_4708}), .b ({signal_8439, signal_5162}), .c ({signal_8611, signal_5324}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5089 ( .a ({signal_8441, signal_5164}), .b ({signal_8442, signal_5165}), .c ({signal_8612, signal_5325}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5094 ( .a ({signal_8002, signal_4718}), .b ({signal_8446, signal_5169}), .c ({signal_8617, signal_5330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5095 ( .a ({signal_8448, signal_5171}), .b ({signal_8449, signal_5172}), .c ({signal_8618, signal_5331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5105 ( .a ({signal_8012, signal_4736}), .b ({signal_8453, signal_5182}), .c ({signal_8623, signal_5341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5106 ( .a ({signal_8455, signal_5184}), .b ({signal_8456, signal_5185}), .c ({signal_8624, signal_5342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5111 ( .a ({signal_8022, signal_4746}), .b ({signal_8460, signal_5189}), .c ({signal_8629, signal_5347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5112 ( .a ({signal_8462, signal_5191}), .b ({signal_8463, signal_5192}), .c ({signal_8630, signal_5348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5117 ( .a ({signal_8032, signal_4756}), .b ({signal_8467, signal_5196}), .c ({signal_8635, signal_5353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5118 ( .a ({signal_8469, signal_5198}), .b ({signal_8470, signal_5199}), .c ({signal_8636, signal_5354}) ) ;
    ClockGatingController #(9) cell_7581 ( .clk (clk), .rst (reset), .GatedClk (signal_12469), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4569 ( .a ({signal_8073, signal_4689}), .b ({signal_8075, signal_4691}), .clk (clk), .r (Fresh[0]), .c ({signal_8253, signal_4805}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4570 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_8078, signal_4694}), .clk (clk), .r (Fresh[1]), .c ({signal_8254, signal_4806}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4571 ( .a ({signal_7883, signal_4551}), .b ({signal_8077, signal_4693}), .clk (clk), .r (Fresh[2]), .c ({signal_8255, signal_4807}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4572 ( .a ({signal_8074, signal_4690}), .b ({signal_8079, signal_4695}), .clk (clk), .r (Fresh[3]), .c ({signal_8256, signal_4808}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4573 ( .a ({signal_7881, signal_4549}), .b ({signal_8076, signal_4692}), .clk (clk), .r (Fresh[4]), .c ({signal_8257, signal_4809}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4574 ( .a ({signal_7884, signal_4552}), .b ({signal_8080, signal_4696}), .clk (clk), .r (Fresh[5]), .c ({signal_8258, signal_4810}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4575 ( .a ({signal_8081, signal_4727}), .b ({signal_8083, signal_4729}), .clk (clk), .r (Fresh[6]), .c ({signal_8259, signal_4811}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4576 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_8086, signal_4732}), .clk (clk), .r (Fresh[7]), .c ({signal_8260, signal_4812}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4577 ( .a ({signal_7893, signal_4561}), .b ({signal_8085, signal_4731}), .clk (clk), .r (Fresh[8]), .c ({signal_8261, signal_4813}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4578 ( .a ({signal_8082, signal_4728}), .b ({signal_8087, signal_4733}), .clk (clk), .r (Fresh[9]), .c ({signal_8262, signal_4814}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4579 ( .a ({signal_7891, signal_4559}), .b ({signal_8084, signal_4730}), .clk (clk), .r (Fresh[10]), .c ({signal_8263, signal_4815}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4580 ( .a ({signal_7894, signal_4562}), .b ({signal_8088, signal_4734}), .clk (clk), .r (Fresh[11]), .c ({signal_8264, signal_4816}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4581 ( .a ({signal_8089, signal_4765}), .b ({signal_8091, signal_4767}), .clk (clk), .r (Fresh[12]), .c ({signal_8265, signal_4817}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4582 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_8094, signal_4770}), .clk (clk), .r (Fresh[13]), .c ({signal_8266, signal_4818}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4583 ( .a ({signal_7903, signal_4571}), .b ({signal_8093, signal_4769}), .clk (clk), .r (Fresh[14]), .c ({signal_8267, signal_4819}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4584 ( .a ({signal_8090, signal_4766}), .b ({signal_8095, signal_4771}), .clk (clk), .r (Fresh[15]), .c ({signal_8268, signal_4820}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4585 ( .a ({signal_7901, signal_4569}), .b ({signal_8092, signal_4768}), .clk (clk), .r (Fresh[16]), .c ({signal_8269, signal_4821}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4586 ( .a ({signal_7904, signal_4572}), .b ({signal_8096, signal_4772}), .clk (clk), .r (Fresh[17]), .c ({signal_8270, signal_4822}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4587 ( .a ({signal_8041, signal_4773}), .b ({signal_8043, signal_4775}), .clk (clk), .r (Fresh[18]), .c ({signal_8097, signal_4823}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4588 ( .a ({signal_7610, signal_4362}), .b ({signal_8046, signal_4778}), .clk (clk), .r (Fresh[19]), .c ({signal_8098, signal_4824}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4589 ( .a ({signal_7843, signal_4581}), .b ({signal_8045, signal_4777}), .clk (clk), .r (Fresh[20]), .c ({signal_8099, signal_4825}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4590 ( .a ({signal_8042, signal_4774}), .b ({signal_8047, signal_4779}), .clk (clk), .r (Fresh[21]), .c ({signal_8100, signal_4826}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4591 ( .a ({signal_7841, signal_4579}), .b ({signal_8044, signal_4776}), .clk (clk), .r (Fresh[22]), .c ({signal_8101, signal_4827}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4592 ( .a ({signal_7844, signal_4582}), .b ({signal_8048, signal_4780}), .clk (clk), .r (Fresh[23]), .c ({signal_8102, signal_4828}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4593 ( .a ({signal_8049, signal_4781}), .b ({signal_8051, signal_4783}), .clk (clk), .r (Fresh[24]), .c ({signal_8103, signal_4829}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4594 ( .a ({signal_7823, signal_4370}), .b ({signal_8054, signal_4786}), .clk (clk), .r (Fresh[25]), .c ({signal_8104, signal_4830}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4595 ( .a ({signal_7853, signal_4591}), .b ({signal_8053, signal_4785}), .clk (clk), .r (Fresh[26]), .c ({signal_8105, signal_4831}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4596 ( .a ({signal_8050, signal_4782}), .b ({signal_8055, signal_4787}), .clk (clk), .r (Fresh[27]), .c ({signal_8106, signal_4832}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4597 ( .a ({signal_7851, signal_4589}), .b ({signal_8052, signal_4784}), .clk (clk), .r (Fresh[28]), .c ({signal_8107, signal_4833}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4598 ( .a ({signal_7854, signal_4592}), .b ({signal_8056, signal_4788}), .clk (clk), .r (Fresh[29]), .c ({signal_8108, signal_4834}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4599 ( .a ({signal_8057, signal_4789}), .b ({signal_8059, signal_4791}), .clk (clk), .r (Fresh[30]), .c ({signal_8109, signal_4835}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4600 ( .a ({signal_7529, signal_4378}), .b ({signal_8062, signal_4794}), .clk (clk), .r (Fresh[31]), .c ({signal_8110, signal_4836}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4601 ( .a ({signal_7863, signal_4601}), .b ({signal_8061, signal_4793}), .clk (clk), .r (Fresh[32]), .c ({signal_8111, signal_4837}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4602 ( .a ({signal_8058, signal_4790}), .b ({signal_8063, signal_4795}), .clk (clk), .r (Fresh[33]), .c ({signal_8112, signal_4838}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4603 ( .a ({signal_7861, signal_4599}), .b ({signal_8060, signal_4792}), .clk (clk), .r (Fresh[34]), .c ({signal_8113, signal_4839}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4604 ( .a ({signal_7864, signal_4602}), .b ({signal_8064, signal_4796}), .clk (clk), .r (Fresh[35]), .c ({signal_8114, signal_4840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4605 ( .a ({signal_8065, signal_4797}), .b ({signal_8067, signal_4799}), .clk (clk), .r (Fresh[36]), .c ({signal_8115, signal_4841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4606 ( .a ({signal_7637, signal_4354}), .b ({signal_8070, signal_4802}), .clk (clk), .r (Fresh[37]), .c ({signal_8116, signal_4842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4607 ( .a ({signal_7873, signal_4611}), .b ({signal_8069, signal_4801}), .clk (clk), .r (Fresh[38]), .c ({signal_8117, signal_4843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4608 ( .a ({signal_8066, signal_4798}), .b ({signal_8071, signal_4803}), .clk (clk), .r (Fresh[39]), .c ({signal_8118, signal_4844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4609 ( .a ({signal_7871, signal_4609}), .b ({signal_8068, signal_4800}), .clk (clk), .r (Fresh[40]), .c ({signal_8119, signal_4845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4610 ( .a ({signal_7874, signal_4612}), .b ({signal_8072, signal_4804}), .clk (clk), .r (Fresh[41]), .c ({signal_8120, signal_4846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4764 ( .a ({signal_8121, signal_4847}), .b ({signal_8123, signal_4849}), .clk (clk), .r (Fresh[42]), .c ({signal_8292, signal_5000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4765 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_8126, signal_4852}), .clk (clk), .r (Fresh[43]), .c ({signal_8293, signal_5001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4766 ( .a ({signal_7913, signal_4621}), .b ({signal_8125, signal_4851}), .clk (clk), .r (Fresh[44]), .c ({signal_8294, signal_5002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4767 ( .a ({signal_8122, signal_4848}), .b ({signal_8127, signal_4853}), .clk (clk), .r (Fresh[45]), .c ({signal_8295, signal_5003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4768 ( .a ({signal_7911, signal_4619}), .b ({signal_8124, signal_4850}), .clk (clk), .r (Fresh[46]), .c ({signal_8296, signal_5004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4769 ( .a ({signal_7914, signal_4622}), .b ({signal_8128, signal_4854}), .clk (clk), .r (Fresh[47]), .c ({signal_8297, signal_5005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4770 ( .a ({signal_8129, signal_4855}), .b ({signal_8131, signal_4857}), .clk (clk), .r (Fresh[48]), .c ({signal_8298, signal_5006}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4771 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_8134, signal_4860}), .clk (clk), .r (Fresh[49]), .c ({signal_8299, signal_5007}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4772 ( .a ({signal_7923, signal_4631}), .b ({signal_8133, signal_4859}), .clk (clk), .r (Fresh[50]), .c ({signal_8300, signal_5008}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4773 ( .a ({signal_8130, signal_4856}), .b ({signal_8135, signal_4861}), .clk (clk), .r (Fresh[51]), .c ({signal_8301, signal_5009}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4774 ( .a ({signal_7921, signal_4629}), .b ({signal_8132, signal_4858}), .clk (clk), .r (Fresh[52]), .c ({signal_8302, signal_5010}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4775 ( .a ({signal_7924, signal_4632}), .b ({signal_8136, signal_4862}), .clk (clk), .r (Fresh[53]), .c ({signal_8303, signal_5011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4776 ( .a ({signal_8137, signal_4863}), .b ({signal_8139, signal_4865}), .clk (clk), .r (Fresh[54]), .c ({signal_8304, signal_5012}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4777 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_8142, signal_4868}), .clk (clk), .r (Fresh[55]), .c ({signal_8305, signal_5013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4778 ( .a ({signal_7933, signal_4641}), .b ({signal_8141, signal_4867}), .clk (clk), .r (Fresh[56]), .c ({signal_8306, signal_5014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4779 ( .a ({signal_8138, signal_4864}), .b ({signal_8143, signal_4869}), .clk (clk), .r (Fresh[57]), .c ({signal_8307, signal_5015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4780 ( .a ({signal_7931, signal_4639}), .b ({signal_8140, signal_4866}), .clk (clk), .r (Fresh[58]), .c ({signal_8308, signal_5016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4781 ( .a ({signal_7934, signal_4642}), .b ({signal_8144, signal_4870}), .clk (clk), .r (Fresh[59]), .c ({signal_8309, signal_5017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4782 ( .a ({signal_8145, signal_4871}), .b ({signal_8147, signal_4873}), .clk (clk), .r (Fresh[60]), .c ({signal_8310, signal_5018}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4783 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_8150, signal_4876}), .clk (clk), .r (Fresh[61]), .c ({signal_8311, signal_5019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4784 ( .a ({signal_7943, signal_4651}), .b ({signal_8149, signal_4875}), .clk (clk), .r (Fresh[62]), .c ({signal_8312, signal_5020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4785 ( .a ({signal_8146, signal_4872}), .b ({signal_8151, signal_4877}), .clk (clk), .r (Fresh[63]), .c ({signal_8313, signal_5021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4786 ( .a ({signal_7941, signal_4649}), .b ({signal_8148, signal_4874}), .clk (clk), .r (Fresh[64]), .c ({signal_8314, signal_5022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4787 ( .a ({signal_7944, signal_4652}), .b ({signal_8152, signal_4878}), .clk (clk), .r (Fresh[65]), .c ({signal_8315, signal_5023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4788 ( .a ({signal_8153, signal_4879}), .b ({signal_8155, signal_4881}), .clk (clk), .r (Fresh[66]), .c ({signal_8316, signal_5024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4789 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_8158, signal_4884}), .clk (clk), .r (Fresh[67]), .c ({signal_8317, signal_5025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4790 ( .a ({signal_7953, signal_4661}), .b ({signal_8157, signal_4883}), .clk (clk), .r (Fresh[68]), .c ({signal_8318, signal_5026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4791 ( .a ({signal_8154, signal_4880}), .b ({signal_8159, signal_4885}), .clk (clk), .r (Fresh[69]), .c ({signal_8319, signal_5027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4792 ( .a ({signal_7951, signal_4659}), .b ({signal_8156, signal_4882}), .clk (clk), .r (Fresh[70]), .c ({signal_8320, signal_5028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4793 ( .a ({signal_7954, signal_4662}), .b ({signal_8160, signal_4886}), .clk (clk), .r (Fresh[71]), .c ({signal_8321, signal_5029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4794 ( .a ({signal_8161, signal_4887}), .b ({signal_8163, signal_4889}), .clk (clk), .r (Fresh[72]), .c ({signal_8322, signal_5030}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4795 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_8166, signal_4892}), .clk (clk), .r (Fresh[73]), .c ({signal_8323, signal_5031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4796 ( .a ({signal_7963, signal_4671}), .b ({signal_8165, signal_4891}), .clk (clk), .r (Fresh[74]), .c ({signal_8324, signal_5032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4797 ( .a ({signal_8162, signal_4888}), .b ({signal_8167, signal_4893}), .clk (clk), .r (Fresh[75]), .c ({signal_8325, signal_5033}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4798 ( .a ({signal_7961, signal_4669}), .b ({signal_8164, signal_4890}), .clk (clk), .r (Fresh[76]), .c ({signal_8326, signal_5034}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4799 ( .a ({signal_7964, signal_4672}), .b ({signal_8168, signal_4894}), .clk (clk), .r (Fresh[77]), .c ({signal_8327, signal_5035}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4800 ( .a ({signal_8169, signal_4895}), .b ({signal_8171, signal_4897}), .clk (clk), .r (Fresh[78]), .c ({signal_8328, signal_5036}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4801 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_8174, signal_4900}), .clk (clk), .r (Fresh[79]), .c ({signal_8329, signal_5037}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4802 ( .a ({signal_7973, signal_4681}), .b ({signal_8173, signal_4899}), .clk (clk), .r (Fresh[80]), .c ({signal_8330, signal_5038}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4803 ( .a ({signal_8170, signal_4896}), .b ({signal_8175, signal_4901}), .clk (clk), .r (Fresh[81]), .c ({signal_8331, signal_5039}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4804 ( .a ({signal_7971, signal_4679}), .b ({signal_8172, signal_4898}), .clk (clk), .r (Fresh[82]), .c ({signal_8332, signal_5040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4805 ( .a ({signal_7974, signal_4682}), .b ({signal_8176, signal_4902}), .clk (clk), .r (Fresh[83]), .c ({signal_8333, signal_5041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4806 ( .a ({signal_8271, signal_4903}), .b ({signal_8276, signal_4908}), .clk (clk), .r (Fresh[84]), .c ({signal_8497, signal_5042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4807 ( .a ({signal_8274, signal_4906}), .b ({signal_8275, signal_4907}), .clk (clk), .r (Fresh[85]), .c ({signal_8498, signal_5043}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4808 ( .a ({signal_7882, signal_4550}), .b ({signal_8272, signal_4904}), .clk (clk), .r (Fresh[86]), .c ({signal_8499, signal_5044}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4809 ( .a ({signal_8177, signal_4910}), .b ({signal_8179, signal_4912}), .clk (clk), .r (Fresh[87]), .c ({signal_8334, signal_5045}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4810 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_8182, signal_4915}), .clk (clk), .r (Fresh[88]), .c ({signal_8335, signal_5046}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4811 ( .a ({signal_7983, signal_4699}), .b ({signal_8181, signal_4914}), .clk (clk), .r (Fresh[89]), .c ({signal_8336, signal_5047}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4812 ( .a ({signal_8178, signal_4911}), .b ({signal_8183, signal_4916}), .clk (clk), .r (Fresh[90]), .c ({signal_8337, signal_5048}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4813 ( .a ({signal_7981, signal_4697}), .b ({signal_8180, signal_4913}), .clk (clk), .r (Fresh[91]), .c ({signal_8338, signal_5049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4814 ( .a ({signal_7984, signal_4700}), .b ({signal_8184, signal_4917}), .clk (clk), .r (Fresh[92]), .c ({signal_8339, signal_5050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4815 ( .a ({signal_8185, signal_4918}), .b ({signal_8187, signal_4920}), .clk (clk), .r (Fresh[93]), .c ({signal_8340, signal_5051}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4816 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_8190, signal_4923}), .clk (clk), .r (Fresh[94]), .c ({signal_8341, signal_5052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4817 ( .a ({signal_7993, signal_4709}), .b ({signal_8189, signal_4922}), .clk (clk), .r (Fresh[95]), .c ({signal_8342, signal_5053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4818 ( .a ({signal_8186, signal_4919}), .b ({signal_8191, signal_4924}), .clk (clk), .r (Fresh[96]), .c ({signal_8343, signal_5054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4819 ( .a ({signal_7991, signal_4707}), .b ({signal_8188, signal_4921}), .clk (clk), .r (Fresh[97]), .c ({signal_8344, signal_5055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4820 ( .a ({signal_7994, signal_4710}), .b ({signal_8192, signal_4925}), .clk (clk), .r (Fresh[98]), .c ({signal_8345, signal_5056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4821 ( .a ({signal_8193, signal_4926}), .b ({signal_8195, signal_4928}), .clk (clk), .r (Fresh[99]), .c ({signal_8346, signal_5057}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4822 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_8198, signal_4931}), .clk (clk), .r (Fresh[100]), .c ({signal_8347, signal_5058}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4823 ( .a ({signal_8003, signal_4719}), .b ({signal_8197, signal_4930}), .clk (clk), .r (Fresh[101]), .c ({signal_8348, signal_5059}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4824 ( .a ({signal_8194, signal_4927}), .b ({signal_8199, signal_4932}), .clk (clk), .r (Fresh[102]), .c ({signal_8349, signal_5060}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4825 ( .a ({signal_8001, signal_4717}), .b ({signal_8196, signal_4929}), .clk (clk), .r (Fresh[103]), .c ({signal_8350, signal_5061}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4826 ( .a ({signal_8004, signal_4720}), .b ({signal_8200, signal_4933}), .clk (clk), .r (Fresh[104]), .c ({signal_8351, signal_5062}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4827 ( .a ({signal_8278, signal_4934}), .b ({signal_8283, signal_4939}), .clk (clk), .r (Fresh[105]), .c ({signal_8500, signal_5063}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4828 ( .a ({signal_8281, signal_4937}), .b ({signal_8282, signal_4938}), .clk (clk), .r (Fresh[106]), .c ({signal_8501, signal_5064}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4829 ( .a ({signal_7892, signal_4560}), .b ({signal_8279, signal_4935}), .clk (clk), .r (Fresh[107]), .c ({signal_8502, signal_5065}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4830 ( .a ({signal_8201, signal_4941}), .b ({signal_8203, signal_4943}), .clk (clk), .r (Fresh[108]), .c ({signal_8352, signal_5066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4831 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_8206, signal_4946}), .clk (clk), .r (Fresh[109]), .c ({signal_8353, signal_5067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4832 ( .a ({signal_8013, signal_4737}), .b ({signal_8205, signal_4945}), .clk (clk), .r (Fresh[110]), .c ({signal_8354, signal_5068}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4833 ( .a ({signal_8202, signal_4942}), .b ({signal_8207, signal_4947}), .clk (clk), .r (Fresh[111]), .c ({signal_8355, signal_5069}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4834 ( .a ({signal_8011, signal_4735}), .b ({signal_8204, signal_4944}), .clk (clk), .r (Fresh[112]), .c ({signal_8356, signal_5070}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4835 ( .a ({signal_8014, signal_4738}), .b ({signal_8208, signal_4948}), .clk (clk), .r (Fresh[113]), .c ({signal_8357, signal_5071}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4836 ( .a ({signal_8209, signal_4949}), .b ({signal_8211, signal_4951}), .clk (clk), .r (Fresh[114]), .c ({signal_8358, signal_5072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4837 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_8214, signal_4954}), .clk (clk), .r (Fresh[115]), .c ({signal_8359, signal_5073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4838 ( .a ({signal_8023, signal_4747}), .b ({signal_8213, signal_4953}), .clk (clk), .r (Fresh[116]), .c ({signal_8360, signal_5074}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4839 ( .a ({signal_8210, signal_4950}), .b ({signal_8215, signal_4955}), .clk (clk), .r (Fresh[117]), .c ({signal_8361, signal_5075}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4840 ( .a ({signal_8021, signal_4745}), .b ({signal_8212, signal_4952}), .clk (clk), .r (Fresh[118]), .c ({signal_8362, signal_5076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4841 ( .a ({signal_8024, signal_4748}), .b ({signal_8216, signal_4956}), .clk (clk), .r (Fresh[119]), .c ({signal_8363, signal_5077}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4842 ( .a ({signal_8217, signal_4957}), .b ({signal_8219, signal_4959}), .clk (clk), .r (Fresh[120]), .c ({signal_8364, signal_5078}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4843 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_8222, signal_4962}), .clk (clk), .r (Fresh[121]), .c ({signal_8365, signal_5079}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4844 ( .a ({signal_8033, signal_4757}), .b ({signal_8221, signal_4961}), .clk (clk), .r (Fresh[122]), .c ({signal_8366, signal_5080}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4845 ( .a ({signal_8218, signal_4958}), .b ({signal_8223, signal_4963}), .clk (clk), .r (Fresh[123]), .c ({signal_8367, signal_5081}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4846 ( .a ({signal_8031, signal_4755}), .b ({signal_8220, signal_4960}), .clk (clk), .r (Fresh[124]), .c ({signal_8368, signal_5082}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4847 ( .a ({signal_8034, signal_4758}), .b ({signal_8224, signal_4964}), .clk (clk), .r (Fresh[125]), .c ({signal_8369, signal_5083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4848 ( .a ({signal_8285, signal_4965}), .b ({signal_8290, signal_4970}), .clk (clk), .r (Fresh[126]), .c ({signal_8503, signal_5084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4849 ( .a ({signal_8288, signal_4968}), .b ({signal_8289, signal_4969}), .clk (clk), .r (Fresh[127]), .c ({signal_8504, signal_5085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4850 ( .a ({signal_7902, signal_4570}), .b ({signal_8286, signal_4966}), .clk (clk), .r (Fresh[128]), .c ({signal_8505, signal_5086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4851 ( .a ({signal_8225, signal_4972}), .b ({signal_8230, signal_4977}), .clk (clk), .r (Fresh[129]), .c ({signal_8370, signal_5087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4852 ( .a ({signal_8228, signal_4975}), .b ({signal_8229, signal_4976}), .clk (clk), .r (Fresh[130]), .c ({signal_8371, signal_5088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4853 ( .a ({signal_7842, signal_4580}), .b ({signal_8226, signal_4973}), .clk (clk), .r (Fresh[131]), .c ({signal_8372, signal_5089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4854 ( .a ({signal_8232, signal_4979}), .b ({signal_8237, signal_4984}), .clk (clk), .r (Fresh[132]), .c ({signal_8373, signal_5090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4855 ( .a ({signal_8235, signal_4982}), .b ({signal_8236, signal_4983}), .clk (clk), .r (Fresh[133]), .c ({signal_8374, signal_5091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4856 ( .a ({signal_7852, signal_4590}), .b ({signal_8233, signal_4980}), .clk (clk), .r (Fresh[134]), .c ({signal_8375, signal_5092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4857 ( .a ({signal_8239, signal_4986}), .b ({signal_8244, signal_4991}), .clk (clk), .r (Fresh[135]), .c ({signal_8376, signal_5093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4858 ( .a ({signal_8242, signal_4989}), .b ({signal_8243, signal_4990}), .clk (clk), .r (Fresh[136]), .c ({signal_8377, signal_5094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4859 ( .a ({signal_7862, signal_4600}), .b ({signal_8240, signal_4987}), .clk (clk), .r (Fresh[137]), .c ({signal_8378, signal_5095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4860 ( .a ({signal_8246, signal_4993}), .b ({signal_8251, signal_4998}), .clk (clk), .r (Fresh[138]), .c ({signal_8379, signal_5096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4861 ( .a ({signal_8249, signal_4996}), .b ({signal_8250, signal_4997}), .clk (clk), .r (Fresh[139]), .c ({signal_8380, signal_5097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4862 ( .a ({signal_7872, signal_4610}), .b ({signal_8247, signal_4994}), .clk (clk), .r (Fresh[140]), .c ({signal_8381, signal_5098}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4914 ( .a ({signal_8273, signal_4905}), .b ({signal_8253, signal_4805}), .c ({signal_8508, signal_5150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4915 ( .a ({signal_8253, signal_4805}), .b ({signal_8254, signal_4806}), .c ({signal_8509, signal_5151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4916 ( .a ({signal_8277, signal_4909}), .b ({signal_8255, signal_4807}), .c ({signal_8510, signal_5152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4917 ( .a ({signal_8257, signal_4809}), .b ({signal_8258, signal_4810}), .c ({signal_8511, signal_5153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4941 ( .a ({signal_8280, signal_4936}), .b ({signal_8259, signal_4811}), .c ({signal_8514, signal_5177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4942 ( .a ({signal_8259, signal_4811}), .b ({signal_8260, signal_4812}), .c ({signal_8515, signal_5178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4943 ( .a ({signal_8284, signal_4940}), .b ({signal_8261, signal_4813}), .c ({signal_8516, signal_5179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4944 ( .a ({signal_8263, signal_4815}), .b ({signal_8264, signal_4816}), .c ({signal_8517, signal_5180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4968 ( .a ({signal_8287, signal_4967}), .b ({signal_8265, signal_4817}), .c ({signal_8520, signal_5204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4969 ( .a ({signal_8265, signal_4817}), .b ({signal_8266, signal_4818}), .c ({signal_8521, signal_5205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4970 ( .a ({signal_8291, signal_4971}), .b ({signal_8267, signal_4819}), .c ({signal_8522, signal_5206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4971 ( .a ({signal_8269, signal_4821}), .b ({signal_8270, signal_4822}), .c ({signal_8523, signal_5207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4974 ( .a ({signal_8227, signal_4974}), .b ({signal_8097, signal_4823}), .c ({signal_8475, signal_5210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4975 ( .a ({signal_8097, signal_4823}), .b ({signal_8098, signal_4824}), .c ({signal_8476, signal_5211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4976 ( .a ({signal_8231, signal_4978}), .b ({signal_8099, signal_4825}), .c ({signal_8477, signal_5212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4977 ( .a ({signal_8101, signal_4827}), .b ({signal_8102, signal_4828}), .c ({signal_8478, signal_5213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4980 ( .a ({signal_8234, signal_4981}), .b ({signal_8103, signal_4829}), .c ({signal_8481, signal_5216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4981 ( .a ({signal_8103, signal_4829}), .b ({signal_8104, signal_4830}), .c ({signal_8482, signal_5217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4982 ( .a ({signal_8238, signal_4985}), .b ({signal_8105, signal_4831}), .c ({signal_8483, signal_5218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4983 ( .a ({signal_8107, signal_4833}), .b ({signal_8108, signal_4834}), .c ({signal_8484, signal_5219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4986 ( .a ({signal_8241, signal_4988}), .b ({signal_8109, signal_4835}), .c ({signal_8487, signal_5222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4987 ( .a ({signal_8109, signal_4835}), .b ({signal_8110, signal_4836}), .c ({signal_8488, signal_5223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4988 ( .a ({signal_8245, signal_4992}), .b ({signal_8111, signal_4837}), .c ({signal_8489, signal_5224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4989 ( .a ({signal_8113, signal_4839}), .b ({signal_8114, signal_4840}), .c ({signal_8490, signal_5225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4992 ( .a ({signal_8248, signal_4995}), .b ({signal_8115, signal_4841}), .c ({signal_8493, signal_5228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4993 ( .a ({signal_8115, signal_4841}), .b ({signal_8116, signal_4842}), .c ({signal_8494, signal_5229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4994 ( .a ({signal_8252, signal_4999}), .b ({signal_8117, signal_4843}), .c ({signal_8495, signal_5230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_4995 ( .a ({signal_8119, signal_4845}), .b ({signal_8120, signal_4846}), .c ({signal_8496, signal_5231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4996 ( .a ({signal_8382, signal_5099}), .b ({signal_8387, signal_5104}), .clk (clk), .r (Fresh[141]), .c ({signal_8524, signal_5232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4997 ( .a ({signal_8385, signal_5102}), .b ({signal_8386, signal_5103}), .clk (clk), .r (Fresh[142]), .c ({signal_8525, signal_5233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4998 ( .a ({signal_7912, signal_4620}), .b ({signal_8383, signal_5100}), .clk (clk), .r (Fresh[143]), .c ({signal_8526, signal_5234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_4999 ( .a ({signal_8389, signal_5106}), .b ({signal_8394, signal_5111}), .clk (clk), .r (Fresh[144]), .c ({signal_8527, signal_5235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5000 ( .a ({signal_8392, signal_5109}), .b ({signal_8393, signal_5110}), .clk (clk), .r (Fresh[145]), .c ({signal_8528, signal_5236}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5001 ( .a ({signal_7922, signal_4630}), .b ({signal_8390, signal_5107}), .clk (clk), .r (Fresh[146]), .c ({signal_8529, signal_5237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5002 ( .a ({signal_8396, signal_5113}), .b ({signal_8401, signal_5118}), .clk (clk), .r (Fresh[147]), .c ({signal_8530, signal_5238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5003 ( .a ({signal_8399, signal_5116}), .b ({signal_8400, signal_5117}), .clk (clk), .r (Fresh[148]), .c ({signal_8531, signal_5239}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5004 ( .a ({signal_7932, signal_4640}), .b ({signal_8397, signal_5114}), .clk (clk), .r (Fresh[149]), .c ({signal_8532, signal_5240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5005 ( .a ({signal_8403, signal_5120}), .b ({signal_8408, signal_5125}), .clk (clk), .r (Fresh[150]), .c ({signal_8533, signal_5241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5006 ( .a ({signal_8406, signal_5123}), .b ({signal_8407, signal_5124}), .clk (clk), .r (Fresh[151]), .c ({signal_8534, signal_5242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5007 ( .a ({signal_7942, signal_4650}), .b ({signal_8404, signal_5121}), .clk (clk), .r (Fresh[152]), .c ({signal_8535, signal_5243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5008 ( .a ({signal_8410, signal_5127}), .b ({signal_8415, signal_5132}), .clk (clk), .r (Fresh[153]), .c ({signal_8536, signal_5244}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5009 ( .a ({signal_8413, signal_5130}), .b ({signal_8414, signal_5131}), .clk (clk), .r (Fresh[154]), .c ({signal_8537, signal_5245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5010 ( .a ({signal_7952, signal_4660}), .b ({signal_8411, signal_5128}), .clk (clk), .r (Fresh[155]), .c ({signal_8538, signal_5246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5011 ( .a ({signal_8417, signal_5134}), .b ({signal_8422, signal_5139}), .clk (clk), .r (Fresh[156]), .c ({signal_8539, signal_5247}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5012 ( .a ({signal_8420, signal_5137}), .b ({signal_8421, signal_5138}), .clk (clk), .r (Fresh[157]), .c ({signal_8540, signal_5248}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5013 ( .a ({signal_7962, signal_4670}), .b ({signal_8418, signal_5135}), .clk (clk), .r (Fresh[158]), .c ({signal_8541, signal_5249}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5014 ( .a ({signal_8424, signal_5141}), .b ({signal_8429, signal_5146}), .clk (clk), .r (Fresh[159]), .c ({signal_8542, signal_5250}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5015 ( .a ({signal_8427, signal_5144}), .b ({signal_8428, signal_5145}), .clk (clk), .r (Fresh[160]), .c ({signal_8543, signal_5251}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5016 ( .a ({signal_7972, signal_4680}), .b ({signal_8425, signal_5142}), .clk (clk), .r (Fresh[161]), .c ({signal_8544, signal_5252}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5017 ( .a ({signal_8431, signal_5154}), .b ({signal_8436, signal_5159}), .clk (clk), .r (Fresh[162]), .c ({signal_8545, signal_5253}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5018 ( .a ({signal_8434, signal_5157}), .b ({signal_8435, signal_5158}), .clk (clk), .r (Fresh[163]), .c ({signal_8546, signal_5254}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5019 ( .a ({signal_7982, signal_4698}), .b ({signal_8432, signal_5155}), .clk (clk), .r (Fresh[164]), .c ({signal_8547, signal_5255}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5020 ( .a ({signal_8438, signal_5161}), .b ({signal_8443, signal_5166}), .clk (clk), .r (Fresh[165]), .c ({signal_8548, signal_5256}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5021 ( .a ({signal_8441, signal_5164}), .b ({signal_8442, signal_5165}), .clk (clk), .r (Fresh[166]), .c ({signal_8549, signal_5257}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5022 ( .a ({signal_7992, signal_4708}), .b ({signal_8439, signal_5162}), .clk (clk), .r (Fresh[167]), .c ({signal_8550, signal_5258}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5023 ( .a ({signal_8445, signal_5168}), .b ({signal_8450, signal_5173}), .clk (clk), .r (Fresh[168]), .c ({signal_8551, signal_5259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5024 ( .a ({signal_8448, signal_5171}), .b ({signal_8449, signal_5172}), .clk (clk), .r (Fresh[169]), .c ({signal_8552, signal_5260}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5025 ( .a ({signal_8002, signal_4718}), .b ({signal_8446, signal_5169}), .clk (clk), .r (Fresh[170]), .c ({signal_8553, signal_5261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5026 ( .a ({signal_8452, signal_5181}), .b ({signal_8457, signal_5186}), .clk (clk), .r (Fresh[171]), .c ({signal_8554, signal_5262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5027 ( .a ({signal_8455, signal_5184}), .b ({signal_8456, signal_5185}), .clk (clk), .r (Fresh[172]), .c ({signal_8555, signal_5263}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5028 ( .a ({signal_8012, signal_4736}), .b ({signal_8453, signal_5182}), .clk (clk), .r (Fresh[173]), .c ({signal_8556, signal_5264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5029 ( .a ({signal_8459, signal_5188}), .b ({signal_8464, signal_5193}), .clk (clk), .r (Fresh[174]), .c ({signal_8557, signal_5265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5030 ( .a ({signal_8462, signal_5191}), .b ({signal_8463, signal_5192}), .clk (clk), .r (Fresh[175]), .c ({signal_8558, signal_5266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5031 ( .a ({signal_8022, signal_4746}), .b ({signal_8460, signal_5189}), .clk (clk), .r (Fresh[176]), .c ({signal_8559, signal_5267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5032 ( .a ({signal_8466, signal_5195}), .b ({signal_8471, signal_5200}), .clk (clk), .r (Fresh[177]), .c ({signal_8560, signal_5268}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5033 ( .a ({signal_8469, signal_5198}), .b ({signal_8470, signal_5199}), .clk (clk), .r (Fresh[178]), .c ({signal_8561, signal_5269}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5034 ( .a ({signal_8032, signal_4756}), .b ({signal_8467, signal_5196}), .clk (clk), .r (Fresh[179]), .c ({signal_8562, signal_5270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5037 ( .a ({signal_8384, signal_5101}), .b ({signal_8292, signal_5000}), .c ({signal_8565, signal_5273}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5038 ( .a ({signal_8292, signal_5000}), .b ({signal_8293, signal_5001}), .c ({signal_8566, signal_5274}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5039 ( .a ({signal_8388, signal_5105}), .b ({signal_8294, signal_5002}), .c ({signal_8567, signal_5275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5040 ( .a ({signal_8296, signal_5004}), .b ({signal_8297, signal_5005}), .c ({signal_8568, signal_5276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5043 ( .a ({signal_8391, signal_5108}), .b ({signal_8298, signal_5006}), .c ({signal_8571, signal_5279}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5044 ( .a ({signal_8298, signal_5006}), .b ({signal_8299, signal_5007}), .c ({signal_8572, signal_5280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5045 ( .a ({signal_8395, signal_5112}), .b ({signal_8300, signal_5008}), .c ({signal_8573, signal_5281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5046 ( .a ({signal_8302, signal_5010}), .b ({signal_8303, signal_5011}), .c ({signal_8574, signal_5282}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5049 ( .a ({signal_8398, signal_5115}), .b ({signal_8304, signal_5012}), .c ({signal_8577, signal_5285}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5050 ( .a ({signal_8304, signal_5012}), .b ({signal_8305, signal_5013}), .c ({signal_8578, signal_5286}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5051 ( .a ({signal_8402, signal_5119}), .b ({signal_8306, signal_5014}), .c ({signal_8579, signal_5287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5052 ( .a ({signal_8308, signal_5016}), .b ({signal_8309, signal_5017}), .c ({signal_8580, signal_5288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5055 ( .a ({signal_8405, signal_5122}), .b ({signal_8310, signal_5018}), .c ({signal_8583, signal_5291}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5056 ( .a ({signal_8310, signal_5018}), .b ({signal_8311, signal_5019}), .c ({signal_8584, signal_5292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5057 ( .a ({signal_8409, signal_5126}), .b ({signal_8312, signal_5020}), .c ({signal_8585, signal_5293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5058 ( .a ({signal_8314, signal_5022}), .b ({signal_8315, signal_5023}), .c ({signal_8586, signal_5294}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5061 ( .a ({signal_8412, signal_5129}), .b ({signal_8316, signal_5024}), .c ({signal_8589, signal_5297}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5062 ( .a ({signal_8316, signal_5024}), .b ({signal_8317, signal_5025}), .c ({signal_8590, signal_5298}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5063 ( .a ({signal_8416, signal_5133}), .b ({signal_8318, signal_5026}), .c ({signal_8591, signal_5299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5064 ( .a ({signal_8320, signal_5028}), .b ({signal_8321, signal_5029}), .c ({signal_8592, signal_5300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5067 ( .a ({signal_8419, signal_5136}), .b ({signal_8322, signal_5030}), .c ({signal_8595, signal_5303}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5068 ( .a ({signal_8322, signal_5030}), .b ({signal_8323, signal_5031}), .c ({signal_8596, signal_5304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5069 ( .a ({signal_8423, signal_5140}), .b ({signal_8324, signal_5032}), .c ({signal_8597, signal_5305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5070 ( .a ({signal_8326, signal_5034}), .b ({signal_8327, signal_5035}), .c ({signal_8598, signal_5306}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5073 ( .a ({signal_8426, signal_5143}), .b ({signal_8328, signal_5036}), .c ({signal_8601, signal_5309}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5074 ( .a ({signal_8328, signal_5036}), .b ({signal_8329, signal_5037}), .c ({signal_8602, signal_5310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5075 ( .a ({signal_8430, signal_5147}), .b ({signal_8330, signal_5038}), .c ({signal_8603, signal_5311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5076 ( .a ({signal_8332, signal_5040}), .b ({signal_8333, signal_5041}), .c ({signal_8604, signal_5312}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5077 ( .a ({signal_8255, signal_4807}), .b ({signal_8498, signal_5043}), .c ({signal_8661, signal_5313}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5078 ( .a ({signal_8257, signal_4809}), .b ({signal_8499, signal_5044}), .c ({signal_8662, signal_5314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5079 ( .a ({signal_8497, signal_5042}), .b ({signal_8508, signal_5150}), .c ({signal_8663, signal_5315}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5080 ( .a ({signal_8506, signal_5148}), .b ({signal_8509, signal_5151}), .c ({signal_8664, signal_5316}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5081 ( .a ({signal_8256, signal_4808}), .b ({signal_8510, signal_5152}), .c ({signal_8665, signal_5317}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5084 ( .a ({signal_8433, signal_5156}), .b ({signal_8334, signal_5045}), .c ({signal_8607, signal_5320}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5085 ( .a ({signal_8334, signal_5045}), .b ({signal_8335, signal_5046}), .c ({signal_8608, signal_5321}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5086 ( .a ({signal_8437, signal_5160}), .b ({signal_8336, signal_5047}), .c ({signal_8609, signal_5322}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5087 ( .a ({signal_8338, signal_5049}), .b ({signal_8339, signal_5050}), .c ({signal_8610, signal_5323}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5090 ( .a ({signal_8440, signal_5163}), .b ({signal_8340, signal_5051}), .c ({signal_8613, signal_5326}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5091 ( .a ({signal_8340, signal_5051}), .b ({signal_8341, signal_5052}), .c ({signal_8614, signal_5327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5092 ( .a ({signal_8444, signal_5167}), .b ({signal_8342, signal_5053}), .c ({signal_8615, signal_5328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5093 ( .a ({signal_8344, signal_5055}), .b ({signal_8345, signal_5056}), .c ({signal_8616, signal_5329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5096 ( .a ({signal_8447, signal_5170}), .b ({signal_8346, signal_5057}), .c ({signal_8619, signal_5332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5097 ( .a ({signal_8346, signal_5057}), .b ({signal_8347, signal_5058}), .c ({signal_8620, signal_5333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5098 ( .a ({signal_8451, signal_5174}), .b ({signal_8348, signal_5059}), .c ({signal_8621, signal_5334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5099 ( .a ({signal_8350, signal_5061}), .b ({signal_8351, signal_5062}), .c ({signal_8622, signal_5335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5100 ( .a ({signal_8261, signal_4813}), .b ({signal_8501, signal_5064}), .c ({signal_8666, signal_5336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5101 ( .a ({signal_8263, signal_4815}), .b ({signal_8502, signal_5065}), .c ({signal_8667, signal_5337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5102 ( .a ({signal_8500, signal_5063}), .b ({signal_8514, signal_5177}), .c ({signal_8668, signal_5338}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5103 ( .a ({signal_8512, signal_5175}), .b ({signal_8515, signal_5178}), .c ({signal_8669, signal_5339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5104 ( .a ({signal_8262, signal_4814}), .b ({signal_8516, signal_5179}), .c ({signal_8670, signal_5340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5107 ( .a ({signal_8454, signal_5183}), .b ({signal_8352, signal_5066}), .c ({signal_8625, signal_5343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5108 ( .a ({signal_8352, signal_5066}), .b ({signal_8353, signal_5067}), .c ({signal_8626, signal_5344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5109 ( .a ({signal_8458, signal_5187}), .b ({signal_8354, signal_5068}), .c ({signal_8627, signal_5345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5110 ( .a ({signal_8356, signal_5070}), .b ({signal_8357, signal_5071}), .c ({signal_8628, signal_5346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5113 ( .a ({signal_8461, signal_5190}), .b ({signal_8358, signal_5072}), .c ({signal_8631, signal_5349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5114 ( .a ({signal_8358, signal_5072}), .b ({signal_8359, signal_5073}), .c ({signal_8632, signal_5350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5115 ( .a ({signal_8465, signal_5194}), .b ({signal_8360, signal_5074}), .c ({signal_8633, signal_5351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5116 ( .a ({signal_8362, signal_5076}), .b ({signal_8363, signal_5077}), .c ({signal_8634, signal_5352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5119 ( .a ({signal_8468, signal_5197}), .b ({signal_8364, signal_5078}), .c ({signal_8637, signal_5355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5120 ( .a ({signal_8364, signal_5078}), .b ({signal_8365, signal_5079}), .c ({signal_8638, signal_5356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5121 ( .a ({signal_8472, signal_5201}), .b ({signal_8366, signal_5080}), .c ({signal_8639, signal_5357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5122 ( .a ({signal_8368, signal_5082}), .b ({signal_8369, signal_5083}), .c ({signal_8640, signal_5358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5123 ( .a ({signal_8267, signal_4819}), .b ({signal_8504, signal_5085}), .c ({signal_8671, signal_5359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5124 ( .a ({signal_8269, signal_4821}), .b ({signal_8505, signal_5086}), .c ({signal_8672, signal_5360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5125 ( .a ({signal_8503, signal_5084}), .b ({signal_8520, signal_5204}), .c ({signal_8673, signal_5361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5126 ( .a ({signal_8518, signal_5202}), .b ({signal_8521, signal_5205}), .c ({signal_8674, signal_5362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5127 ( .a ({signal_8268, signal_4820}), .b ({signal_8522, signal_5206}), .c ({signal_8675, signal_5363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5128 ( .a ({signal_8099, signal_4825}), .b ({signal_8371, signal_5088}), .c ({signal_8641, signal_5364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5129 ( .a ({signal_8101, signal_4827}), .b ({signal_8372, signal_5089}), .c ({signal_8642, signal_5365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5130 ( .a ({signal_8370, signal_5087}), .b ({signal_8475, signal_5210}), .c ({signal_8643, signal_5366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5131 ( .a ({signal_8473, signal_5208}), .b ({signal_8476, signal_5211}), .c ({signal_8644, signal_5367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5132 ( .a ({signal_8100, signal_4826}), .b ({signal_8477, signal_5212}), .c ({signal_8645, signal_5368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5133 ( .a ({signal_8105, signal_4831}), .b ({signal_8374, signal_5091}), .c ({signal_8646, signal_5369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5134 ( .a ({signal_8107, signal_4833}), .b ({signal_8375, signal_5092}), .c ({signal_8647, signal_5370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5135 ( .a ({signal_8373, signal_5090}), .b ({signal_8481, signal_5216}), .c ({signal_8648, signal_5371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5136 ( .a ({signal_8479, signal_5214}), .b ({signal_8482, signal_5217}), .c ({signal_8649, signal_5372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5137 ( .a ({signal_8106, signal_4832}), .b ({signal_8483, signal_5218}), .c ({signal_8650, signal_5373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5138 ( .a ({signal_8111, signal_4837}), .b ({signal_8377, signal_5094}), .c ({signal_8651, signal_5374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5139 ( .a ({signal_8113, signal_4839}), .b ({signal_8378, signal_5095}), .c ({signal_8652, signal_5375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5140 ( .a ({signal_8376, signal_5093}), .b ({signal_8487, signal_5222}), .c ({signal_8653, signal_5376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5141 ( .a ({signal_8485, signal_5220}), .b ({signal_8488, signal_5223}), .c ({signal_8654, signal_5377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5142 ( .a ({signal_8112, signal_4838}), .b ({signal_8489, signal_5224}), .c ({signal_8655, signal_5378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5143 ( .a ({signal_8117, signal_4843}), .b ({signal_8380, signal_5097}), .c ({signal_8656, signal_5379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5144 ( .a ({signal_8119, signal_4845}), .b ({signal_8381, signal_5098}), .c ({signal_8657, signal_5380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5145 ( .a ({signal_8379, signal_5096}), .b ({signal_8493, signal_5228}), .c ({signal_8658, signal_5381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5146 ( .a ({signal_8491, signal_5226}), .b ({signal_8494, signal_5229}), .c ({signal_8659, signal_5382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5147 ( .a ({signal_8118, signal_4844}), .b ({signal_8495, signal_5230}), .c ({signal_8660, signal_5383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5148 ( .a ({signal_8294, signal_5002}), .b ({signal_8525, signal_5233}), .c ({signal_8676, signal_5384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5149 ( .a ({signal_8296, signal_5004}), .b ({signal_8526, signal_5234}), .c ({signal_8677, signal_5385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5150 ( .a ({signal_8524, signal_5232}), .b ({signal_8565, signal_5273}), .c ({signal_8678, signal_5386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5151 ( .a ({signal_8563, signal_5271}), .b ({signal_8566, signal_5274}), .c ({signal_8679, signal_5387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5152 ( .a ({signal_8295, signal_5003}), .b ({signal_8567, signal_5275}), .c ({signal_8680, signal_5388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5153 ( .a ({signal_8300, signal_5008}), .b ({signal_8528, signal_5236}), .c ({signal_8681, signal_5389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5154 ( .a ({signal_8302, signal_5010}), .b ({signal_8529, signal_5237}), .c ({signal_8682, signal_5390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5155 ( .a ({signal_8527, signal_5235}), .b ({signal_8571, signal_5279}), .c ({signal_8683, signal_5391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5156 ( .a ({signal_8569, signal_5277}), .b ({signal_8572, signal_5280}), .c ({signal_8684, signal_5392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5157 ( .a ({signal_8301, signal_5009}), .b ({signal_8573, signal_5281}), .c ({signal_8685, signal_5393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5158 ( .a ({signal_8306, signal_5014}), .b ({signal_8531, signal_5239}), .c ({signal_8686, signal_5394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5159 ( .a ({signal_8308, signal_5016}), .b ({signal_8532, signal_5240}), .c ({signal_8687, signal_5395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5160 ( .a ({signal_8530, signal_5238}), .b ({signal_8577, signal_5285}), .c ({signal_8688, signal_5396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5161 ( .a ({signal_8575, signal_5283}), .b ({signal_8578, signal_5286}), .c ({signal_8689, signal_5397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5162 ( .a ({signal_8307, signal_5015}), .b ({signal_8579, signal_5287}), .c ({signal_8690, signal_5398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5163 ( .a ({signal_8312, signal_5020}), .b ({signal_8534, signal_5242}), .c ({signal_8691, signal_5399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5164 ( .a ({signal_8314, signal_5022}), .b ({signal_8535, signal_5243}), .c ({signal_8692, signal_5400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5165 ( .a ({signal_8533, signal_5241}), .b ({signal_8583, signal_5291}), .c ({signal_8693, signal_5401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5166 ( .a ({signal_8581, signal_5289}), .b ({signal_8584, signal_5292}), .c ({signal_8694, signal_5402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5167 ( .a ({signal_8313, signal_5021}), .b ({signal_8585, signal_5293}), .c ({signal_8695, signal_5403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5168 ( .a ({signal_8318, signal_5026}), .b ({signal_8537, signal_5245}), .c ({signal_8696, signal_5404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5169 ( .a ({signal_8320, signal_5028}), .b ({signal_8538, signal_5246}), .c ({signal_8697, signal_5405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5170 ( .a ({signal_8536, signal_5244}), .b ({signal_8589, signal_5297}), .c ({signal_8698, signal_5406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5171 ( .a ({signal_8587, signal_5295}), .b ({signal_8590, signal_5298}), .c ({signal_8699, signal_5407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5172 ( .a ({signal_8319, signal_5027}), .b ({signal_8591, signal_5299}), .c ({signal_8700, signal_5408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5173 ( .a ({signal_8324, signal_5032}), .b ({signal_8540, signal_5248}), .c ({signal_8701, signal_5409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5174 ( .a ({signal_8326, signal_5034}), .b ({signal_8541, signal_5249}), .c ({signal_8702, signal_5410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5175 ( .a ({signal_8539, signal_5247}), .b ({signal_8595, signal_5303}), .c ({signal_8703, signal_5411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5176 ( .a ({signal_8593, signal_5301}), .b ({signal_8596, signal_5304}), .c ({signal_8704, signal_5412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5177 ( .a ({signal_8325, signal_5033}), .b ({signal_8597, signal_5305}), .c ({signal_8705, signal_5413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5178 ( .a ({signal_8330, signal_5038}), .b ({signal_8543, signal_5251}), .c ({signal_8706, signal_5414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5179 ( .a ({signal_8332, signal_5040}), .b ({signal_8544, signal_5252}), .c ({signal_8707, signal_5415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5180 ( .a ({signal_8542, signal_5250}), .b ({signal_8601, signal_5309}), .c ({signal_8708, signal_5416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5181 ( .a ({signal_8599, signal_5307}), .b ({signal_8602, signal_5310}), .c ({signal_8709, signal_5417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5182 ( .a ({signal_8331, signal_5039}), .b ({signal_8603, signal_5311}), .c ({signal_8710, signal_5418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5183 ( .a ({signal_8661, signal_5313}), .b ({signal_8662, signal_5314}), .c ({signal_8757, signal_5419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5184 ( .a ({signal_8511, signal_5153}), .b ({signal_8663, signal_5315}), .c ({signal_8758, signal_5420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5185 ( .a ({signal_8662, signal_5314}), .b ({signal_8664, signal_5316}), .c ({signal_8759, signal_5421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5186 ( .a ({signal_8511, signal_5153}), .b ({signal_8665, signal_5317}), .c ({signal_8760, signal_5422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5187 ( .a ({signal_8336, signal_5047}), .b ({signal_8546, signal_5254}), .c ({signal_8711, signal_5423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5188 ( .a ({signal_8338, signal_5049}), .b ({signal_8547, signal_5255}), .c ({signal_8712, signal_5424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5189 ( .a ({signal_8545, signal_5253}), .b ({signal_8607, signal_5320}), .c ({signal_8713, signal_5425}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5190 ( .a ({signal_8605, signal_5318}), .b ({signal_8608, signal_5321}), .c ({signal_8714, signal_5426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5191 ( .a ({signal_8337, signal_5048}), .b ({signal_8609, signal_5322}), .c ({signal_8715, signal_5427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5192 ( .a ({signal_8342, signal_5053}), .b ({signal_8549, signal_5257}), .c ({signal_8716, signal_5428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5193 ( .a ({signal_8344, signal_5055}), .b ({signal_8550, signal_5258}), .c ({signal_8717, signal_5429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5194 ( .a ({signal_8548, signal_5256}), .b ({signal_8613, signal_5326}), .c ({signal_8718, signal_5430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5195 ( .a ({signal_8611, signal_5324}), .b ({signal_8614, signal_5327}), .c ({signal_8719, signal_5431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5196 ( .a ({signal_8343, signal_5054}), .b ({signal_8615, signal_5328}), .c ({signal_8720, signal_5432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5197 ( .a ({signal_8348, signal_5059}), .b ({signal_8552, signal_5260}), .c ({signal_8721, signal_5433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5198 ( .a ({signal_8350, signal_5061}), .b ({signal_8553, signal_5261}), .c ({signal_8722, signal_5434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5199 ( .a ({signal_8551, signal_5259}), .b ({signal_8619, signal_5332}), .c ({signal_8723, signal_5435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5200 ( .a ({signal_8617, signal_5330}), .b ({signal_8620, signal_5333}), .c ({signal_8724, signal_5436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5201 ( .a ({signal_8349, signal_5060}), .b ({signal_8621, signal_5334}), .c ({signal_8725, signal_5437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5202 ( .a ({signal_8666, signal_5336}), .b ({signal_8667, signal_5337}), .c ({signal_8761, signal_5438}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5203 ( .a ({signal_8517, signal_5180}), .b ({signal_8668, signal_5338}), .c ({signal_8762, signal_5439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5204 ( .a ({signal_8667, signal_5337}), .b ({signal_8669, signal_5339}), .c ({signal_8763, signal_5440}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5205 ( .a ({signal_8517, signal_5180}), .b ({signal_8670, signal_5340}), .c ({signal_8764, signal_5441}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5206 ( .a ({signal_8354, signal_5068}), .b ({signal_8555, signal_5263}), .c ({signal_8726, signal_5442}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5207 ( .a ({signal_8356, signal_5070}), .b ({signal_8556, signal_5264}), .c ({signal_8727, signal_5443}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5208 ( .a ({signal_8554, signal_5262}), .b ({signal_8625, signal_5343}), .c ({signal_8728, signal_5444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5209 ( .a ({signal_8623, signal_5341}), .b ({signal_8626, signal_5344}), .c ({signal_8729, signal_5445}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5210 ( .a ({signal_8355, signal_5069}), .b ({signal_8627, signal_5345}), .c ({signal_8730, signal_5446}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5211 ( .a ({signal_8360, signal_5074}), .b ({signal_8558, signal_5266}), .c ({signal_8731, signal_5447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5212 ( .a ({signal_8362, signal_5076}), .b ({signal_8559, signal_5267}), .c ({signal_8732, signal_5448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5213 ( .a ({signal_8557, signal_5265}), .b ({signal_8631, signal_5349}), .c ({signal_8733, signal_5449}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5214 ( .a ({signal_8629, signal_5347}), .b ({signal_8632, signal_5350}), .c ({signal_8734, signal_5450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5215 ( .a ({signal_8361, signal_5075}), .b ({signal_8633, signal_5351}), .c ({signal_8735, signal_5451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5216 ( .a ({signal_8366, signal_5080}), .b ({signal_8561, signal_5269}), .c ({signal_8736, signal_5452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5217 ( .a ({signal_8368, signal_5082}), .b ({signal_8562, signal_5270}), .c ({signal_8737, signal_5453}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5218 ( .a ({signal_8560, signal_5268}), .b ({signal_8637, signal_5355}), .c ({signal_8738, signal_5454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5219 ( .a ({signal_8635, signal_5353}), .b ({signal_8638, signal_5356}), .c ({signal_8739, signal_5455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5220 ( .a ({signal_8367, signal_5081}), .b ({signal_8639, signal_5357}), .c ({signal_8740, signal_5456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5221 ( .a ({signal_8671, signal_5359}), .b ({signal_8672, signal_5360}), .c ({signal_8765, signal_5457}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5222 ( .a ({signal_8523, signal_5207}), .b ({signal_8673, signal_5361}), .c ({signal_8766, signal_5458}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5223 ( .a ({signal_8672, signal_5360}), .b ({signal_8674, signal_5362}), .c ({signal_8767, signal_5459}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5224 ( .a ({signal_8523, signal_5207}), .b ({signal_8675, signal_5363}), .c ({signal_8768, signal_5460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5225 ( .a ({signal_8641, signal_5364}), .b ({signal_8642, signal_5365}), .c ({signal_8741, signal_5461}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5226 ( .a ({signal_8478, signal_5213}), .b ({signal_8643, signal_5366}), .c ({signal_8742, signal_5462}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5227 ( .a ({signal_8642, signal_5365}), .b ({signal_8644, signal_5367}), .c ({signal_8743, signal_5463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5228 ( .a ({signal_8478, signal_5213}), .b ({signal_8645, signal_5368}), .c ({signal_8744, signal_5464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5229 ( .a ({signal_8646, signal_5369}), .b ({signal_8647, signal_5370}), .c ({signal_8745, signal_5465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5230 ( .a ({signal_8484, signal_5219}), .b ({signal_8648, signal_5371}), .c ({signal_8746, signal_5466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5231 ( .a ({signal_8647, signal_5370}), .b ({signal_8649, signal_5372}), .c ({signal_8747, signal_5467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5232 ( .a ({signal_8484, signal_5219}), .b ({signal_8650, signal_5373}), .c ({signal_8748, signal_5468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5233 ( .a ({signal_8651, signal_5374}), .b ({signal_8652, signal_5375}), .c ({signal_8749, signal_5469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5234 ( .a ({signal_8490, signal_5225}), .b ({signal_8653, signal_5376}), .c ({signal_8750, signal_5470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5235 ( .a ({signal_8652, signal_5375}), .b ({signal_8654, signal_5377}), .c ({signal_8751, signal_5471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5236 ( .a ({signal_8490, signal_5225}), .b ({signal_8655, signal_5378}), .c ({signal_8752, signal_5472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5237 ( .a ({signal_8656, signal_5379}), .b ({signal_8657, signal_5380}), .c ({signal_8753, signal_5473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5238 ( .a ({signal_8496, signal_5231}), .b ({signal_8658, signal_5381}), .c ({signal_8754, signal_5474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5239 ( .a ({signal_8657, signal_5380}), .b ({signal_8659, signal_5382}), .c ({signal_8755, signal_5475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5240 ( .a ({signal_8496, signal_5231}), .b ({signal_8660, signal_5383}), .c ({signal_8756, signal_5476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5255 ( .a ({signal_8676, signal_5384}), .b ({signal_8677, signal_5385}), .c ({signal_8777, signal_5491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5256 ( .a ({signal_8568, signal_5276}), .b ({signal_8678, signal_5386}), .c ({signal_8778, signal_5492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5257 ( .a ({signal_8677, signal_5385}), .b ({signal_8679, signal_5387}), .c ({signal_8779, signal_5493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5258 ( .a ({signal_8568, signal_5276}), .b ({signal_8680, signal_5388}), .c ({signal_8780, signal_5494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5259 ( .a ({signal_8681, signal_5389}), .b ({signal_8682, signal_5390}), .c ({signal_8781, signal_5495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5260 ( .a ({signal_8574, signal_5282}), .b ({signal_8683, signal_5391}), .c ({signal_8782, signal_5496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5261 ( .a ({signal_8682, signal_5390}), .b ({signal_8684, signal_5392}), .c ({signal_8783, signal_5497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5262 ( .a ({signal_8574, signal_5282}), .b ({signal_8685, signal_5393}), .c ({signal_8784, signal_5498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5263 ( .a ({signal_8686, signal_5394}), .b ({signal_8687, signal_5395}), .c ({signal_8785, signal_5499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5264 ( .a ({signal_8580, signal_5288}), .b ({signal_8688, signal_5396}), .c ({signal_8786, signal_5500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5265 ( .a ({signal_8687, signal_5395}), .b ({signal_8689, signal_5397}), .c ({signal_8787, signal_5501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5266 ( .a ({signal_8580, signal_5288}), .b ({signal_8690, signal_5398}), .c ({signal_8788, signal_5502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5267 ( .a ({signal_8691, signal_5399}), .b ({signal_8692, signal_5400}), .c ({signal_8789, signal_5503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5268 ( .a ({signal_8586, signal_5294}), .b ({signal_8693, signal_5401}), .c ({signal_8790, signal_5504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5269 ( .a ({signal_8692, signal_5400}), .b ({signal_8694, signal_5402}), .c ({signal_8791, signal_5505}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5270 ( .a ({signal_8586, signal_5294}), .b ({signal_8695, signal_5403}), .c ({signal_8792, signal_5506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5271 ( .a ({signal_8696, signal_5404}), .b ({signal_8697, signal_5405}), .c ({signal_8793, signal_5507}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5272 ( .a ({signal_8592, signal_5300}), .b ({signal_8698, signal_5406}), .c ({signal_8794, signal_5508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5273 ( .a ({signal_8697, signal_5405}), .b ({signal_8699, signal_5407}), .c ({signal_8795, signal_5509}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5274 ( .a ({signal_8592, signal_5300}), .b ({signal_8700, signal_5408}), .c ({signal_8796, signal_5510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5275 ( .a ({signal_8701, signal_5409}), .b ({signal_8702, signal_5410}), .c ({signal_8797, signal_5511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5276 ( .a ({signal_8598, signal_5306}), .b ({signal_8703, signal_5411}), .c ({signal_8798, signal_5512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5277 ( .a ({signal_8702, signal_5410}), .b ({signal_8704, signal_5412}), .c ({signal_8799, signal_5513}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5278 ( .a ({signal_8598, signal_5306}), .b ({signal_8705, signal_5413}), .c ({signal_8800, signal_5514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5279 ( .a ({signal_8706, signal_5414}), .b ({signal_8707, signal_5415}), .c ({signal_8801, signal_5515}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5280 ( .a ({signal_8604, signal_5312}), .b ({signal_8708, signal_5416}), .c ({signal_8802, signal_5516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5281 ( .a ({signal_8707, signal_5415}), .b ({signal_8709, signal_5417}), .c ({signal_8803, signal_5517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5282 ( .a ({signal_8604, signal_5312}), .b ({signal_8710, signal_5418}), .c ({signal_8804, signal_5518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5283 ( .a ({signal_8507, signal_5149}), .b ({signal_8757, signal_5419}), .c ({signal_8843, signal_5519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5284 ( .a ({signal_8758, signal_5420}), .b ({signal_8759, signal_5421}), .c ({signal_8844, signal_5520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5285 ( .a ({signal_8711, signal_5423}), .b ({signal_8712, signal_5424}), .c ({signal_8805, signal_5521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5286 ( .a ({signal_8610, signal_5323}), .b ({signal_8713, signal_5425}), .c ({signal_8806, signal_5522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5287 ( .a ({signal_8712, signal_5424}), .b ({signal_8714, signal_5426}), .c ({signal_8807, signal_5523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5288 ( .a ({signal_8610, signal_5323}), .b ({signal_8715, signal_5427}), .c ({signal_8808, signal_5524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5289 ( .a ({signal_8716, signal_5428}), .b ({signal_8717, signal_5429}), .c ({signal_8809, signal_5525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5290 ( .a ({signal_8616, signal_5329}), .b ({signal_8718, signal_5430}), .c ({signal_8810, signal_5526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5291 ( .a ({signal_8717, signal_5429}), .b ({signal_8719, signal_5431}), .c ({signal_8811, signal_5527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5292 ( .a ({signal_8616, signal_5329}), .b ({signal_8720, signal_5432}), .c ({signal_8812, signal_5528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5293 ( .a ({signal_8721, signal_5433}), .b ({signal_8722, signal_5434}), .c ({signal_8813, signal_5529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5294 ( .a ({signal_8622, signal_5335}), .b ({signal_8723, signal_5435}), .c ({signal_8814, signal_5530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5295 ( .a ({signal_8722, signal_5434}), .b ({signal_8724, signal_5436}), .c ({signal_8815, signal_5531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5296 ( .a ({signal_8622, signal_5335}), .b ({signal_8725, signal_5437}), .c ({signal_8816, signal_5532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5297 ( .a ({signal_8513, signal_5176}), .b ({signal_8761, signal_5438}), .c ({signal_8845, signal_5533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5298 ( .a ({signal_8762, signal_5439}), .b ({signal_8763, signal_5440}), .c ({signal_8846, signal_5534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5299 ( .a ({signal_8726, signal_5442}), .b ({signal_8727, signal_5443}), .c ({signal_8817, signal_5535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5300 ( .a ({signal_8628, signal_5346}), .b ({signal_8728, signal_5444}), .c ({signal_8818, signal_5536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5301 ( .a ({signal_8727, signal_5443}), .b ({signal_8729, signal_5445}), .c ({signal_8819, signal_5537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5302 ( .a ({signal_8628, signal_5346}), .b ({signal_8730, signal_5446}), .c ({signal_8820, signal_5538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5303 ( .a ({signal_8731, signal_5447}), .b ({signal_8732, signal_5448}), .c ({signal_8821, signal_5539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5304 ( .a ({signal_8634, signal_5352}), .b ({signal_8733, signal_5449}), .c ({signal_8822, signal_5540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5305 ( .a ({signal_8732, signal_5448}), .b ({signal_8734, signal_5450}), .c ({signal_8823, signal_5541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5306 ( .a ({signal_8634, signal_5352}), .b ({signal_8735, signal_5451}), .c ({signal_8824, signal_5542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5307 ( .a ({signal_8736, signal_5452}), .b ({signal_8737, signal_5453}), .c ({signal_8825, signal_5543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5308 ( .a ({signal_8640, signal_5358}), .b ({signal_8738, signal_5454}), .c ({signal_8826, signal_5544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5309 ( .a ({signal_8737, signal_5453}), .b ({signal_8739, signal_5455}), .c ({signal_8827, signal_5545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5310 ( .a ({signal_8640, signal_5358}), .b ({signal_8740, signal_5456}), .c ({signal_8828, signal_5546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5311 ( .a ({signal_8519, signal_5203}), .b ({signal_8765, signal_5457}), .c ({signal_8847, signal_5547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5312 ( .a ({signal_8766, signal_5458}), .b ({signal_8767, signal_5459}), .c ({signal_8848, signal_5548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5313 ( .a ({signal_8474, signal_5209}), .b ({signal_8741, signal_5461}), .c ({signal_8829, signal_5549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5314 ( .a ({signal_8742, signal_5462}), .b ({signal_8743, signal_5463}), .c ({signal_8830, signal_5550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5315 ( .a ({signal_8480, signal_5215}), .b ({signal_8745, signal_5465}), .c ({signal_8831, signal_5551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5316 ( .a ({signal_8746, signal_5466}), .b ({signal_8747, signal_5467}), .c ({signal_8832, signal_5552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5317 ( .a ({signal_8486, signal_5221}), .b ({signal_8749, signal_5469}), .c ({signal_8833, signal_5553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5318 ( .a ({signal_8750, signal_5470}), .b ({signal_8751, signal_5471}), .c ({signal_8834, signal_5554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5319 ( .a ({signal_8492, signal_5227}), .b ({signal_8753, signal_5473}), .c ({signal_8835, signal_5555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5320 ( .a ({signal_8754, signal_5474}), .b ({signal_8755, signal_5475}), .c ({signal_8836, signal_5556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5354 ( .a ({signal_8564, signal_5272}), .b ({signal_8777, signal_5491}), .c ({signal_8879, signal_5590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5355 ( .a ({signal_8778, signal_5492}), .b ({signal_8779, signal_5493}), .c ({signal_8880, signal_5591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5356 ( .a ({signal_8570, signal_5278}), .b ({signal_8781, signal_5495}), .c ({signal_8881, signal_5592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5357 ( .a ({signal_8782, signal_5496}), .b ({signal_8783, signal_5497}), .c ({signal_8882, signal_5593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5358 ( .a ({signal_8576, signal_5284}), .b ({signal_8785, signal_5499}), .c ({signal_8883, signal_5594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5359 ( .a ({signal_8786, signal_5500}), .b ({signal_8787, signal_5501}), .c ({signal_8884, signal_5595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5360 ( .a ({signal_8582, signal_5290}), .b ({signal_8789, signal_5503}), .c ({signal_8885, signal_5596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5361 ( .a ({signal_8790, signal_5504}), .b ({signal_8791, signal_5505}), .c ({signal_8886, signal_5597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5362 ( .a ({signal_8588, signal_5296}), .b ({signal_8793, signal_5507}), .c ({signal_8887, signal_5598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5363 ( .a ({signal_8794, signal_5508}), .b ({signal_8795, signal_5509}), .c ({signal_8888, signal_5599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5364 ( .a ({signal_8594, signal_5302}), .b ({signal_8797, signal_5511}), .c ({signal_8889, signal_5600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5365 ( .a ({signal_8798, signal_5512}), .b ({signal_8799, signal_5513}), .c ({signal_8890, signal_5601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5366 ( .a ({signal_8600, signal_5308}), .b ({signal_8801, signal_5515}), .c ({signal_8891, signal_5602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5367 ( .a ({signal_8802, signal_5516}), .b ({signal_8803, signal_5517}), .c ({signal_8892, signal_5603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5368 ( .a ({signal_8760, signal_5422}), .b ({signal_8843, signal_5519}), .c ({signal_8924, signal_5604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5372 ( .a ({signal_8606, signal_5319}), .b ({signal_8805, signal_5521}), .c ({signal_8893, signal_5608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5373 ( .a ({signal_8806, signal_5522}), .b ({signal_8807, signal_5523}), .c ({signal_8894, signal_5609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5374 ( .a ({signal_8612, signal_5325}), .b ({signal_8809, signal_5525}), .c ({signal_8895, signal_5610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5375 ( .a ({signal_8810, signal_5526}), .b ({signal_8811, signal_5527}), .c ({signal_8896, signal_5611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5376 ( .a ({signal_8618, signal_5331}), .b ({signal_8813, signal_5529}), .c ({signal_8897, signal_5612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5377 ( .a ({signal_8814, signal_5530}), .b ({signal_8815, signal_5531}), .c ({signal_8898, signal_5613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5378 ( .a ({signal_8764, signal_5441}), .b ({signal_8845, signal_5533}), .c ({signal_8928, signal_5614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5382 ( .a ({signal_8624, signal_5342}), .b ({signal_8817, signal_5535}), .c ({signal_8899, signal_5618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5383 ( .a ({signal_8818, signal_5536}), .b ({signal_8819, signal_5537}), .c ({signal_8900, signal_5619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5384 ( .a ({signal_8630, signal_5348}), .b ({signal_8821, signal_5539}), .c ({signal_8901, signal_5620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5385 ( .a ({signal_8822, signal_5540}), .b ({signal_8823, signal_5541}), .c ({signal_8902, signal_5621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5386 ( .a ({signal_8636, signal_5354}), .b ({signal_8825, signal_5543}), .c ({signal_8903, signal_5622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5387 ( .a ({signal_8826, signal_5544}), .b ({signal_8827, signal_5545}), .c ({signal_8904, signal_5623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5388 ( .a ({signal_8768, signal_5460}), .b ({signal_8847, signal_5547}), .c ({signal_8932, signal_5624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5392 ( .a ({signal_8744, signal_5464}), .b ({signal_8829, signal_5549}), .c ({signal_8905, signal_5628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5396 ( .a ({signal_8748, signal_5468}), .b ({signal_8831, signal_5551}), .c ({signal_8909, signal_5632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5400 ( .a ({signal_8752, signal_5472}), .b ({signal_8833, signal_5553}), .c ({signal_8913, signal_5636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5404 ( .a ({signal_8756, signal_5476}), .b ({signal_8835, signal_5555}), .c ({signal_8917, signal_5640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5449 ( .a ({signal_8780, signal_5494}), .b ({signal_8879, signal_5590}), .c ({signal_8965, signal_5685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5453 ( .a ({signal_8784, signal_5498}), .b ({signal_8881, signal_5592}), .c ({signal_8969, signal_5689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5457 ( .a ({signal_8788, signal_5502}), .b ({signal_8883, signal_5594}), .c ({signal_8973, signal_5693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5461 ( .a ({signal_8792, signal_5506}), .b ({signal_8885, signal_5596}), .c ({signal_8977, signal_5697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5465 ( .a ({signal_8796, signal_5510}), .b ({signal_8887, signal_5598}), .c ({signal_8981, signal_5701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5469 ( .a ({signal_8800, signal_5514}), .b ({signal_8889, signal_5600}), .c ({signal_8985, signal_5705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5473 ( .a ({signal_8804, signal_5518}), .b ({signal_8891, signal_5602}), .c ({signal_8989, signal_5709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5478 ( .a ({signal_8808, signal_5524}), .b ({signal_8893, signal_5608}), .c ({signal_8993, signal_5714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5482 ( .a ({signal_8812, signal_5528}), .b ({signal_8895, signal_5610}), .c ({signal_8997, signal_5718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5486 ( .a ({signal_8816, signal_5532}), .b ({signal_8897, signal_5612}), .c ({signal_9001, signal_5722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5491 ( .a ({signal_8820, signal_5538}), .b ({signal_8899, signal_5618}), .c ({signal_9005, signal_5727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5495 ( .a ({signal_8824, signal_5542}), .b ({signal_8901, signal_5620}), .c ({signal_9009, signal_5731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5499 ( .a ({signal_8828, signal_5546}), .b ({signal_8903, signal_5622}), .c ({signal_9013, signal_5735}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5241 ( .a ({signal_8758, signal_5420}), .b ({signal_8760, signal_5422}), .clk (clk), .r (Fresh[180]), .c ({signal_8837, signal_5477}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5242 ( .a ({signal_8759, signal_5421}), .b ({signal_8760, signal_5422}), .clk (clk), .r (Fresh[181]), .c ({signal_8838, signal_5478}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5243 ( .a ({signal_8762, signal_5439}), .b ({signal_8764, signal_5441}), .clk (clk), .r (Fresh[182]), .c ({signal_8839, signal_5479}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5244 ( .a ({signal_8763, signal_5440}), .b ({signal_8764, signal_5441}), .clk (clk), .r (Fresh[183]), .c ({signal_8840, signal_5480}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5245 ( .a ({signal_8766, signal_5458}), .b ({signal_8768, signal_5460}), .clk (clk), .r (Fresh[184]), .c ({signal_8841, signal_5481}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5246 ( .a ({signal_8767, signal_5459}), .b ({signal_8768, signal_5460}), .clk (clk), .r (Fresh[185]), .c ({signal_8842, signal_5482}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5247 ( .a ({signal_8742, signal_5462}), .b ({signal_8744, signal_5464}), .clk (clk), .r (Fresh[186]), .c ({signal_8769, signal_5483}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5248 ( .a ({signal_8743, signal_5463}), .b ({signal_8744, signal_5464}), .clk (clk), .r (Fresh[187]), .c ({signal_8770, signal_5484}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5249 ( .a ({signal_8746, signal_5466}), .b ({signal_8748, signal_5468}), .clk (clk), .r (Fresh[188]), .c ({signal_8771, signal_5485}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5250 ( .a ({signal_8747, signal_5467}), .b ({signal_8748, signal_5468}), .clk (clk), .r (Fresh[189]), .c ({signal_8772, signal_5486}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5251 ( .a ({signal_8750, signal_5470}), .b ({signal_8752, signal_5472}), .clk (clk), .r (Fresh[190]), .c ({signal_8773, signal_5487}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5252 ( .a ({signal_8751, signal_5471}), .b ({signal_8752, signal_5472}), .clk (clk), .r (Fresh[191]), .c ({signal_8774, signal_5488}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5253 ( .a ({signal_8754, signal_5474}), .b ({signal_8756, signal_5476}), .clk (clk), .r (Fresh[192]), .c ({signal_8775, signal_5489}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5254 ( .a ({signal_8755, signal_5475}), .b ({signal_8756, signal_5476}), .clk (clk), .r (Fresh[193]), .c ({signal_8776, signal_5490}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5321 ( .a ({signal_8778, signal_5492}), .b ({signal_8780, signal_5494}), .clk (clk), .r (Fresh[194]), .c ({signal_8849, signal_5557}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5322 ( .a ({signal_8779, signal_5493}), .b ({signal_8780, signal_5494}), .clk (clk), .r (Fresh[195]), .c ({signal_8850, signal_5558}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5323 ( .a ({signal_8782, signal_5496}), .b ({signal_8784, signal_5498}), .clk (clk), .r (Fresh[196]), .c ({signal_8851, signal_5559}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5324 ( .a ({signal_8783, signal_5497}), .b ({signal_8784, signal_5498}), .clk (clk), .r (Fresh[197]), .c ({signal_8852, signal_5560}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5325 ( .a ({signal_8786, signal_5500}), .b ({signal_8788, signal_5502}), .clk (clk), .r (Fresh[198]), .c ({signal_8853, signal_5561}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5326 ( .a ({signal_8787, signal_5501}), .b ({signal_8788, signal_5502}), .clk (clk), .r (Fresh[199]), .c ({signal_8854, signal_5562}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5327 ( .a ({signal_8790, signal_5504}), .b ({signal_8792, signal_5506}), .clk (clk), .r (Fresh[200]), .c ({signal_8855, signal_5563}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5328 ( .a ({signal_8791, signal_5505}), .b ({signal_8792, signal_5506}), .clk (clk), .r (Fresh[201]), .c ({signal_8856, signal_5564}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5329 ( .a ({signal_8794, signal_5508}), .b ({signal_8796, signal_5510}), .clk (clk), .r (Fresh[202]), .c ({signal_8857, signal_5565}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5330 ( .a ({signal_8795, signal_5509}), .b ({signal_8796, signal_5510}), .clk (clk), .r (Fresh[203]), .c ({signal_8858, signal_5566}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5331 ( .a ({signal_8798, signal_5512}), .b ({signal_8800, signal_5514}), .clk (clk), .r (Fresh[204]), .c ({signal_8859, signal_5567}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5332 ( .a ({signal_8799, signal_5513}), .b ({signal_8800, signal_5514}), .clk (clk), .r (Fresh[205]), .c ({signal_8860, signal_5568}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5333 ( .a ({signal_8802, signal_5516}), .b ({signal_8804, signal_5518}), .clk (clk), .r (Fresh[206]), .c ({signal_8861, signal_5569}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5334 ( .a ({signal_8803, signal_5517}), .b ({signal_8804, signal_5518}), .clk (clk), .r (Fresh[207]), .c ({signal_8862, signal_5570}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5335 ( .a ({signal_8758, signal_5420}), .b ({signal_8843, signal_5519}), .clk (clk), .r (Fresh[208]), .c ({signal_8921, signal_5571}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5336 ( .a ({signal_8806, signal_5522}), .b ({signal_8808, signal_5524}), .clk (clk), .r (Fresh[209]), .c ({signal_8863, signal_5572}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5337 ( .a ({signal_8807, signal_5523}), .b ({signal_8808, signal_5524}), .clk (clk), .r (Fresh[210]), .c ({signal_8864, signal_5573}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5338 ( .a ({signal_8810, signal_5526}), .b ({signal_8812, signal_5528}), .clk (clk), .r (Fresh[211]), .c ({signal_8865, signal_5574}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5339 ( .a ({signal_8811, signal_5527}), .b ({signal_8812, signal_5528}), .clk (clk), .r (Fresh[212]), .c ({signal_8866, signal_5575}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5340 ( .a ({signal_8814, signal_5530}), .b ({signal_8816, signal_5532}), .clk (clk), .r (Fresh[213]), .c ({signal_8867, signal_5576}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5341 ( .a ({signal_8815, signal_5531}), .b ({signal_8816, signal_5532}), .clk (clk), .r (Fresh[214]), .c ({signal_8868, signal_5577}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5342 ( .a ({signal_8762, signal_5439}), .b ({signal_8845, signal_5533}), .clk (clk), .r (Fresh[215]), .c ({signal_8922, signal_5578}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5343 ( .a ({signal_8818, signal_5536}), .b ({signal_8820, signal_5538}), .clk (clk), .r (Fresh[216]), .c ({signal_8869, signal_5579}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5344 ( .a ({signal_8819, signal_5537}), .b ({signal_8820, signal_5538}), .clk (clk), .r (Fresh[217]), .c ({signal_8870, signal_5580}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5345 ( .a ({signal_8822, signal_5540}), .b ({signal_8824, signal_5542}), .clk (clk), .r (Fresh[218]), .c ({signal_8871, signal_5581}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5346 ( .a ({signal_8823, signal_5541}), .b ({signal_8824, signal_5542}), .clk (clk), .r (Fresh[219]), .c ({signal_8872, signal_5582}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5347 ( .a ({signal_8826, signal_5544}), .b ({signal_8828, signal_5546}), .clk (clk), .r (Fresh[220]), .c ({signal_8873, signal_5583}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5348 ( .a ({signal_8827, signal_5545}), .b ({signal_8828, signal_5546}), .clk (clk), .r (Fresh[221]), .c ({signal_8874, signal_5584}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5349 ( .a ({signal_8766, signal_5458}), .b ({signal_8847, signal_5547}), .clk (clk), .r (Fresh[222]), .c ({signal_8923, signal_5585}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5350 ( .a ({signal_8742, signal_5462}), .b ({signal_8829, signal_5549}), .clk (clk), .r (Fresh[223]), .c ({signal_8875, signal_5586}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5351 ( .a ({signal_8746, signal_5466}), .b ({signal_8831, signal_5551}), .clk (clk), .r (Fresh[224]), .c ({signal_8876, signal_5587}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5352 ( .a ({signal_8750, signal_5470}), .b ({signal_8833, signal_5553}), .clk (clk), .r (Fresh[225]), .c ({signal_8877, signal_5588}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5353 ( .a ({signal_8754, signal_5474}), .b ({signal_8835, signal_5555}), .clk (clk), .r (Fresh[226]), .c ({signal_8878, signal_5589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5369 ( .a ({signal_8759, signal_5421}), .b ({signal_8837, signal_5477}), .c ({signal_8925, signal_5605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5370 ( .a ({signal_8843, signal_5519}), .b ({signal_8837, signal_5477}), .c ({signal_8926, signal_5606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5371 ( .a ({signal_8837, signal_5477}), .b ({signal_8844, signal_5520}), .c ({signal_8927, signal_5607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5379 ( .a ({signal_8763, signal_5440}), .b ({signal_8839, signal_5479}), .c ({signal_8929, signal_5615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5380 ( .a ({signal_8845, signal_5533}), .b ({signal_8839, signal_5479}), .c ({signal_8930, signal_5616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5381 ( .a ({signal_8839, signal_5479}), .b ({signal_8846, signal_5534}), .c ({signal_8931, signal_5617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5389 ( .a ({signal_8767, signal_5459}), .b ({signal_8841, signal_5481}), .c ({signal_8933, signal_5625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5390 ( .a ({signal_8847, signal_5547}), .b ({signal_8841, signal_5481}), .c ({signal_8934, signal_5626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5391 ( .a ({signal_8841, signal_5481}), .b ({signal_8848, signal_5548}), .c ({signal_8935, signal_5627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5393 ( .a ({signal_8743, signal_5463}), .b ({signal_8769, signal_5483}), .c ({signal_8906, signal_5629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5394 ( .a ({signal_8829, signal_5549}), .b ({signal_8769, signal_5483}), .c ({signal_8907, signal_5630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5395 ( .a ({signal_8769, signal_5483}), .b ({signal_8830, signal_5550}), .c ({signal_8908, signal_5631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5397 ( .a ({signal_8747, signal_5467}), .b ({signal_8771, signal_5485}), .c ({signal_8910, signal_5633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5398 ( .a ({signal_8831, signal_5551}), .b ({signal_8771, signal_5485}), .c ({signal_8911, signal_5634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5399 ( .a ({signal_8771, signal_5485}), .b ({signal_8832, signal_5552}), .c ({signal_8912, signal_5635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5401 ( .a ({signal_8751, signal_5471}), .b ({signal_8773, signal_5487}), .c ({signal_8914, signal_5637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5402 ( .a ({signal_8833, signal_5553}), .b ({signal_8773, signal_5487}), .c ({signal_8915, signal_5638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5403 ( .a ({signal_8773, signal_5487}), .b ({signal_8834, signal_5554}), .c ({signal_8916, signal_5639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5405 ( .a ({signal_8755, signal_5475}), .b ({signal_8775, signal_5489}), .c ({signal_8918, signal_5641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5406 ( .a ({signal_8835, signal_5555}), .b ({signal_8775, signal_5489}), .c ({signal_8919, signal_5642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5407 ( .a ({signal_8775, signal_5489}), .b ({signal_8836, signal_5556}), .c ({signal_8920, signal_5643}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5408 ( .a ({signal_8778, signal_5492}), .b ({signal_8879, signal_5590}), .clk (clk), .r (Fresh[227]), .c ({signal_8936, signal_5644}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5409 ( .a ({signal_8782, signal_5496}), .b ({signal_8881, signal_5592}), .clk (clk), .r (Fresh[228]), .c ({signal_8937, signal_5645}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5410 ( .a ({signal_8786, signal_5500}), .b ({signal_8883, signal_5594}), .clk (clk), .r (Fresh[229]), .c ({signal_8938, signal_5646}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5411 ( .a ({signal_8790, signal_5504}), .b ({signal_8885, signal_5596}), .clk (clk), .r (Fresh[230]), .c ({signal_8939, signal_5647}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5412 ( .a ({signal_8794, signal_5508}), .b ({signal_8887, signal_5598}), .clk (clk), .r (Fresh[231]), .c ({signal_8940, signal_5648}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5413 ( .a ({signal_8798, signal_5512}), .b ({signal_8889, signal_5600}), .clk (clk), .r (Fresh[232]), .c ({signal_8941, signal_5649}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5414 ( .a ({signal_8802, signal_5516}), .b ({signal_8891, signal_5602}), .clk (clk), .r (Fresh[233]), .c ({signal_8942, signal_5650}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5419 ( .a ({signal_8806, signal_5522}), .b ({signal_8893, signal_5608}), .clk (clk), .r (Fresh[234]), .c ({signal_8943, signal_5655}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5420 ( .a ({signal_8810, signal_5526}), .b ({signal_8895, signal_5610}), .clk (clk), .r (Fresh[235]), .c ({signal_8944, signal_5656}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5421 ( .a ({signal_8814, signal_5530}), .b ({signal_8897, signal_5612}), .clk (clk), .r (Fresh[236]), .c ({signal_8945, signal_5657}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5426 ( .a ({signal_8818, signal_5536}), .b ({signal_8899, signal_5618}), .clk (clk), .r (Fresh[237]), .c ({signal_8946, signal_5662}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5427 ( .a ({signal_8822, signal_5540}), .b ({signal_8901, signal_5620}), .clk (clk), .r (Fresh[238]), .c ({signal_8947, signal_5663}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5428 ( .a ({signal_8826, signal_5544}), .b ({signal_8903, signal_5622}), .clk (clk), .r (Fresh[239]), .c ({signal_8948, signal_5664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5450 ( .a ({signal_8779, signal_5493}), .b ({signal_8849, signal_5557}), .c ({signal_8966, signal_5686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5451 ( .a ({signal_8879, signal_5590}), .b ({signal_8849, signal_5557}), .c ({signal_8967, signal_5687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5452 ( .a ({signal_8849, signal_5557}), .b ({signal_8880, signal_5591}), .c ({signal_8968, signal_5688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5454 ( .a ({signal_8783, signal_5497}), .b ({signal_8851, signal_5559}), .c ({signal_8970, signal_5690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5455 ( .a ({signal_8881, signal_5592}), .b ({signal_8851, signal_5559}), .c ({signal_8971, signal_5691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5456 ( .a ({signal_8851, signal_5559}), .b ({signal_8882, signal_5593}), .c ({signal_8972, signal_5692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5458 ( .a ({signal_8787, signal_5501}), .b ({signal_8853, signal_5561}), .c ({signal_8974, signal_5694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5459 ( .a ({signal_8883, signal_5594}), .b ({signal_8853, signal_5561}), .c ({signal_8975, signal_5695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5460 ( .a ({signal_8853, signal_5561}), .b ({signal_8884, signal_5595}), .c ({signal_8976, signal_5696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5462 ( .a ({signal_8791, signal_5505}), .b ({signal_8855, signal_5563}), .c ({signal_8978, signal_5698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5463 ( .a ({signal_8885, signal_5596}), .b ({signal_8855, signal_5563}), .c ({signal_8979, signal_5699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5464 ( .a ({signal_8855, signal_5563}), .b ({signal_8886, signal_5597}), .c ({signal_8980, signal_5700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5466 ( .a ({signal_8795, signal_5509}), .b ({signal_8857, signal_5565}), .c ({signal_8982, signal_5702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5467 ( .a ({signal_8887, signal_5598}), .b ({signal_8857, signal_5565}), .c ({signal_8983, signal_5703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5468 ( .a ({signal_8857, signal_5565}), .b ({signal_8888, signal_5599}), .c ({signal_8984, signal_5704}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5470 ( .a ({signal_8799, signal_5513}), .b ({signal_8859, signal_5567}), .c ({signal_8986, signal_5706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5471 ( .a ({signal_8889, signal_5600}), .b ({signal_8859, signal_5567}), .c ({signal_8987, signal_5707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5472 ( .a ({signal_8859, signal_5567}), .b ({signal_8890, signal_5601}), .c ({signal_8988, signal_5708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5474 ( .a ({signal_8803, signal_5517}), .b ({signal_8861, signal_5569}), .c ({signal_8990, signal_5710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5475 ( .a ({signal_8891, signal_5602}), .b ({signal_8861, signal_5569}), .c ({signal_8991, signal_5711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5476 ( .a ({signal_8861, signal_5569}), .b ({signal_8892, signal_5603}), .c ({signal_8992, signal_5712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5477 ( .a ({signal_8837, signal_5477}), .b ({signal_8924, signal_5604}), .c ({signal_9033, signal_5713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5479 ( .a ({signal_8807, signal_5523}), .b ({signal_8863, signal_5572}), .c ({signal_8994, signal_5715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5480 ( .a ({signal_8893, signal_5608}), .b ({signal_8863, signal_5572}), .c ({signal_8995, signal_5716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5481 ( .a ({signal_8863, signal_5572}), .b ({signal_8894, signal_5609}), .c ({signal_8996, signal_5717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5483 ( .a ({signal_8811, signal_5527}), .b ({signal_8865, signal_5574}), .c ({signal_8998, signal_5719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5484 ( .a ({signal_8895, signal_5610}), .b ({signal_8865, signal_5574}), .c ({signal_8999, signal_5720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5485 ( .a ({signal_8865, signal_5574}), .b ({signal_8896, signal_5611}), .c ({signal_9000, signal_5721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5487 ( .a ({signal_8815, signal_5531}), .b ({signal_8867, signal_5576}), .c ({signal_9002, signal_5723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5488 ( .a ({signal_8897, signal_5612}), .b ({signal_8867, signal_5576}), .c ({signal_9003, signal_5724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5489 ( .a ({signal_8867, signal_5576}), .b ({signal_8898, signal_5613}), .c ({signal_9004, signal_5725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5490 ( .a ({signal_8839, signal_5479}), .b ({signal_8928, signal_5614}), .c ({signal_9034, signal_5726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5492 ( .a ({signal_8819, signal_5537}), .b ({signal_8869, signal_5579}), .c ({signal_9006, signal_5728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5493 ( .a ({signal_8899, signal_5618}), .b ({signal_8869, signal_5579}), .c ({signal_9007, signal_5729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5494 ( .a ({signal_8869, signal_5579}), .b ({signal_8900, signal_5619}), .c ({signal_9008, signal_5730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5496 ( .a ({signal_8823, signal_5541}), .b ({signal_8871, signal_5581}), .c ({signal_9010, signal_5732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5497 ( .a ({signal_8901, signal_5620}), .b ({signal_8871, signal_5581}), .c ({signal_9011, signal_5733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5498 ( .a ({signal_8871, signal_5581}), .b ({signal_8902, signal_5621}), .c ({signal_9012, signal_5734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5500 ( .a ({signal_8827, signal_5545}), .b ({signal_8873, signal_5583}), .c ({signal_9014, signal_5736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5501 ( .a ({signal_8903, signal_5622}), .b ({signal_8873, signal_5583}), .c ({signal_9015, signal_5737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5502 ( .a ({signal_8873, signal_5583}), .b ({signal_8904, signal_5623}), .c ({signal_9016, signal_5738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5503 ( .a ({signal_8841, signal_5481}), .b ({signal_8932, signal_5624}), .c ({signal_9035, signal_5739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5504 ( .a ({signal_8769, signal_5483}), .b ({signal_8905, signal_5628}), .c ({signal_9017, signal_5740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5505 ( .a ({signal_8771, signal_5485}), .b ({signal_8909, signal_5632}), .c ({signal_9018, signal_5741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5506 ( .a ({signal_8773, signal_5487}), .b ({signal_8913, signal_5636}), .c ({signal_9019, signal_5742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5507 ( .a ({signal_8775, signal_5489}), .b ({signal_8917, signal_5640}), .c ({signal_9020, signal_5743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5560 ( .a ({signal_8849, signal_5557}), .b ({signal_8965, signal_5685}), .c ({signal_9088, signal_5796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5561 ( .a ({signal_8851, signal_5559}), .b ({signal_8969, signal_5689}), .c ({signal_9089, signal_5797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5562 ( .a ({signal_8853, signal_5561}), .b ({signal_8973, signal_5693}), .c ({signal_9090, signal_5798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5563 ( .a ({signal_8855, signal_5563}), .b ({signal_8977, signal_5697}), .c ({signal_9091, signal_5799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5564 ( .a ({signal_8857, signal_5565}), .b ({signal_8981, signal_5701}), .c ({signal_9092, signal_5800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5565 ( .a ({signal_8859, signal_5567}), .b ({signal_8985, signal_5705}), .c ({signal_9093, signal_5801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5566 ( .a ({signal_8861, signal_5569}), .b ({signal_8989, signal_5709}), .c ({signal_9094, signal_5802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5571 ( .a ({signal_8863, signal_5572}), .b ({signal_8993, signal_5714}), .c ({signal_9095, signal_5807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5572 ( .a ({signal_8865, signal_5574}), .b ({signal_8997, signal_5718}), .c ({signal_9096, signal_5808}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5573 ( .a ({signal_8867, signal_5576}), .b ({signal_9001, signal_5722}), .c ({signal_9097, signal_5809}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5578 ( .a ({signal_8869, signal_5579}), .b ({signal_9005, signal_5727}), .c ({signal_9098, signal_5814}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5579 ( .a ({signal_8871, signal_5581}), .b ({signal_9009, signal_5731}), .c ({signal_9099, signal_5815}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5580 ( .a ({signal_8873, signal_5583}), .b ({signal_9013, signal_5735}), .c ({signal_9100, signal_5816}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5415 ( .a ({signal_8844, signal_5520}), .b ({signal_8926, signal_5606}), .clk (clk), .r (Fresh[240]), .c ({signal_9021, signal_5651}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5416 ( .a ({signal_8924, signal_5604}), .b ({signal_8925, signal_5605}), .clk (clk), .r (Fresh[241]), .c ({signal_9022, signal_5652}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5417 ( .a ({signal_8844, signal_5520}), .b ({signal_8921, signal_5571}), .clk (clk), .r (Fresh[242]), .c ({signal_9023, signal_5653}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5418 ( .a ({signal_8838, signal_5478}), .b ({signal_8924, signal_5604}), .clk (clk), .r (Fresh[243]), .c ({signal_9024, signal_5654}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5422 ( .a ({signal_8846, signal_5534}), .b ({signal_8930, signal_5616}), .clk (clk), .r (Fresh[244]), .c ({signal_9025, signal_5658}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5423 ( .a ({signal_8928, signal_5614}), .b ({signal_8929, signal_5615}), .clk (clk), .r (Fresh[245]), .c ({signal_9026, signal_5659}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5424 ( .a ({signal_8846, signal_5534}), .b ({signal_8922, signal_5578}), .clk (clk), .r (Fresh[246]), .c ({signal_9027, signal_5660}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5425 ( .a ({signal_8840, signal_5480}), .b ({signal_8928, signal_5614}), .clk (clk), .r (Fresh[247]), .c ({signal_9028, signal_5661}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5429 ( .a ({signal_8848, signal_5548}), .b ({signal_8934, signal_5626}), .clk (clk), .r (Fresh[248]), .c ({signal_9029, signal_5665}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5430 ( .a ({signal_8932, signal_5624}), .b ({signal_8933, signal_5625}), .clk (clk), .r (Fresh[249]), .c ({signal_9030, signal_5666}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5431 ( .a ({signal_8848, signal_5548}), .b ({signal_8923, signal_5585}), .clk (clk), .r (Fresh[250]), .c ({signal_9031, signal_5667}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5432 ( .a ({signal_8842, signal_5482}), .b ({signal_8932, signal_5624}), .clk (clk), .r (Fresh[251]), .c ({signal_9032, signal_5668}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5433 ( .a ({signal_8830, signal_5550}), .b ({signal_8907, signal_5630}), .clk (clk), .r (Fresh[252]), .c ({signal_8949, signal_5669}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5434 ( .a ({signal_8905, signal_5628}), .b ({signal_8906, signal_5629}), .clk (clk), .r (Fresh[253]), .c ({signal_8950, signal_5670}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5435 ( .a ({signal_8830, signal_5550}), .b ({signal_8875, signal_5586}), .clk (clk), .r (Fresh[254]), .c ({signal_8951, signal_5671}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5436 ( .a ({signal_8770, signal_5484}), .b ({signal_8905, signal_5628}), .clk (clk), .r (Fresh[255]), .c ({signal_8952, signal_5672}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5437 ( .a ({signal_8832, signal_5552}), .b ({signal_8911, signal_5634}), .clk (clk), .r (Fresh[256]), .c ({signal_8953, signal_5673}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5438 ( .a ({signal_8909, signal_5632}), .b ({signal_8910, signal_5633}), .clk (clk), .r (Fresh[257]), .c ({signal_8954, signal_5674}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5439 ( .a ({signal_8832, signal_5552}), .b ({signal_8876, signal_5587}), .clk (clk), .r (Fresh[258]), .c ({signal_8955, signal_5675}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5440 ( .a ({signal_8772, signal_5486}), .b ({signal_8909, signal_5632}), .clk (clk), .r (Fresh[259]), .c ({signal_8956, signal_5676}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5441 ( .a ({signal_8834, signal_5554}), .b ({signal_8915, signal_5638}), .clk (clk), .r (Fresh[260]), .c ({signal_8957, signal_5677}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5442 ( .a ({signal_8913, signal_5636}), .b ({signal_8914, signal_5637}), .clk (clk), .r (Fresh[261]), .c ({signal_8958, signal_5678}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5443 ( .a ({signal_8834, signal_5554}), .b ({signal_8877, signal_5588}), .clk (clk), .r (Fresh[262]), .c ({signal_8959, signal_5679}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5444 ( .a ({signal_8774, signal_5488}), .b ({signal_8913, signal_5636}), .clk (clk), .r (Fresh[263]), .c ({signal_8960, signal_5680}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5445 ( .a ({signal_8836, signal_5556}), .b ({signal_8919, signal_5642}), .clk (clk), .r (Fresh[264]), .c ({signal_8961, signal_5681}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5446 ( .a ({signal_8917, signal_5640}), .b ({signal_8918, signal_5641}), .clk (clk), .r (Fresh[265]), .c ({signal_8962, signal_5682}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5447 ( .a ({signal_8836, signal_5556}), .b ({signal_8878, signal_5589}), .clk (clk), .r (Fresh[266]), .c ({signal_8963, signal_5683}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5448 ( .a ({signal_8776, signal_5490}), .b ({signal_8917, signal_5640}), .clk (clk), .r (Fresh[267]), .c ({signal_8964, signal_5684}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5508 ( .a ({signal_8880, signal_5591}), .b ({signal_8967, signal_5687}), .clk (clk), .r (Fresh[268]), .c ({signal_9036, signal_5744}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5509 ( .a ({signal_8965, signal_5685}), .b ({signal_8966, signal_5686}), .clk (clk), .r (Fresh[269]), .c ({signal_9037, signal_5745}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5510 ( .a ({signal_8880, signal_5591}), .b ({signal_8936, signal_5644}), .clk (clk), .r (Fresh[270]), .c ({signal_9038, signal_5746}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5511 ( .a ({signal_8850, signal_5558}), .b ({signal_8965, signal_5685}), .clk (clk), .r (Fresh[271]), .c ({signal_9039, signal_5747}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5512 ( .a ({signal_8882, signal_5593}), .b ({signal_8971, signal_5691}), .clk (clk), .r (Fresh[272]), .c ({signal_9040, signal_5748}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5513 ( .a ({signal_8969, signal_5689}), .b ({signal_8970, signal_5690}), .clk (clk), .r (Fresh[273]), .c ({signal_9041, signal_5749}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5514 ( .a ({signal_8882, signal_5593}), .b ({signal_8937, signal_5645}), .clk (clk), .r (Fresh[274]), .c ({signal_9042, signal_5750}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5515 ( .a ({signal_8852, signal_5560}), .b ({signal_8969, signal_5689}), .clk (clk), .r (Fresh[275]), .c ({signal_9043, signal_5751}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5516 ( .a ({signal_8884, signal_5595}), .b ({signal_8975, signal_5695}), .clk (clk), .r (Fresh[276]), .c ({signal_9044, signal_5752}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5517 ( .a ({signal_8973, signal_5693}), .b ({signal_8974, signal_5694}), .clk (clk), .r (Fresh[277]), .c ({signal_9045, signal_5753}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5518 ( .a ({signal_8884, signal_5595}), .b ({signal_8938, signal_5646}), .clk (clk), .r (Fresh[278]), .c ({signal_9046, signal_5754}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5519 ( .a ({signal_8854, signal_5562}), .b ({signal_8973, signal_5693}), .clk (clk), .r (Fresh[279]), .c ({signal_9047, signal_5755}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5520 ( .a ({signal_8886, signal_5597}), .b ({signal_8979, signal_5699}), .clk (clk), .r (Fresh[280]), .c ({signal_9048, signal_5756}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5521 ( .a ({signal_8977, signal_5697}), .b ({signal_8978, signal_5698}), .clk (clk), .r (Fresh[281]), .c ({signal_9049, signal_5757}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5522 ( .a ({signal_8886, signal_5597}), .b ({signal_8939, signal_5647}), .clk (clk), .r (Fresh[282]), .c ({signal_9050, signal_5758}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5523 ( .a ({signal_8856, signal_5564}), .b ({signal_8977, signal_5697}), .clk (clk), .r (Fresh[283]), .c ({signal_9051, signal_5759}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5524 ( .a ({signal_8888, signal_5599}), .b ({signal_8983, signal_5703}), .clk (clk), .r (Fresh[284]), .c ({signal_9052, signal_5760}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5525 ( .a ({signal_8981, signal_5701}), .b ({signal_8982, signal_5702}), .clk (clk), .r (Fresh[285]), .c ({signal_9053, signal_5761}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5526 ( .a ({signal_8888, signal_5599}), .b ({signal_8940, signal_5648}), .clk (clk), .r (Fresh[286]), .c ({signal_9054, signal_5762}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5527 ( .a ({signal_8858, signal_5566}), .b ({signal_8981, signal_5701}), .clk (clk), .r (Fresh[287]), .c ({signal_9055, signal_5763}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5528 ( .a ({signal_8890, signal_5601}), .b ({signal_8987, signal_5707}), .clk (clk), .r (Fresh[288]), .c ({signal_9056, signal_5764}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5529 ( .a ({signal_8985, signal_5705}), .b ({signal_8986, signal_5706}), .clk (clk), .r (Fresh[289]), .c ({signal_9057, signal_5765}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5530 ( .a ({signal_8890, signal_5601}), .b ({signal_8941, signal_5649}), .clk (clk), .r (Fresh[290]), .c ({signal_9058, signal_5766}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5531 ( .a ({signal_8860, signal_5568}), .b ({signal_8985, signal_5705}), .clk (clk), .r (Fresh[291]), .c ({signal_9059, signal_5767}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5532 ( .a ({signal_8892, signal_5603}), .b ({signal_8991, signal_5711}), .clk (clk), .r (Fresh[292]), .c ({signal_9060, signal_5768}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5533 ( .a ({signal_8989, signal_5709}), .b ({signal_8990, signal_5710}), .clk (clk), .r (Fresh[293]), .c ({signal_9061, signal_5769}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5534 ( .a ({signal_8892, signal_5603}), .b ({signal_8942, signal_5650}), .clk (clk), .r (Fresh[294]), .c ({signal_9062, signal_5770}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5535 ( .a ({signal_8862, signal_5570}), .b ({signal_8989, signal_5709}), .clk (clk), .r (Fresh[295]), .c ({signal_9063, signal_5771}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5536 ( .a ({signal_8894, signal_5609}), .b ({signal_8995, signal_5716}), .clk (clk), .r (Fresh[296]), .c ({signal_9064, signal_5772}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5537 ( .a ({signal_8993, signal_5714}), .b ({signal_8994, signal_5715}), .clk (clk), .r (Fresh[297]), .c ({signal_9065, signal_5773}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5538 ( .a ({signal_8894, signal_5609}), .b ({signal_8943, signal_5655}), .clk (clk), .r (Fresh[298]), .c ({signal_9066, signal_5774}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5539 ( .a ({signal_8864, signal_5573}), .b ({signal_8993, signal_5714}), .clk (clk), .r (Fresh[299]), .c ({signal_9067, signal_5775}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5540 ( .a ({signal_8896, signal_5611}), .b ({signal_8999, signal_5720}), .clk (clk), .r (Fresh[300]), .c ({signal_9068, signal_5776}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5541 ( .a ({signal_8997, signal_5718}), .b ({signal_8998, signal_5719}), .clk (clk), .r (Fresh[301]), .c ({signal_9069, signal_5777}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5542 ( .a ({signal_8896, signal_5611}), .b ({signal_8944, signal_5656}), .clk (clk), .r (Fresh[302]), .c ({signal_9070, signal_5778}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5543 ( .a ({signal_8866, signal_5575}), .b ({signal_8997, signal_5718}), .clk (clk), .r (Fresh[303]), .c ({signal_9071, signal_5779}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5544 ( .a ({signal_8898, signal_5613}), .b ({signal_9003, signal_5724}), .clk (clk), .r (Fresh[304]), .c ({signal_9072, signal_5780}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5545 ( .a ({signal_9001, signal_5722}), .b ({signal_9002, signal_5723}), .clk (clk), .r (Fresh[305]), .c ({signal_9073, signal_5781}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5546 ( .a ({signal_8898, signal_5613}), .b ({signal_8945, signal_5657}), .clk (clk), .r (Fresh[306]), .c ({signal_9074, signal_5782}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5547 ( .a ({signal_8868, signal_5577}), .b ({signal_9001, signal_5722}), .clk (clk), .r (Fresh[307]), .c ({signal_9075, signal_5783}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5548 ( .a ({signal_8900, signal_5619}), .b ({signal_9007, signal_5729}), .clk (clk), .r (Fresh[308]), .c ({signal_9076, signal_5784}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5549 ( .a ({signal_9005, signal_5727}), .b ({signal_9006, signal_5728}), .clk (clk), .r (Fresh[309]), .c ({signal_9077, signal_5785}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5550 ( .a ({signal_8900, signal_5619}), .b ({signal_8946, signal_5662}), .clk (clk), .r (Fresh[310]), .c ({signal_9078, signal_5786}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5551 ( .a ({signal_8870, signal_5580}), .b ({signal_9005, signal_5727}), .clk (clk), .r (Fresh[311]), .c ({signal_9079, signal_5787}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5552 ( .a ({signal_8902, signal_5621}), .b ({signal_9011, signal_5733}), .clk (clk), .r (Fresh[312]), .c ({signal_9080, signal_5788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5553 ( .a ({signal_9009, signal_5731}), .b ({signal_9010, signal_5732}), .clk (clk), .r (Fresh[313]), .c ({signal_9081, signal_5789}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5554 ( .a ({signal_8902, signal_5621}), .b ({signal_8947, signal_5663}), .clk (clk), .r (Fresh[314]), .c ({signal_9082, signal_5790}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5555 ( .a ({signal_8872, signal_5582}), .b ({signal_9009, signal_5731}), .clk (clk), .r (Fresh[315]), .c ({signal_9083, signal_5791}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5556 ( .a ({signal_8904, signal_5623}), .b ({signal_9015, signal_5737}), .clk (clk), .r (Fresh[316]), .c ({signal_9084, signal_5792}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5557 ( .a ({signal_9013, signal_5735}), .b ({signal_9014, signal_5736}), .clk (clk), .r (Fresh[317]), .c ({signal_9085, signal_5793}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5558 ( .a ({signal_8904, signal_5623}), .b ({signal_8948, signal_5664}), .clk (clk), .r (Fresh[318]), .c ({signal_9086, signal_5794}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5559 ( .a ({signal_8874, signal_5584}), .b ({signal_9013, signal_5735}), .clk (clk), .r (Fresh[319]), .c ({signal_9087, signal_5795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5567 ( .a ({signal_8759, signal_5421}), .b ({signal_9021, signal_5651}), .c ({signal_9117, signal_5803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5568 ( .a ({signal_8927, signal_5607}), .b ({signal_9023, signal_5653}), .c ({signal_9118, signal_5804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5569 ( .a ({signal_8843, signal_5519}), .b ({signal_9022, signal_5652}), .c ({signal_9119, signal_5805}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5570 ( .a ({signal_9024, signal_5654}), .b ({signal_9033, signal_5713}), .c ({signal_9120, signal_5806}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5574 ( .a ({signal_8763, signal_5440}), .b ({signal_9025, signal_5658}), .c ({signal_9121, signal_5810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5575 ( .a ({signal_8931, signal_5617}), .b ({signal_9027, signal_5660}), .c ({signal_9122, signal_5811}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5576 ( .a ({signal_8845, signal_5533}), .b ({signal_9026, signal_5659}), .c ({signal_9123, signal_5812}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5577 ( .a ({signal_9028, signal_5661}), .b ({signal_9034, signal_5726}), .c ({signal_9124, signal_5813}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5581 ( .a ({signal_8767, signal_5459}), .b ({signal_9029, signal_5665}), .c ({signal_9125, signal_5817}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5582 ( .a ({signal_8935, signal_5627}), .b ({signal_9031, signal_5667}), .c ({signal_9126, signal_5818}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5583 ( .a ({signal_8847, signal_5547}), .b ({signal_9030, signal_5666}), .c ({signal_9127, signal_5819}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5584 ( .a ({signal_9032, signal_5668}), .b ({signal_9035, signal_5739}), .c ({signal_9128, signal_5820}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5585 ( .a ({signal_8743, signal_5463}), .b ({signal_8949, signal_5669}), .c ({signal_9101, signal_5821}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5586 ( .a ({signal_8908, signal_5631}), .b ({signal_8951, signal_5671}), .c ({signal_9102, signal_5822}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5587 ( .a ({signal_8829, signal_5549}), .b ({signal_8950, signal_5670}), .c ({signal_9103, signal_5823}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5588 ( .a ({signal_8952, signal_5672}), .b ({signal_9017, signal_5740}), .c ({signal_9104, signal_5824}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5589 ( .a ({signal_8747, signal_5467}), .b ({signal_8953, signal_5673}), .c ({signal_9105, signal_5825}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5590 ( .a ({signal_8912, signal_5635}), .b ({signal_8955, signal_5675}), .c ({signal_9106, signal_5826}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5591 ( .a ({signal_8831, signal_5551}), .b ({signal_8954, signal_5674}), .c ({signal_9107, signal_5827}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5592 ( .a ({signal_8956, signal_5676}), .b ({signal_9018, signal_5741}), .c ({signal_9108, signal_5828}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5593 ( .a ({signal_8751, signal_5471}), .b ({signal_8957, signal_5677}), .c ({signal_9109, signal_5829}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5594 ( .a ({signal_8916, signal_5639}), .b ({signal_8959, signal_5679}), .c ({signal_9110, signal_5830}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5595 ( .a ({signal_8833, signal_5553}), .b ({signal_8958, signal_5678}), .c ({signal_9111, signal_5831}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5596 ( .a ({signal_8960, signal_5680}), .b ({signal_9019, signal_5742}), .c ({signal_9112, signal_5832}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5597 ( .a ({signal_8755, signal_5475}), .b ({signal_8961, signal_5681}), .c ({signal_9113, signal_5833}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5598 ( .a ({signal_8920, signal_5643}), .b ({signal_8963, signal_5683}), .c ({signal_9114, signal_5834}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5599 ( .a ({signal_8835, signal_5555}), .b ({signal_8962, signal_5682}), .c ({signal_9115, signal_5835}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5600 ( .a ({signal_8964, signal_5684}), .b ({signal_9020, signal_5743}), .c ({signal_9116, signal_5836}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5657 ( .a ({signal_8779, signal_5493}), .b ({signal_9036, signal_5744}), .c ({signal_9161, signal_5893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5658 ( .a ({signal_8968, signal_5688}), .b ({signal_9038, signal_5746}), .c ({signal_9162, signal_5894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5659 ( .a ({signal_8879, signal_5590}), .b ({signal_9037, signal_5745}), .c ({signal_9163, signal_5895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5660 ( .a ({signal_9039, signal_5747}), .b ({signal_9088, signal_5796}), .c ({signal_9164, signal_5896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5661 ( .a ({signal_8783, signal_5497}), .b ({signal_9040, signal_5748}), .c ({signal_9165, signal_5897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5662 ( .a ({signal_8972, signal_5692}), .b ({signal_9042, signal_5750}), .c ({signal_9166, signal_5898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5663 ( .a ({signal_8881, signal_5592}), .b ({signal_9041, signal_5749}), .c ({signal_9167, signal_5899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5664 ( .a ({signal_9043, signal_5751}), .b ({signal_9089, signal_5797}), .c ({signal_9168, signal_5900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5665 ( .a ({signal_8787, signal_5501}), .b ({signal_9044, signal_5752}), .c ({signal_9169, signal_5901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5666 ( .a ({signal_8976, signal_5696}), .b ({signal_9046, signal_5754}), .c ({signal_9170, signal_5902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5667 ( .a ({signal_8883, signal_5594}), .b ({signal_9045, signal_5753}), .c ({signal_9171, signal_5903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5668 ( .a ({signal_9047, signal_5755}), .b ({signal_9090, signal_5798}), .c ({signal_9172, signal_5904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5669 ( .a ({signal_8791, signal_5505}), .b ({signal_9048, signal_5756}), .c ({signal_9173, signal_5905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5670 ( .a ({signal_8980, signal_5700}), .b ({signal_9050, signal_5758}), .c ({signal_9174, signal_5906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5671 ( .a ({signal_8885, signal_5596}), .b ({signal_9049, signal_5757}), .c ({signal_9175, signal_5907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5672 ( .a ({signal_9051, signal_5759}), .b ({signal_9091, signal_5799}), .c ({signal_9176, signal_5908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5673 ( .a ({signal_8795, signal_5509}), .b ({signal_9052, signal_5760}), .c ({signal_9177, signal_5909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5674 ( .a ({signal_8984, signal_5704}), .b ({signal_9054, signal_5762}), .c ({signal_9178, signal_5910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5675 ( .a ({signal_8887, signal_5598}), .b ({signal_9053, signal_5761}), .c ({signal_9179, signal_5911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5676 ( .a ({signal_9055, signal_5763}), .b ({signal_9092, signal_5800}), .c ({signal_9180, signal_5912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5677 ( .a ({signal_8799, signal_5513}), .b ({signal_9056, signal_5764}), .c ({signal_9181, signal_5913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5678 ( .a ({signal_8988, signal_5708}), .b ({signal_9058, signal_5766}), .c ({signal_9182, signal_5914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5679 ( .a ({signal_8889, signal_5600}), .b ({signal_9057, signal_5765}), .c ({signal_9183, signal_5915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5680 ( .a ({signal_9059, signal_5767}), .b ({signal_9093, signal_5801}), .c ({signal_9184, signal_5916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5681 ( .a ({signal_8803, signal_5517}), .b ({signal_9060, signal_5768}), .c ({signal_9185, signal_5917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5682 ( .a ({signal_8992, signal_5712}), .b ({signal_9062, signal_5770}), .c ({signal_9186, signal_5918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5683 ( .a ({signal_8891, signal_5602}), .b ({signal_9061, signal_5769}), .c ({signal_9187, signal_5919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5684 ( .a ({signal_9063, signal_5771}), .b ({signal_9094, signal_5802}), .c ({signal_9188, signal_5920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5685 ( .a ({signal_9118, signal_5804}), .b ({signal_9120, signal_5806}), .c ({signal_9253, signal_5921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5686 ( .a ({signal_9117, signal_5803}), .b ({signal_9119, signal_5805}), .c ({signal_9254, signal_5922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5687 ( .a ({signal_9117, signal_5803}), .b ({signal_9118, signal_5804}), .c ({signal_9255, signal_5923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5688 ( .a ({signal_9119, signal_5805}), .b ({signal_9120, signal_5806}), .c ({signal_9256, signal_5924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5689 ( .a ({signal_8807, signal_5523}), .b ({signal_9064, signal_5772}), .c ({signal_9189, signal_5925}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5690 ( .a ({signal_8996, signal_5717}), .b ({signal_9066, signal_5774}), .c ({signal_9190, signal_5926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5691 ( .a ({signal_8893, signal_5608}), .b ({signal_9065, signal_5773}), .c ({signal_9191, signal_5927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5692 ( .a ({signal_9067, signal_5775}), .b ({signal_9095, signal_5807}), .c ({signal_9192, signal_5928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5693 ( .a ({signal_8811, signal_5527}), .b ({signal_9068, signal_5776}), .c ({signal_9193, signal_5929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5694 ( .a ({signal_9000, signal_5721}), .b ({signal_9070, signal_5778}), .c ({signal_9194, signal_5930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5695 ( .a ({signal_8895, signal_5610}), .b ({signal_9069, signal_5777}), .c ({signal_9195, signal_5931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5696 ( .a ({signal_9071, signal_5779}), .b ({signal_9096, signal_5808}), .c ({signal_9196, signal_5932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5697 ( .a ({signal_8815, signal_5531}), .b ({signal_9072, signal_5780}), .c ({signal_9197, signal_5933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5698 ( .a ({signal_9004, signal_5725}), .b ({signal_9074, signal_5782}), .c ({signal_9198, signal_5934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5699 ( .a ({signal_8897, signal_5612}), .b ({signal_9073, signal_5781}), .c ({signal_9199, signal_5935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5700 ( .a ({signal_9075, signal_5783}), .b ({signal_9097, signal_5809}), .c ({signal_9200, signal_5936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5701 ( .a ({signal_9122, signal_5811}), .b ({signal_9124, signal_5813}), .c ({signal_9257, signal_5937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5702 ( .a ({signal_9121, signal_5810}), .b ({signal_9123, signal_5812}), .c ({signal_9258, signal_5938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5703 ( .a ({signal_9121, signal_5810}), .b ({signal_9122, signal_5811}), .c ({signal_9259, signal_5939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5704 ( .a ({signal_9123, signal_5812}), .b ({signal_9124, signal_5813}), .c ({signal_9260, signal_5940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5705 ( .a ({signal_8819, signal_5537}), .b ({signal_9076, signal_5784}), .c ({signal_9201, signal_5941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5706 ( .a ({signal_9008, signal_5730}), .b ({signal_9078, signal_5786}), .c ({signal_9202, signal_5942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5707 ( .a ({signal_8899, signal_5618}), .b ({signal_9077, signal_5785}), .c ({signal_9203, signal_5943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5708 ( .a ({signal_9079, signal_5787}), .b ({signal_9098, signal_5814}), .c ({signal_9204, signal_5944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5709 ( .a ({signal_8823, signal_5541}), .b ({signal_9080, signal_5788}), .c ({signal_9205, signal_5945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5710 ( .a ({signal_9012, signal_5734}), .b ({signal_9082, signal_5790}), .c ({signal_9206, signal_5946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5711 ( .a ({signal_8901, signal_5620}), .b ({signal_9081, signal_5789}), .c ({signal_9207, signal_5947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5712 ( .a ({signal_9083, signal_5791}), .b ({signal_9099, signal_5815}), .c ({signal_9208, signal_5948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5713 ( .a ({signal_8827, signal_5545}), .b ({signal_9084, signal_5792}), .c ({signal_9209, signal_5949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5714 ( .a ({signal_9016, signal_5738}), .b ({signal_9086, signal_5794}), .c ({signal_9210, signal_5950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5715 ( .a ({signal_8903, signal_5622}), .b ({signal_9085, signal_5793}), .c ({signal_9211, signal_5951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5716 ( .a ({signal_9087, signal_5795}), .b ({signal_9100, signal_5816}), .c ({signal_9212, signal_5952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5717 ( .a ({signal_9126, signal_5818}), .b ({signal_9128, signal_5820}), .c ({signal_9261, signal_5953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5718 ( .a ({signal_9125, signal_5817}), .b ({signal_9127, signal_5819}), .c ({signal_9262, signal_5954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5719 ( .a ({signal_9125, signal_5817}), .b ({signal_9126, signal_5818}), .c ({signal_9263, signal_5955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5720 ( .a ({signal_9127, signal_5819}), .b ({signal_9128, signal_5820}), .c ({signal_9264, signal_5956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5721 ( .a ({signal_9102, signal_5822}), .b ({signal_9104, signal_5824}), .c ({signal_9213, signal_5957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5722 ( .a ({signal_9101, signal_5821}), .b ({signal_9103, signal_5823}), .c ({signal_9214, signal_5958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5723 ( .a ({signal_9101, signal_5821}), .b ({signal_9102, signal_5822}), .c ({signal_9215, signal_5959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5724 ( .a ({signal_9103, signal_5823}), .b ({signal_9104, signal_5824}), .c ({signal_9216, signal_5960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5725 ( .a ({signal_9106, signal_5826}), .b ({signal_9108, signal_5828}), .c ({signal_9217, signal_5961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5726 ( .a ({signal_9105, signal_5825}), .b ({signal_9107, signal_5827}), .c ({signal_9218, signal_5962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5727 ( .a ({signal_9105, signal_5825}), .b ({signal_9106, signal_5826}), .c ({signal_9219, signal_5963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5728 ( .a ({signal_9107, signal_5827}), .b ({signal_9108, signal_5828}), .c ({signal_9220, signal_5964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5729 ( .a ({signal_9110, signal_5830}), .b ({signal_9112, signal_5832}), .c ({signal_9221, signal_5965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5730 ( .a ({signal_9109, signal_5829}), .b ({signal_9111, signal_5831}), .c ({signal_9222, signal_5966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5731 ( .a ({signal_9109, signal_5829}), .b ({signal_9110, signal_5830}), .c ({signal_9223, signal_5967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5732 ( .a ({signal_9111, signal_5831}), .b ({signal_9112, signal_5832}), .c ({signal_9224, signal_5968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5733 ( .a ({signal_9114, signal_5834}), .b ({signal_9116, signal_5836}), .c ({signal_9225, signal_5969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5734 ( .a ({signal_9113, signal_5833}), .b ({signal_9115, signal_5835}), .c ({signal_9226, signal_5970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5735 ( .a ({signal_9113, signal_5833}), .b ({signal_9114, signal_5834}), .c ({signal_9227, signal_5971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5736 ( .a ({signal_9115, signal_5835}), .b ({signal_9116, signal_5836}), .c ({signal_9228, signal_5972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5897 ( .a ({signal_9162, signal_5894}), .b ({signal_9164, signal_5896}), .c ({signal_9401, signal_6133}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5898 ( .a ({signal_9161, signal_5893}), .b ({signal_9163, signal_5895}), .c ({signal_9402, signal_6134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5899 ( .a ({signal_9161, signal_5893}), .b ({signal_9162, signal_5894}), .c ({signal_9403, signal_6135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5900 ( .a ({signal_9163, signal_5895}), .b ({signal_9164, signal_5896}), .c ({signal_9404, signal_6136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5901 ( .a ({signal_9166, signal_5898}), .b ({signal_9168, signal_5900}), .c ({signal_9405, signal_6137}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5902 ( .a ({signal_9165, signal_5897}), .b ({signal_9167, signal_5899}), .c ({signal_9406, signal_6138}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5903 ( .a ({signal_9165, signal_5897}), .b ({signal_9166, signal_5898}), .c ({signal_9407, signal_6139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5904 ( .a ({signal_9167, signal_5899}), .b ({signal_9168, signal_5900}), .c ({signal_9408, signal_6140}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5905 ( .a ({signal_9170, signal_5902}), .b ({signal_9172, signal_5904}), .c ({signal_9409, signal_6141}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5906 ( .a ({signal_9169, signal_5901}), .b ({signal_9171, signal_5903}), .c ({signal_9410, signal_6142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5907 ( .a ({signal_9169, signal_5901}), .b ({signal_9170, signal_5902}), .c ({signal_9411, signal_6143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5908 ( .a ({signal_9171, signal_5903}), .b ({signal_9172, signal_5904}), .c ({signal_9412, signal_6144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5909 ( .a ({signal_9174, signal_5906}), .b ({signal_9176, signal_5908}), .c ({signal_9413, signal_6145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5910 ( .a ({signal_9173, signal_5905}), .b ({signal_9175, signal_5907}), .c ({signal_9414, signal_6146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5911 ( .a ({signal_9173, signal_5905}), .b ({signal_9174, signal_5906}), .c ({signal_9415, signal_6147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5912 ( .a ({signal_9175, signal_5907}), .b ({signal_9176, signal_5908}), .c ({signal_9416, signal_6148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5913 ( .a ({signal_9178, signal_5910}), .b ({signal_9180, signal_5912}), .c ({signal_9417, signal_6149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5914 ( .a ({signal_9177, signal_5909}), .b ({signal_9179, signal_5911}), .c ({signal_9418, signal_6150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5915 ( .a ({signal_9177, signal_5909}), .b ({signal_9178, signal_5910}), .c ({signal_9419, signal_6151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5916 ( .a ({signal_9179, signal_5911}), .b ({signal_9180, signal_5912}), .c ({signal_9420, signal_6152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5917 ( .a ({signal_9182, signal_5914}), .b ({signal_9184, signal_5916}), .c ({signal_9421, signal_6153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5918 ( .a ({signal_9181, signal_5913}), .b ({signal_9183, signal_5915}), .c ({signal_9422, signal_6154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5919 ( .a ({signal_9181, signal_5913}), .b ({signal_9182, signal_5914}), .c ({signal_9423, signal_6155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5920 ( .a ({signal_9183, signal_5915}), .b ({signal_9184, signal_5916}), .c ({signal_9424, signal_6156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5921 ( .a ({signal_9186, signal_5918}), .b ({signal_9188, signal_5920}), .c ({signal_9425, signal_6157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5922 ( .a ({signal_9185, signal_5917}), .b ({signal_9187, signal_5919}), .c ({signal_9426, signal_6158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5923 ( .a ({signal_9185, signal_5917}), .b ({signal_9186, signal_5918}), .c ({signal_9427, signal_6159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5924 ( .a ({signal_9187, signal_5919}), .b ({signal_9188, signal_5920}), .c ({signal_9428, signal_6160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5925 ( .a ({signal_9253, signal_5921}), .b ({signal_9254, signal_5922}), .c ({signal_9493, signal_6161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5929 ( .a ({signal_9190, signal_5926}), .b ({signal_9192, signal_5928}), .c ({signal_9429, signal_6165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5930 ( .a ({signal_9189, signal_5925}), .b ({signal_9191, signal_5927}), .c ({signal_9430, signal_6166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5931 ( .a ({signal_9189, signal_5925}), .b ({signal_9190, signal_5926}), .c ({signal_9431, signal_6167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5932 ( .a ({signal_9191, signal_5927}), .b ({signal_9192, signal_5928}), .c ({signal_9432, signal_6168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5933 ( .a ({signal_9194, signal_5930}), .b ({signal_9196, signal_5932}), .c ({signal_9433, signal_6169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5934 ( .a ({signal_9193, signal_5929}), .b ({signal_9195, signal_5931}), .c ({signal_9434, signal_6170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5935 ( .a ({signal_9193, signal_5929}), .b ({signal_9194, signal_5930}), .c ({signal_9435, signal_6171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5936 ( .a ({signal_9195, signal_5931}), .b ({signal_9196, signal_5932}), .c ({signal_9436, signal_6172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5937 ( .a ({signal_9198, signal_5934}), .b ({signal_9200, signal_5936}), .c ({signal_9437, signal_6173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5938 ( .a ({signal_9197, signal_5933}), .b ({signal_9199, signal_5935}), .c ({signal_9438, signal_6174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5939 ( .a ({signal_9197, signal_5933}), .b ({signal_9198, signal_5934}), .c ({signal_9439, signal_6175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5940 ( .a ({signal_9199, signal_5935}), .b ({signal_9200, signal_5936}), .c ({signal_9440, signal_6176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5941 ( .a ({signal_9257, signal_5937}), .b ({signal_9258, signal_5938}), .c ({signal_9497, signal_6177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5945 ( .a ({signal_9202, signal_5942}), .b ({signal_9204, signal_5944}), .c ({signal_9441, signal_6181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5946 ( .a ({signal_9201, signal_5941}), .b ({signal_9203, signal_5943}), .c ({signal_9442, signal_6182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5947 ( .a ({signal_9201, signal_5941}), .b ({signal_9202, signal_5942}), .c ({signal_9443, signal_6183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5948 ( .a ({signal_9203, signal_5943}), .b ({signal_9204, signal_5944}), .c ({signal_9444, signal_6184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5949 ( .a ({signal_9206, signal_5946}), .b ({signal_9208, signal_5948}), .c ({signal_9445, signal_6185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5950 ( .a ({signal_9205, signal_5945}), .b ({signal_9207, signal_5947}), .c ({signal_9446, signal_6186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5951 ( .a ({signal_9205, signal_5945}), .b ({signal_9206, signal_5946}), .c ({signal_9447, signal_6187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5952 ( .a ({signal_9207, signal_5947}), .b ({signal_9208, signal_5948}), .c ({signal_9448, signal_6188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5953 ( .a ({signal_9210, signal_5950}), .b ({signal_9212, signal_5952}), .c ({signal_9449, signal_6189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5954 ( .a ({signal_9209, signal_5949}), .b ({signal_9211, signal_5951}), .c ({signal_9450, signal_6190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5955 ( .a ({signal_9209, signal_5949}), .b ({signal_9210, signal_5950}), .c ({signal_9451, signal_6191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5956 ( .a ({signal_9211, signal_5951}), .b ({signal_9212, signal_5952}), .c ({signal_9452, signal_6192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5957 ( .a ({signal_9261, signal_5953}), .b ({signal_9262, signal_5954}), .c ({signal_9501, signal_6193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5961 ( .a ({signal_9213, signal_5957}), .b ({signal_9214, signal_5958}), .c ({signal_9453, signal_6197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5965 ( .a ({signal_9217, signal_5961}), .b ({signal_9218, signal_5962}), .c ({signal_9457, signal_6201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5969 ( .a ({signal_9221, signal_5965}), .b ({signal_9222, signal_5966}), .c ({signal_9461, signal_6205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5973 ( .a ({signal_9225, signal_5969}), .b ({signal_9226, signal_5970}), .c ({signal_9465, signal_6209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6095 ( .a ({signal_9401, signal_6133}), .b ({signal_9402, signal_6134}), .c ({signal_9617, signal_6331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6099 ( .a ({signal_9405, signal_6137}), .b ({signal_9406, signal_6138}), .c ({signal_9621, signal_6335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6103 ( .a ({signal_9409, signal_6141}), .b ({signal_9410, signal_6142}), .c ({signal_9625, signal_6339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6107 ( .a ({signal_9413, signal_6145}), .b ({signal_9414, signal_6146}), .c ({signal_9629, signal_6343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6111 ( .a ({signal_9417, signal_6149}), .b ({signal_9418, signal_6150}), .c ({signal_9633, signal_6347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6115 ( .a ({signal_9421, signal_6153}), .b ({signal_9422, signal_6154}), .c ({signal_9637, signal_6351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6119 ( .a ({signal_9425, signal_6157}), .b ({signal_9426, signal_6158}), .c ({signal_9641, signal_6355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6131 ( .a ({signal_9429, signal_6165}), .b ({signal_9430, signal_6166}), .c ({signal_9645, signal_6367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6135 ( .a ({signal_9433, signal_6169}), .b ({signal_9434, signal_6170}), .c ({signal_9649, signal_6371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6139 ( .a ({signal_9437, signal_6173}), .b ({signal_9438, signal_6174}), .c ({signal_9653, signal_6375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6151 ( .a ({signal_9441, signal_6181}), .b ({signal_9442, signal_6182}), .c ({signal_9657, signal_6387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6155 ( .a ({signal_9445, signal_6185}), .b ({signal_9446, signal_6186}), .c ({signal_9661, signal_6391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6159 ( .a ({signal_9449, signal_6189}), .b ({signal_9450, signal_6190}), .c ({signal_9665, signal_6395}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(0)) cell_28 ( .s (signal_402), .b ({signal_10326, signal_3994}), .a ({signal_11320, signal_4122}), .c ({signal_11378, signal_3742}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_29 ( .s (signal_402), .b ({signal_10344, signal_4415}), .a ({signal_11331, signal_4022}), .c ({signal_11379, signal_3642}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_30 ( .s (signal_402), .b ({signal_10516, signal_4414}), .a ({signal_11278, signal_4021}), .c ({signal_11380, signal_3641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_31 ( .s (signal_402), .b ({signal_10515, signal_4413}), .a ({signal_11277, signal_4020}), .c ({signal_11381, signal_3640}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_32 ( .s (signal_402), .b ({signal_10341, signal_4420}), .a ({signal_11025, signal_4019}), .c ({signal_11169, signal_3639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_33 ( .s (signal_402), .b ({signal_10327, signal_3890}), .a ({signal_11276, signal_4018}), .c ({signal_11382, signal_3638}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_34 ( .s (signal_402), .b ({signal_10532, signal_4410}), .a ({signal_11559, signal_4017}), .c ({signal_11575, signal_3637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_35 ( .s (signal_402), .b ({signal_10381, signal_3888}), .a ({signal_11052, signal_4016}), .c ({signal_11170, signal_3636}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_36 ( .s (signal_396), .b ({signal_10380, signal_3887}), .a ({signal_11341, signal_4015}), .c ({signal_11383, signal_3635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_37 ( .s (signal_397), .b ({signal_10379, signal_4407}), .a ({signal_11340, signal_4014}), .c ({signal_11384, signal_3634}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_38 ( .s (signal_398), .b ({signal_10531, signal_4406}), .a ({signal_11285, signal_4013}), .c ({signal_11385, signal_3633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_39 ( .s (signal_399), .b ({signal_10402, signal_3984}), .a ({signal_11146, signal_4112}), .c ({signal_11171, signal_3732}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_40 ( .s (signal_400), .b ({signal_10530, signal_4405}), .a ({signal_11284, signal_4012}), .c ({signal_11386, signal_3632}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_41 ( .s (signal_401), .b ({signal_10376, signal_4412}), .a ({signal_11047, signal_4011}), .c ({signal_11172, signal_3631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_42 ( .s (signal_400), .b ({signal_10331, signal_3882}), .a ({signal_11283, signal_4010}), .c ({signal_11387, signal_3630}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_43 ( .s (signal_399), .b ({signal_10544, signal_4402}), .a ({signal_11562, signal_4009}), .c ({signal_11576, signal_3629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_44 ( .s (signal_399), .b ({signal_10409, signal_3880}), .a ({signal_11044, signal_4008}), .c ({signal_11173, signal_3628}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_45 ( .s (signal_396), .b ({signal_10408, signal_3879}), .a ({signal_11338, signal_4007}), .c ({signal_11388, signal_3627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_46 ( .s (signal_397), .b ({signal_10407, signal_4399}), .a ({signal_11336, signal_4006}), .c ({signal_11389, signal_3626}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_47 ( .s (signal_398), .b ({signal_10543, signal_4398}), .a ({signal_11282, signal_4005}), .c ({signal_11390, signal_3625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_48 ( .s (signal_400), .b ({signal_10542, signal_4397}), .a ({signal_11281, signal_4004}), .c ({signal_11391, signal_3624}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_49 ( .s (signal_401), .b ({signal_10404, signal_4404}), .a ({signal_11038, signal_4003}), .c ({signal_11174, signal_3623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_50 ( .s (signal_401), .b ({signal_10401, signal_3983}), .a ({signal_11377, signal_4111}), .c ({signal_11392, signal_3731}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_51 ( .s (signal_400), .b ({signal_10300, signal_3874}), .a ({signal_11273, signal_4002}), .c ({signal_11393, signal_3622}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_52 ( .s (signal_399), .b ({signal_10502, signal_4394}), .a ({signal_11560, signal_4001}), .c ({signal_11577, signal_3621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_53 ( .s (signal_400), .b ({signal_10320, signal_3872}), .a ({signal_11036, signal_4000}), .c ({signal_11175, signal_3620}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_54 ( .s (signal_401), .b ({signal_10319, signal_3871}), .a ({signal_11334, signal_3999}), .c ({signal_11394, signal_3619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_55 ( .s (signal_397), .b ({signal_10318, signal_4391}), .a ({signal_11333, signal_3998}), .c ({signal_11395, signal_3618}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_56 ( .s (signal_401), .b ({signal_10501, signal_4390}), .a ({signal_11280, signal_3997}), .c ({signal_11396, signal_3617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_57 ( .s (signal_397), .b ({signal_10500, signal_4389}), .a ({signal_11279, signal_3996}), .c ({signal_11397, signal_3616}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_58 ( .s (signal_398), .b ({signal_10315, signal_4396}), .a ({signal_11030, signal_3995}), .c ({signal_11176, signal_3615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_59 ( .s (signal_396), .b ({signal_10400, signal_4503}), .a ({signal_11376, signal_4110}), .c ({signal_11398, signal_3730}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_60 ( .s (signal_398), .b ({signal_10540, signal_4502}), .a ({signal_11319, signal_4109}), .c ({signal_11399, signal_3729}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_61 ( .s (signal_397), .b ({signal_10539, signal_4501}), .a ({signal_11318, signal_4108}), .c ({signal_11400, signal_3728}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_62 ( .s (signal_398), .b ({signal_10397, signal_4508}), .a ({signal_11141, signal_4107}), .c ({signal_11177, signal_3727}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_63 ( .s (signal_396), .b ({signal_10334, signal_3978}), .a ({signal_11317, signal_4106}), .c ({signal_11401, signal_3726}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_64 ( .s (signal_399), .b ({signal_10553, signal_4498}), .a ({signal_11574, signal_4105}), .c ({signal_11578, signal_3725}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_65 ( .s (signal_400), .b ({signal_10430, signal_3976}), .a ({signal_11138, signal_4104}), .c ({signal_11178, signal_3724}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_66 ( .s (signal_401), .b ({signal_10429, signal_3975}), .a ({signal_11374, signal_4103}), .c ({signal_11402, signal_3723}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_67 ( .s (signal_399), .b ({signal_10529, signal_4514}), .a ({signal_11573, signal_4121}), .c ({signal_11579, signal_3741}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_68 ( .s (signal_400), .b ({signal_10428, signal_4495}), .a ({signal_11372, signal_4102}), .c ({signal_11403, signal_3722}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_69 ( .s (signal_397), .b ({signal_10552, signal_4494}), .a ({signal_11316, signal_4101}), .c ({signal_11404, signal_3721}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_70 ( .s (signal_398), .b ({signal_10551, signal_4493}), .a ({signal_11315, signal_4100}), .c ({signal_11405, signal_3720}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_71 ( .s (signal_396), .b ({signal_10425, signal_4500}), .a ({signal_11132, signal_4099}), .c ({signal_11179, signal_3719}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_72 ( .s (signal_401), .b ({signal_10325, signal_3970}), .a ({signal_11314, signal_4098}), .c ({signal_11406, signal_3718}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_73 ( .s (signal_399), .b ({signal_10526, signal_4490}), .a ({signal_11572, signal_4097}), .c ({signal_11580, signal_3717}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_74 ( .s (signal_397), .b ({signal_10367, signal_3968}), .a ({signal_11129, signal_4096}), .c ({signal_11180, signal_3716}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_75 ( .s (signal_398), .b ({signal_10366, signal_3967}), .a ({signal_11370, signal_4095}), .c ({signal_11407, signal_3715}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_76 ( .s (signal_396), .b ({signal_10365, signal_4487}), .a ({signal_11369, signal_4094}), .c ({signal_11408, signal_3714}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_77 ( .s (signal_400), .b ({signal_10525, signal_4486}), .a ({signal_11313, signal_4093}), .c ({signal_11409, signal_3713}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_78 ( .s (signal_396), .b ({signal_10374, signal_3992}), .a ({signal_11125, signal_4120}), .c ({signal_11181, signal_3740}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_79 ( .s (signal_401), .b ({signal_10524, signal_4485}), .a ({signal_11312, signal_4092}), .c ({signal_11410, signal_3712}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_80 ( .s (signal_399), .b ({signal_10362, signal_4492}), .a ({signal_11123, signal_4091}), .c ({signal_11182, signal_3711}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_81 ( .s (signal_397), .b ({signal_10329, signal_3962}), .a ({signal_11308, signal_4090}), .c ({signal_11411, signal_3710}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_82 ( .s (signal_398), .b ({signal_10538, signal_4482}), .a ({signal_11569, signal_4089}), .c ({signal_11581, signal_3709}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_83 ( .s (signal_396), .b ({signal_10395, signal_3960}), .a ({signal_11094, signal_4088}), .c ({signal_11183, signal_3708}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_84 ( .s (signal_401), .b ({signal_10394, signal_3959}), .a ({signal_11356, signal_4087}), .c ({signal_11412, signal_3707}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_85 ( .s (signal_401), .b ({signal_10393, signal_4479}), .a ({signal_11355, signal_4086}), .c ({signal_11413, signal_3706}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_86 ( .s (signal_401), .b ({signal_10537, signal_4478}), .a ({signal_11300, signal_4085}), .c ({signal_11414, signal_3705}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_87 ( .s (signal_401), .b ({signal_10536, signal_4477}), .a ({signal_11299, signal_4084}), .c ({signal_11415, signal_3704}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_88 ( .s (signal_401), .b ({signal_10390, signal_4484}), .a ({signal_11087, signal_4083}), .c ({signal_11184, signal_3703}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_89 ( .s (signal_401), .b ({signal_10373, signal_3991}), .a ({signal_11368, signal_4119}), .c ({signal_11416, signal_3739}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_90 ( .s (signal_401), .b ({signal_10333, signal_3954}), .a ({signal_11298, signal_4082}), .c ({signal_11417, signal_3702}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_91 ( .s (signal_401), .b ({signal_10550, signal_4474}), .a ({signal_11567, signal_4081}), .c ({signal_11582, signal_3701}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_92 ( .s (signal_401), .b ({signal_10423, signal_3952}), .a ({signal_11114, signal_4080}), .c ({signal_11185, signal_3700}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_93 ( .s (signal_401), .b ({signal_10422, signal_3951}), .a ({signal_11365, signal_4079}), .c ({signal_11418, signal_3699}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_94 ( .s (signal_401), .b ({signal_10421, signal_4471}), .a ({signal_11364, signal_4078}), .c ({signal_11419, signal_3698}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_95 ( .s (signal_401), .b ({signal_10549, signal_4470}), .a ({signal_11307, signal_4077}), .c ({signal_11420, signal_3697}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_96 ( .s (signal_400), .b ({signal_10548, signal_4469}), .a ({signal_11306, signal_4076}), .c ({signal_11421, signal_3696}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_97 ( .s (signal_400), .b ({signal_10418, signal_4476}), .a ({signal_11109, signal_4075}), .c ({signal_11186, signal_3695}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_98 ( .s (signal_400), .b ({signal_10324, signal_3946}), .a ({signal_11305, signal_4074}), .c ({signal_11422, signal_3694}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_99 ( .s (signal_400), .b ({signal_10523, signal_4466}), .a ({signal_11570, signal_4073}), .c ({signal_11583, signal_3693}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_100 ( .s (signal_400), .b ({signal_10372, signal_4511}), .a ({signal_11367, signal_4118}), .c ({signal_11423, signal_3738}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_101 ( .s (signal_400), .b ({signal_10360, signal_3944}), .a ({signal_11106, signal_4072}), .c ({signal_11187, signal_3692}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_102 ( .s (signal_400), .b ({signal_10359, signal_3943}), .a ({signal_11362, signal_4071}), .c ({signal_11424, signal_3691}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_103 ( .s (signal_400), .b ({signal_10358, signal_4463}), .a ({signal_11360, signal_4070}), .c ({signal_11425, signal_3690}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_104 ( .s (signal_400), .b ({signal_10522, signal_4462}), .a ({signal_11304, signal_4069}), .c ({signal_11426, signal_3689}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_105 ( .s (signal_400), .b ({signal_10521, signal_4461}), .a ({signal_11303, signal_4068}), .c ({signal_11427, signal_3688}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_106 ( .s (signal_400), .b ({signal_10355, signal_4468}), .a ({signal_11100, signal_4067}), .c ({signal_11188, signal_3687}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_107 ( .s (signal_400), .b ({signal_10298, signal_3938}), .a ({signal_11275, signal_4066}), .c ({signal_11428, signal_3686}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_108 ( .s (signal_399), .b ({signal_10496, signal_4458}), .a ({signal_11568, signal_4065}), .c ({signal_11584, signal_3685}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_109 ( .s (signal_399), .b ({signal_10306, signal_3936}), .a ({signal_11098, signal_4064}), .c ({signal_11189, signal_3684}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_110 ( .s (signal_399), .b ({signal_10305, signal_3935}), .a ({signal_11358, signal_4063}), .c ({signal_11429, signal_3683}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_111 ( .s (signal_399), .b ({signal_10528, signal_4510}), .a ({signal_11311, signal_4117}), .c ({signal_11430, signal_3737}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_112 ( .s (signal_399), .b ({signal_10304, signal_4455}), .a ({signal_11357, signal_4062}), .c ({signal_11431, signal_3682}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_113 ( .s (signal_399), .b ({signal_10495, signal_4454}), .a ({signal_11302, signal_4061}), .c ({signal_11432, signal_3681}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_114 ( .s (signal_399), .b ({signal_10494, signal_4453}), .a ({signal_11301, signal_4060}), .c ({signal_11433, signal_3680}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_115 ( .s (signal_399), .b ({signal_10301, signal_4460}), .a ({signal_11092, signal_4059}), .c ({signal_11190, signal_3679}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_116 ( .s (signal_399), .b ({signal_10332, signal_3930}), .a ({signal_11297, signal_4058}), .c ({signal_11434, signal_3678}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_117 ( .s (signal_399), .b ({signal_10547, signal_4450}), .a ({signal_11565, signal_4057}), .c ({signal_11585, signal_3677}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_118 ( .s (signal_399), .b ({signal_10416, signal_3928}), .a ({signal_11063, signal_4056}), .c ({signal_11191, signal_3676}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_119 ( .s (signal_399), .b ({signal_10415, signal_3927}), .a ({signal_11344, signal_4055}), .c ({signal_11435, signal_3675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_120 ( .s (signal_398), .b ({signal_10414, signal_4447}), .a ({signal_11343, signal_4054}), .c ({signal_11436, signal_3674}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_121 ( .s (signal_398), .b ({signal_10546, signal_4446}), .a ({signal_11289, signal_4053}), .c ({signal_11437, signal_3673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_122 ( .s (signal_398), .b ({signal_10527, signal_4509}), .a ({signal_11310, signal_4116}), .c ({signal_11438, signal_3736}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_123 ( .s (signal_398), .b ({signal_10545, signal_4445}), .a ({signal_11288, signal_4052}), .c ({signal_11439, signal_3672}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_124 ( .s (signal_398), .b ({signal_10411, signal_4452}), .a ({signal_11056, signal_4051}), .c ({signal_11192, signal_3671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_125 ( .s (signal_398), .b ({signal_10323, signal_3922}), .a ({signal_11287, signal_4050}), .c ({signal_11440, signal_3670}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_126 ( .s (signal_398), .b ({signal_10520, signal_4442}), .a ({signal_11563, signal_4049}), .c ({signal_11586, signal_3669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_127 ( .s (signal_398), .b ({signal_10353, signal_3920}), .a ({signal_11083, signal_4048}), .c ({signal_11193, signal_3668}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_128 ( .s (signal_398), .b ({signal_10352, signal_3919}), .a ({signal_11353, signal_4047}), .c ({signal_11441, signal_3667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_129 ( .s (signal_398), .b ({signal_10351, signal_4439}), .a ({signal_11352, signal_4046}), .c ({signal_11442, signal_3666}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_130 ( .s (signal_398), .b ({signal_10519, signal_4438}), .a ({signal_11296, signal_4045}), .c ({signal_11443, signal_3665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_131 ( .s (signal_398), .b ({signal_10518, signal_4437}), .a ({signal_11295, signal_4044}), .c ({signal_11444, signal_3664}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_132 ( .s (signal_397), .b ({signal_10348, signal_4444}), .a ({signal_11078, signal_4043}), .c ({signal_11194, signal_3663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_133 ( .s (signal_397), .b ({signal_10369, signal_4516}), .a ({signal_11118, signal_4115}), .c ({signal_11195, signal_3735}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_134 ( .s (signal_397), .b ({signal_10328, signal_3914}), .a ({signal_11294, signal_4042}), .c ({signal_11445, signal_3662}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_135 ( .s (signal_397), .b ({signal_10535, signal_4434}), .a ({signal_11566, signal_4041}), .c ({signal_11587, signal_3661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_136 ( .s (signal_397), .b ({signal_10388, signal_3912}), .a ({signal_11075, signal_4040}), .c ({signal_11196, signal_3660}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_137 ( .s (signal_397), .b ({signal_10387, signal_3911}), .a ({signal_11350, signal_4039}), .c ({signal_11446, signal_3659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_138 ( .s (signal_397), .b ({signal_10386, signal_4431}), .a ({signal_11348, signal_4038}), .c ({signal_11447, signal_3658}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_139 ( .s (signal_397), .b ({signal_10534, signal_4430}), .a ({signal_11293, signal_4037}), .c ({signal_11448, signal_3657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_140 ( .s (signal_397), .b ({signal_10533, signal_4429}), .a ({signal_11292, signal_4036}), .c ({signal_11449, signal_3656}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_141 ( .s (signal_397), .b ({signal_10383, signal_4436}), .a ({signal_11069, signal_4035}), .c ({signal_11197, signal_3655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_142 ( .s (signal_397), .b ({signal_10299, signal_3906}), .a ({signal_11274, signal_4034}), .c ({signal_11450, signal_3654}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_143 ( .s (signal_397), .b ({signal_10499, signal_4426}), .a ({signal_11564, signal_4033}), .c ({signal_11588, signal_3653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_144 ( .s (signal_396), .b ({signal_10330, signal_3986}), .a ({signal_11309, signal_4114}), .c ({signal_11451, signal_3734}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_145 ( .s (signal_396), .b ({signal_10313, signal_3904}), .a ({signal_11067, signal_4032}), .c ({signal_11198, signal_3652}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_146 ( .s (signal_396), .b ({signal_10312, signal_3903}), .a ({signal_11346, signal_4031}), .c ({signal_11452, signal_3651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_147 ( .s (signal_396), .b ({signal_10311, signal_4423}), .a ({signal_11345, signal_4030}), .c ({signal_11453, signal_3650}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_148 ( .s (signal_396), .b ({signal_10498, signal_4422}), .a ({signal_11291, signal_4029}), .c ({signal_11454, signal_3649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_149 ( .s (signal_396), .b ({signal_10497, signal_4421}), .a ({signal_11290, signal_4028}), .c ({signal_11455, signal_3648}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_150 ( .s (signal_396), .b ({signal_10308, signal_4428}), .a ({signal_11061, signal_4027}), .c ({signal_11199, signal_3647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_151 ( .s (signal_396), .b ({signal_10322, signal_3898}), .a ({signal_11286, signal_4026}), .c ({signal_11456, signal_3646}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_152 ( .s (signal_396), .b ({signal_10517, signal_4418}), .a ({signal_11561, signal_4025}), .c ({signal_11589, signal_3645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_153 ( .s (signal_396), .b ({signal_10346, signal_3896}), .a ({signal_11032, signal_4024}), .c ({signal_11200, signal_3644}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_154 ( .s (signal_396), .b ({signal_10345, signal_3895}), .a ({signal_11332, signal_4023}), .c ({signal_11457, signal_3643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_155 ( .s (signal_396), .b ({signal_10541, signal_4506}), .a ({signal_11571, signal_4113}), .c ({signal_11590, signal_3733}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_291 ( .s (reset), .b ({signal_11378, signal_3742}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({signal_11592, signal_421}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_294 ( .s (reset), .b ({signal_11579, signal_3741}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({signal_11758, signal_423}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_297 ( .s (reset), .b ({signal_11181, signal_3740}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({signal_11459, signal_425}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_300 ( .s (reset), .b ({signal_11416, signal_3739}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({signal_11594, signal_427}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_303 ( .s (reset), .b ({signal_11423, signal_3738}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({signal_11596, signal_429}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_306 ( .s (reset), .b ({signal_11430, signal_3737}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({signal_11598, signal_431}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_309 ( .s (reset), .b ({signal_11438, signal_3736}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({signal_11600, signal_433}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_312 ( .s (reset), .b ({signal_11195, signal_3735}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({signal_11461, signal_435}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_315 ( .s (reset), .b ({signal_11451, signal_3734}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({signal_11602, signal_437}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_318 ( .s (reset), .b ({signal_11590, signal_3733}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({signal_11760, signal_439}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_321 ( .s (reset), .b ({signal_11171, signal_3732}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({signal_11463, signal_441}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_324 ( .s (reset), .b ({signal_11392, signal_3731}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({signal_11604, signal_443}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_327 ( .s (reset), .b ({signal_11398, signal_3730}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({signal_11606, signal_445}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_330 ( .s (reset), .b ({signal_11399, signal_3729}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({signal_11608, signal_447}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_333 ( .s (reset), .b ({signal_11400, signal_3728}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({signal_11610, signal_449}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_336 ( .s (reset), .b ({signal_11177, signal_3727}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({signal_11465, signal_451}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_339 ( .s (reset), .b ({signal_11401, signal_3726}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({signal_11612, signal_453}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_342 ( .s (reset), .b ({signal_11578, signal_3725}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({signal_11762, signal_455}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_345 ( .s (reset), .b ({signal_11178, signal_3724}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({signal_11467, signal_457}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_348 ( .s (reset), .b ({signal_11402, signal_3723}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({signal_11614, signal_459}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_351 ( .s (reset), .b ({signal_11403, signal_3722}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({signal_11616, signal_461}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_354 ( .s (reset), .b ({signal_11404, signal_3721}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({signal_11618, signal_463}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_357 ( .s (reset), .b ({signal_11405, signal_3720}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({signal_11620, signal_465}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_360 ( .s (reset), .b ({signal_11179, signal_3719}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({signal_11469, signal_467}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_363 ( .s (reset), .b ({signal_11406, signal_3718}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({signal_11622, signal_469}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_366 ( .s (reset), .b ({signal_11580, signal_3717}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({signal_11764, signal_471}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_369 ( .s (reset), .b ({signal_11180, signal_3716}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({signal_11471, signal_473}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_372 ( .s (reset), .b ({signal_11407, signal_3715}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({signal_11624, signal_475}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_375 ( .s (reset), .b ({signal_11408, signal_3714}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({signal_11626, signal_477}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_378 ( .s (reset), .b ({signal_11409, signal_3713}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({signal_11628, signal_479}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_381 ( .s (reset), .b ({signal_11410, signal_3712}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({signal_11630, signal_481}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_384 ( .s (reset), .b ({signal_11182, signal_3711}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({signal_11473, signal_483}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_387 ( .s (reset), .b ({signal_11411, signal_3710}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_11632, signal_485}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_390 ( .s (reset), .b ({signal_11581, signal_3709}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_11766, signal_487}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_393 ( .s (reset), .b ({signal_11183, signal_3708}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_11475, signal_489}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_396 ( .s (reset), .b ({signal_11412, signal_3707}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_11634, signal_491}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_399 ( .s (reset), .b ({signal_11413, signal_3706}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_11636, signal_493}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_402 ( .s (reset), .b ({signal_11414, signal_3705}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_11638, signal_495}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_405 ( .s (reset), .b ({signal_11415, signal_3704}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_11640, signal_497}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_408 ( .s (reset), .b ({signal_11184, signal_3703}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_11477, signal_499}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_411 ( .s (reset), .b ({signal_11417, signal_3702}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_11642, signal_501}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_414 ( .s (reset), .b ({signal_11582, signal_3701}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_11768, signal_503}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_417 ( .s (reset), .b ({signal_11185, signal_3700}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_11479, signal_505}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_420 ( .s (reset), .b ({signal_11418, signal_3699}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_11644, signal_507}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_423 ( .s (reset), .b ({signal_11419, signal_3698}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_11646, signal_509}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_426 ( .s (reset), .b ({signal_11420, signal_3697}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_11648, signal_511}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_429 ( .s (reset), .b ({signal_11421, signal_3696}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_11650, signal_513}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_432 ( .s (reset), .b ({signal_11186, signal_3695}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_11481, signal_515}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_435 ( .s (reset), .b ({signal_11422, signal_3694}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_11652, signal_517}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_438 ( .s (reset), .b ({signal_11583, signal_3693}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_11770, signal_519}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_441 ( .s (reset), .b ({signal_11187, signal_3692}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_11483, signal_521}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_444 ( .s (reset), .b ({signal_11424, signal_3691}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_11654, signal_523}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_447 ( .s (reset), .b ({signal_11425, signal_3690}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_11656, signal_525}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_450 ( .s (reset), .b ({signal_11426, signal_3689}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_11658, signal_527}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_453 ( .s (reset), .b ({signal_11427, signal_3688}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_11660, signal_529}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_456 ( .s (reset), .b ({signal_11188, signal_3687}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_11485, signal_531}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_459 ( .s (reset), .b ({signal_11428, signal_3686}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_11662, signal_533}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_462 ( .s (reset), .b ({signal_11584, signal_3685}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_11772, signal_535}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_465 ( .s (reset), .b ({signal_11189, signal_3684}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_11487, signal_537}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_468 ( .s (reset), .b ({signal_11429, signal_3683}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_11664, signal_539}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_471 ( .s (reset), .b ({signal_11431, signal_3682}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_11666, signal_541}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_474 ( .s (reset), .b ({signal_11432, signal_3681}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_11668, signal_543}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_477 ( .s (reset), .b ({signal_11433, signal_3680}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_11670, signal_545}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_480 ( .s (reset), .b ({signal_11190, signal_3679}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_11489, signal_547}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_483 ( .s (reset), .b ({signal_11434, signal_3678}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_11672, signal_549}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_486 ( .s (reset), .b ({signal_11585, signal_3677}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_11774, signal_551}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_489 ( .s (reset), .b ({signal_11191, signal_3676}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_11491, signal_553}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_492 ( .s (reset), .b ({signal_11435, signal_3675}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_11674, signal_555}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_495 ( .s (reset), .b ({signal_11436, signal_3674}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_11676, signal_557}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_498 ( .s (reset), .b ({signal_11437, signal_3673}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_11678, signal_559}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_501 ( .s (reset), .b ({signal_11439, signal_3672}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_11680, signal_561}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_504 ( .s (reset), .b ({signal_11192, signal_3671}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_11493, signal_563}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_507 ( .s (reset), .b ({signal_11440, signal_3670}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_11682, signal_565}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_510 ( .s (reset), .b ({signal_11586, signal_3669}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_11776, signal_567}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_513 ( .s (reset), .b ({signal_11193, signal_3668}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_11495, signal_569}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_516 ( .s (reset), .b ({signal_11441, signal_3667}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_11684, signal_571}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_519 ( .s (reset), .b ({signal_11442, signal_3666}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_11686, signal_573}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_522 ( .s (reset), .b ({signal_11443, signal_3665}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_11688, signal_575}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_525 ( .s (reset), .b ({signal_11444, signal_3664}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_11690, signal_577}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_528 ( .s (reset), .b ({signal_11194, signal_3663}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_11497, signal_579}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_531 ( .s (reset), .b ({signal_11445, signal_3662}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_11692, signal_581}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_534 ( .s (reset), .b ({signal_11587, signal_3661}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_11778, signal_583}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_537 ( .s (reset), .b ({signal_11196, signal_3660}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_11499, signal_585}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_540 ( .s (reset), .b ({signal_11446, signal_3659}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_11694, signal_587}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_543 ( .s (reset), .b ({signal_11447, signal_3658}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_11696, signal_589}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_546 ( .s (reset), .b ({signal_11448, signal_3657}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_11698, signal_591}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_549 ( .s (reset), .b ({signal_11449, signal_3656}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_11700, signal_593}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_552 ( .s (reset), .b ({signal_11197, signal_3655}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_11501, signal_595}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_555 ( .s (reset), .b ({signal_11450, signal_3654}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_11702, signal_597}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_558 ( .s (reset), .b ({signal_11588, signal_3653}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_11780, signal_599}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_561 ( .s (reset), .b ({signal_11198, signal_3652}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_11503, signal_601}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_564 ( .s (reset), .b ({signal_11452, signal_3651}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_11704, signal_603}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_567 ( .s (reset), .b ({signal_11453, signal_3650}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_11706, signal_605}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_570 ( .s (reset), .b ({signal_11454, signal_3649}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_11708, signal_607}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_573 ( .s (reset), .b ({signal_11455, signal_3648}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_11710, signal_609}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_576 ( .s (reset), .b ({signal_11199, signal_3647}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_11505, signal_611}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_579 ( .s (reset), .b ({signal_11456, signal_3646}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_11712, signal_613}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_582 ( .s (reset), .b ({signal_11589, signal_3645}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_11782, signal_615}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_585 ( .s (reset), .b ({signal_11200, signal_3644}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_11507, signal_617}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_588 ( .s (reset), .b ({signal_11457, signal_3643}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_11714, signal_619}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_591 ( .s (reset), .b ({signal_11379, signal_3642}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_11716, signal_621}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_594 ( .s (reset), .b ({signal_11380, signal_3641}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_11718, signal_623}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_597 ( .s (reset), .b ({signal_11381, signal_3640}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_11720, signal_625}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_600 ( .s (reset), .b ({signal_11169, signal_3639}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_11509, signal_627}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_603 ( .s (reset), .b ({signal_11382, signal_3638}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_11722, signal_629}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_606 ( .s (reset), .b ({signal_11575, signal_3637}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_11784, signal_631}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_609 ( .s (reset), .b ({signal_11170, signal_3636}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_11511, signal_633}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_612 ( .s (reset), .b ({signal_11383, signal_3635}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_11724, signal_635}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_615 ( .s (reset), .b ({signal_11384, signal_3634}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_11726, signal_637}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_618 ( .s (reset), .b ({signal_11385, signal_3633}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_11728, signal_639}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_621 ( .s (reset), .b ({signal_11386, signal_3632}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_11730, signal_641}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_624 ( .s (reset), .b ({signal_11172, signal_3631}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_11513, signal_643}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_627 ( .s (reset), .b ({signal_11387, signal_3630}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_11732, signal_645}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_630 ( .s (reset), .b ({signal_11576, signal_3629}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_11786, signal_647}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_633 ( .s (reset), .b ({signal_11173, signal_3628}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_11515, signal_649}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_636 ( .s (reset), .b ({signal_11388, signal_3627}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_11734, signal_651}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_639 ( .s (reset), .b ({signal_11389, signal_3626}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_11736, signal_653}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_642 ( .s (reset), .b ({signal_11390, signal_3625}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_11738, signal_655}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_645 ( .s (reset), .b ({signal_11391, signal_3624}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_11740, signal_657}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_648 ( .s (reset), .b ({signal_11174, signal_3623}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_11517, signal_659}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_651 ( .s (reset), .b ({signal_11393, signal_3622}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_11742, signal_661}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_654 ( .s (reset), .b ({signal_11577, signal_3621}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_11788, signal_663}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_657 ( .s (reset), .b ({signal_11175, signal_3620}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_11519, signal_665}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_660 ( .s (reset), .b ({signal_11394, signal_3619}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_11744, signal_667}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_663 ( .s (reset), .b ({signal_11395, signal_3618}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_11746, signal_669}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_666 ( .s (reset), .b ({signal_11396, signal_3617}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_11748, signal_671}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_669 ( .s (reset), .b ({signal_11397, signal_3616}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_11750, signal_673}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_672 ( .s (reset), .b ({signal_11176, signal_3615}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_11521, signal_675}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3155 ( .s (reset), .b ({signal_11022, signal_4250}), .a ({key_s1[0], key_s0[0]}), .c ({signal_11202, signal_2853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3158 ( .s (reset), .b ({signal_11326, signal_4249}), .a ({key_s1[1], key_s0[1]}), .c ({signal_11523, signal_2855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3161 ( .s (reset), .b ({signal_11154, signal_4248}), .a ({key_s1[2], key_s0[2]}), .c ({signal_11204, signal_2857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3164 ( .s (reset), .b ({signal_11153, signal_4247}), .a ({key_s1[3], key_s0[3]}), .c ({signal_11206, signal_2859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3167 ( .s (reset), .b ({signal_11152, signal_4246}), .a ({key_s1[4], key_s0[4]}), .c ({signal_11208, signal_2861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3170 ( .s (reset), .b ({signal_11323, signal_4245}), .a ({key_s1[5], key_s0[5]}), .c ({signal_11525, signal_2863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3173 ( .s (reset), .b ({signal_11322, signal_4244}), .a ({key_s1[6], key_s0[6]}), .c ({signal_11527, signal_2865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3176 ( .s (reset), .b ({signal_11149, signal_4243}), .a ({key_s1[7], key_s0[7]}), .c ({signal_11210, signal_2867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3179 ( .s (reset), .b ({signal_11011, signal_4242}), .a ({key_s1[8], key_s0[8]}), .c ({signal_11212, signal_2869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3182 ( .s (reset), .b ({signal_11321, signal_4241}), .a ({key_s1[9], key_s0[9]}), .c ({signal_11529, signal_2871}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3185 ( .s (reset), .b ({signal_11168, signal_4240}), .a ({key_s1[10], key_s0[10]}), .c ({signal_11214, signal_2873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3188 ( .s (reset), .b ({signal_11167, signal_4239}), .a ({key_s1[11], key_s0[11]}), .c ({signal_11216, signal_2875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3191 ( .s (reset), .b ({signal_11166, signal_4238}), .a ({key_s1[12], key_s0[12]}), .c ({signal_11218, signal_2877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3194 ( .s (reset), .b ({signal_11329, signal_4237}), .a ({key_s1[13], key_s0[13]}), .c ({signal_11531, signal_2879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3197 ( .s (reset), .b ({signal_11328, signal_4236}), .a ({key_s1[14], key_s0[14]}), .c ({signal_11533, signal_2881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3200 ( .s (reset), .b ({signal_11163, signal_4235}), .a ({key_s1[15], key_s0[15]}), .c ({signal_11220, signal_2883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3203 ( .s (reset), .b ({signal_11019, signal_4234}), .a ({key_s1[16], key_s0[16]}), .c ({signal_11222, signal_2885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3206 ( .s (reset), .b ({signal_11327, signal_4233}), .a ({key_s1[17], key_s0[17]}), .c ({signal_11535, signal_2887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3209 ( .s (reset), .b ({signal_11161, signal_4232}), .a ({key_s1[18], key_s0[18]}), .c ({signal_11224, signal_2889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3212 ( .s (reset), .b ({signal_11160, signal_4231}), .a ({key_s1[19], key_s0[19]}), .c ({signal_11226, signal_2891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3215 ( .s (reset), .b ({signal_11158, signal_4230}), .a ({key_s1[20], key_s0[20]}), .c ({signal_11228, signal_2893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3218 ( .s (reset), .b ({signal_11325, signal_4229}), .a ({key_s1[21], key_s0[21]}), .c ({signal_11537, signal_2895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3221 ( .s (reset), .b ({signal_11324, signal_4228}), .a ({key_s1[22], key_s0[22]}), .c ({signal_11539, signal_2897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3224 ( .s (reset), .b ({signal_11155, signal_4227}), .a ({key_s1[23], key_s0[23]}), .c ({signal_11230, signal_2899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3227 ( .s (reset), .b ({signal_11272, signal_4226}), .a ({key_s1[24], key_s0[24]}), .c ({signal_11541, signal_2901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3230 ( .s (reset), .b ({signal_11558, signal_4225}), .a ({key_s1[25], key_s0[25]}), .c ({signal_11752, signal_2903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3233 ( .s (reset), .b ({signal_11270, signal_4224}), .a ({key_s1[26], key_s0[26]}), .c ({signal_11543, signal_2905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3236 ( .s (reset), .b ({signal_11269, signal_4223}), .a ({key_s1[27], key_s0[27]}), .c ({signal_11545, signal_2907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3239 ( .s (reset), .b ({signal_11268, signal_4222}), .a ({key_s1[28], key_s0[28]}), .c ({signal_11547, signal_2909}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3242 ( .s (reset), .b ({signal_11557, signal_4221}), .a ({key_s1[29], key_s0[29]}), .c ({signal_11754, signal_2911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3245 ( .s (reset), .b ({signal_11556, signal_4220}), .a ({key_s1[30], key_s0[30]}), .c ({signal_11756, signal_2913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3248 ( .s (reset), .b ({signal_11265, signal_4219}), .a ({key_s1[31], key_s0[31]}), .c ({signal_11549, signal_2915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3251 ( .s (reset), .b ({signal_10795, signal_4218}), .a ({key_s1[32], key_s0[32]}), .c ({signal_10937, signal_2917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3254 ( .s (reset), .b ({signal_11017, signal_4217}), .a ({key_s1[33], key_s0[33]}), .c ({signal_11232, signal_2919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3257 ( .s (reset), .b ({signal_10919, signal_4216}), .a ({key_s1[34], key_s0[34]}), .c ({signal_10939, signal_2921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3260 ( .s (reset), .b ({signal_10918, signal_4215}), .a ({key_s1[35], key_s0[35]}), .c ({signal_10941, signal_2923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3263 ( .s (reset), .b ({signal_10917, signal_4214}), .a ({key_s1[36], key_s0[36]}), .c ({signal_10943, signal_2925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3266 ( .s (reset), .b ({signal_11014, signal_4213}), .a ({key_s1[37], key_s0[37]}), .c ({signal_11234, signal_2927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3269 ( .s (reset), .b ({signal_11013, signal_4212}), .a ({key_s1[38], key_s0[38]}), .c ({signal_11236, signal_2929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3272 ( .s (reset), .b ({signal_10914, signal_4211}), .a ({key_s1[39], key_s0[39]}), .c ({signal_10945, signal_2931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3275 ( .s (reset), .b ({signal_10785, signal_4210}), .a ({key_s1[40], key_s0[40]}), .c ({signal_10947, signal_2933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3278 ( .s (reset), .b ({signal_11012, signal_4209}), .a ({key_s1[41], key_s0[41]}), .c ({signal_11238, signal_2935}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3281 ( .s (reset), .b ({signal_10934, signal_4208}), .a ({key_s1[42], key_s0[42]}), .c ({signal_10949, signal_2937}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3284 ( .s (reset), .b ({signal_10933, signal_4207}), .a ({key_s1[43], key_s0[43]}), .c ({signal_10951, signal_2939}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3287 ( .s (reset), .b ({signal_10932, signal_4206}), .a ({key_s1[44], key_s0[44]}), .c ({signal_10953, signal_2941}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3290 ( .s (reset), .b ({signal_11021, signal_4205}), .a ({key_s1[45], key_s0[45]}), .c ({signal_11240, signal_2943}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3293 ( .s (reset), .b ({signal_11020, signal_4204}), .a ({key_s1[46], key_s0[46]}), .c ({signal_11242, signal_2945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3296 ( .s (reset), .b ({signal_10929, signal_4203}), .a ({key_s1[47], key_s0[47]}), .c ({signal_10955, signal_2947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3299 ( .s (reset), .b ({signal_10792, signal_4202}), .a ({key_s1[48], key_s0[48]}), .c ({signal_10957, signal_2949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3302 ( .s (reset), .b ({signal_11018, signal_4201}), .a ({key_s1[49], key_s0[49]}), .c ({signal_11244, signal_2951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3305 ( .s (reset), .b ({signal_10926, signal_4200}), .a ({key_s1[50], key_s0[50]}), .c ({signal_10959, signal_2953}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3308 ( .s (reset), .b ({signal_10925, signal_4199}), .a ({key_s1[51], key_s0[51]}), .c ({signal_10961, signal_2955}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3311 ( .s (reset), .b ({signal_10923, signal_4198}), .a ({key_s1[52], key_s0[52]}), .c ({signal_10963, signal_2957}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3314 ( .s (reset), .b ({signal_11016, signal_4197}), .a ({key_s1[53], key_s0[53]}), .c ({signal_11246, signal_2959}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3317 ( .s (reset), .b ({signal_11015, signal_4196}), .a ({key_s1[54], key_s0[54]}), .c ({signal_11248, signal_2961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3320 ( .s (reset), .b ({signal_10920, signal_4195}), .a ({key_s1[55], key_s0[55]}), .c ({signal_10965, signal_2963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3323 ( .s (reset), .b ({signal_11007, signal_4194}), .a ({key_s1[56], key_s0[56]}), .c ({signal_11250, signal_2965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3326 ( .s (reset), .b ({signal_11271, signal_4193}), .a ({key_s1[57], key_s0[57]}), .c ({signal_11551, signal_2967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3329 ( .s (reset), .b ({signal_11005, signal_4192}), .a ({key_s1[58], key_s0[58]}), .c ({signal_11252, signal_2969}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3332 ( .s (reset), .b ({signal_11004, signal_4191}), .a ({key_s1[59], key_s0[59]}), .c ({signal_11254, signal_2971}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3335 ( .s (reset), .b ({signal_11003, signal_4190}), .a ({key_s1[60], key_s0[60]}), .c ({signal_11256, signal_2973}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3338 ( .s (reset), .b ({signal_11267, signal_4189}), .a ({key_s1[61], key_s0[61]}), .c ({signal_11553, signal_2975}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3341 ( .s (reset), .b ({signal_11266, signal_4188}), .a ({key_s1[62], key_s0[62]}), .c ({signal_11555, signal_2977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3344 ( .s (reset), .b ({signal_11000, signal_4187}), .a ({key_s1[63], key_s0[63]}), .c ({signal_11258, signal_2979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3347 ( .s (reset), .b ({signal_10565, signal_4186}), .a ({key_s1[64], key_s0[64]}), .c ({signal_10707, signal_2981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3350 ( .s (reset), .b ({signal_10790, signal_4185}), .a ({key_s1[65], key_s0[65]}), .c ({signal_10967, signal_2983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3353 ( .s (reset), .b ({signal_10689, signal_4184}), .a ({key_s1[66], key_s0[66]}), .c ({signal_10709, signal_2985}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3356 ( .s (reset), .b ({signal_10688, signal_4183}), .a ({key_s1[67], key_s0[67]}), .c ({signal_10711, signal_2987}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3359 ( .s (reset), .b ({signal_10687, signal_4182}), .a ({key_s1[68], key_s0[68]}), .c ({signal_10713, signal_2989}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3362 ( .s (reset), .b ({signal_10787, signal_4181}), .a ({key_s1[69], key_s0[69]}), .c ({signal_10969, signal_2991}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3365 ( .s (reset), .b ({signal_10786, signal_4180}), .a ({key_s1[70], key_s0[70]}), .c ({signal_10971, signal_2993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3368 ( .s (reset), .b ({signal_10684, signal_4179}), .a ({key_s1[71], key_s0[71]}), .c ({signal_10715, signal_2995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3371 ( .s (reset), .b ({signal_10554, signal_4178}), .a ({key_s1[72], key_s0[72]}), .c ({signal_10717, signal_2997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3374 ( .s (reset), .b ({signal_10784, signal_4177}), .a ({key_s1[73], key_s0[73]}), .c ({signal_10973, signal_2999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3377 ( .s (reset), .b ({signal_10704, signal_4176}), .a ({key_s1[74], key_s0[74]}), .c ({signal_10719, signal_3001}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3380 ( .s (reset), .b ({signal_10703, signal_4175}), .a ({key_s1[75], key_s0[75]}), .c ({signal_10721, signal_3003}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3383 ( .s (reset), .b ({signal_10702, signal_4174}), .a ({key_s1[76], key_s0[76]}), .c ({signal_10723, signal_3005}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3386 ( .s (reset), .b ({signal_10794, signal_4173}), .a ({key_s1[77], key_s0[77]}), .c ({signal_10975, signal_3007}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3389 ( .s (reset), .b ({signal_10793, signal_4172}), .a ({key_s1[78], key_s0[78]}), .c ({signal_10977, signal_3009}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3392 ( .s (reset), .b ({signal_10699, signal_4171}), .a ({key_s1[79], key_s0[79]}), .c ({signal_10725, signal_3011}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3395 ( .s (reset), .b ({signal_10556, signal_4170}), .a ({key_s1[80], key_s0[80]}), .c ({signal_10727, signal_3013}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3398 ( .s (reset), .b ({signal_10791, signal_4169}), .a ({key_s1[81], key_s0[81]}), .c ({signal_10979, signal_3015}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3401 ( .s (reset), .b ({signal_10696, signal_4168}), .a ({key_s1[82], key_s0[82]}), .c ({signal_10729, signal_3017}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3404 ( .s (reset), .b ({signal_10695, signal_4167}), .a ({key_s1[83], key_s0[83]}), .c ({signal_10731, signal_3019}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3407 ( .s (reset), .b ({signal_10693, signal_4166}), .a ({key_s1[84], key_s0[84]}), .c ({signal_10733, signal_3021}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3410 ( .s (reset), .b ({signal_10789, signal_4165}), .a ({key_s1[85], key_s0[85]}), .c ({signal_10981, signal_3023}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3413 ( .s (reset), .b ({signal_10788, signal_4164}), .a ({key_s1[86], key_s0[86]}), .c ({signal_10983, signal_3025}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3416 ( .s (reset), .b ({signal_10690, signal_4163}), .a ({key_s1[87], key_s0[87]}), .c ({signal_10735, signal_3027}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3419 ( .s (reset), .b ({signal_10768, signal_4162}), .a ({key_s1[88], key_s0[88]}), .c ({signal_10985, signal_3029}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3422 ( .s (reset), .b ({signal_11006, signal_4161}), .a ({key_s1[89], key_s0[89]}), .c ({signal_11260, signal_3031}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3425 ( .s (reset), .b ({signal_10767, signal_4160}), .a ({key_s1[90], key_s0[90]}), .c ({signal_10987, signal_3033}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3428 ( .s (reset), .b ({signal_10766, signal_4159}), .a ({key_s1[91], key_s0[91]}), .c ({signal_10989, signal_3035}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3431 ( .s (reset), .b ({signal_10765, signal_4158}), .a ({key_s1[92], key_s0[92]}), .c ({signal_10991, signal_3037}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3434 ( .s (reset), .b ({signal_11002, signal_4157}), .a ({key_s1[93], key_s0[93]}), .c ({signal_11262, signal_3039}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3437 ( .s (reset), .b ({signal_11001, signal_4156}), .a ({key_s1[94], key_s0[94]}), .c ({signal_11264, signal_3041}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3440 ( .s (reset), .b ({signal_10764, signal_4155}), .a ({key_s1[95], key_s0[95]}), .c ({signal_10993, signal_3043}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3443 ( .s (reset), .b ({signal_10337, signal_4154}), .a ({key_s1[96], key_s0[96]}), .c ({signal_10457, signal_3045}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3446 ( .s (reset), .b ({signal_10555, signal_4153}), .a ({key_s1[97], key_s0[97]}), .c ({signal_10737, signal_3047}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3449 ( .s (reset), .b ({signal_10434, signal_4152}), .a ({key_s1[98], key_s0[98]}), .c ({signal_10459, signal_3049}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3452 ( .s (reset), .b ({signal_10433, signal_4151}), .a ({key_s1[99], key_s0[99]}), .c ({signal_10461, signal_3051}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3455 ( .s (reset), .b ({signal_10454, signal_4150}), .a ({key_s1[100], key_s0[100]}), .c ({signal_10463, signal_3053}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3458 ( .s (reset), .b ({signal_10564, signal_4149}), .a ({key_s1[101], key_s0[101]}), .c ({signal_10739, signal_3055}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3461 ( .s (reset), .b ({signal_10563, signal_4148}), .a ({key_s1[102], key_s0[102]}), .c ({signal_10741, signal_3057}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3464 ( .s (reset), .b ({signal_10451, signal_4147}), .a ({key_s1[103], key_s0[103]}), .c ({signal_10465, signal_3059}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3467 ( .s (reset), .b ({signal_10336, signal_4146}), .a ({key_s1[104], key_s0[104]}), .c ({signal_10467, signal_3061}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3470 ( .s (reset), .b ({signal_10562, signal_4145}), .a ({key_s1[105], key_s0[105]}), .c ({signal_10743, signal_3063}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3473 ( .s (reset), .b ({signal_10449, signal_4144}), .a ({key_s1[106], key_s0[106]}), .c ({signal_10469, signal_3065}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3476 ( .s (reset), .b ({signal_10448, signal_4143}), .a ({key_s1[107], key_s0[107]}), .c ({signal_10471, signal_3067}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3479 ( .s (reset), .b ({signal_10447, signal_4142}), .a ({key_s1[108], key_s0[108]}), .c ({signal_10473, signal_3069}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3482 ( .s (reset), .b ({signal_10561, signal_4141}), .a ({key_s1[109], key_s0[109]}), .c ({signal_10745, signal_3071}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3485 ( .s (reset), .b ({signal_10560, signal_4140}), .a ({key_s1[110], key_s0[110]}), .c ({signal_10747, signal_3073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3488 ( .s (reset), .b ({signal_10444, signal_4139}), .a ({key_s1[111], key_s0[111]}), .c ({signal_10475, signal_3075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3491 ( .s (reset), .b ({signal_10335, signal_4138}), .a ({key_s1[112], key_s0[112]}), .c ({signal_10477, signal_3077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3494 ( .s (reset), .b ({signal_10559, signal_4137}), .a ({key_s1[113], key_s0[113]}), .c ({signal_10749, signal_3079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3497 ( .s (reset), .b ({signal_10442, signal_4136}), .a ({key_s1[114], key_s0[114]}), .c ({signal_10479, signal_3081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3500 ( .s (reset), .b ({signal_10441, signal_4135}), .a ({key_s1[115], key_s0[115]}), .c ({signal_10481, signal_3083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3503 ( .s (reset), .b ({signal_10440, signal_4134}), .a ({key_s1[116], key_s0[116]}), .c ({signal_10483, signal_3085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3506 ( .s (reset), .b ({signal_10558, signal_4133}), .a ({key_s1[117], key_s0[117]}), .c ({signal_10751, signal_3087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3509 ( .s (reset), .b ({signal_10557, signal_4132}), .a ({key_s1[118], key_s0[118]}), .c ({signal_10753, signal_3089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3512 ( .s (reset), .b ({signal_10437, signal_4131}), .a ({key_s1[119], key_s0[119]}), .c ({signal_10485, signal_3091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3515 ( .s (reset), .b ({signal_10490, signal_4130}), .a ({key_s1[120], key_s0[120]}), .c ({signal_10755, signal_3093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3518 ( .s (reset), .b ({signal_10771, signal_4129}), .a ({key_s1[121], key_s0[121]}), .c ({signal_10995, signal_3095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3521 ( .s (reset), .b ({signal_10489, signal_4128}), .a ({key_s1[122], key_s0[122]}), .c ({signal_10757, signal_3097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3524 ( .s (reset), .b ({signal_10488, signal_4127}), .a ({key_s1[123], key_s0[123]}), .c ({signal_10759, signal_3099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3527 ( .s (reset), .b ({signal_10487, signal_4126}), .a ({key_s1[124], key_s0[124]}), .c ({signal_10761, signal_3101}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3530 ( .s (reset), .b ({signal_10770, signal_4125}), .a ({key_s1[125], key_s0[125]}), .c ({signal_10997, signal_3103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3533 ( .s (reset), .b ({signal_10769, signal_4124}), .a ({key_s1[126], key_s0[126]}), .c ({signal_10999, signal_3105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(0)) cell_3536 ( .s (reset), .b ({signal_10486, signal_4123}), .a ({key_s1[127], key_s0[127]}), .c ({signal_10763, signal_3107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3561 ( .a ({signal_7661, signal_4347}), .b ({signal_11000, signal_4187}), .c ({signal_11265, signal_4219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3562 ( .a ({signal_7503, signal_4315}), .b ({signal_10764, signal_4155}), .c ({signal_11000, signal_4187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3563 ( .a ({signal_7527, signal_4283}), .b ({signal_10486, signal_4123}), .c ({signal_10764, signal_4155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3564 ( .a ({signal_7658, signal_4348}), .b ({signal_11266, signal_4188}), .c ({signal_11556, signal_4220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3565 ( .a ({signal_7500, signal_4316}), .b ({signal_11001, signal_4156}), .c ({signal_11266, signal_4188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3566 ( .a ({signal_7524, signal_4284}), .b ({signal_10769, signal_4124}), .c ({signal_11001, signal_4156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3571 ( .a ({signal_7652, signal_4349}), .b ({signal_11267, signal_4189}), .c ({signal_11557, signal_4221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3572 ( .a ({signal_7497, signal_4317}), .b ({signal_11002, signal_4157}), .c ({signal_11267, signal_4189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3573 ( .a ({signal_7521, signal_4285}), .b ({signal_10770, signal_4125}), .c ({signal_11002, signal_4157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3574 ( .a ({signal_7649, signal_4350}), .b ({signal_11003, signal_4190}), .c ({signal_11268, signal_4222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3575 ( .a ({signal_7494, signal_4318}), .b ({signal_10765, signal_4158}), .c ({signal_11003, signal_4190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3576 ( .a ({signal_7518, signal_4286}), .b ({signal_10487, signal_4126}), .c ({signal_10765, signal_4158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3577 ( .a ({signal_7646, signal_4351}), .b ({signal_11004, signal_4191}), .c ({signal_11269, signal_4223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3578 ( .a ({signal_7491, signal_4319}), .b ({signal_10766, signal_4159}), .c ({signal_11004, signal_4191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3579 ( .a ({signal_7515, signal_4287}), .b ({signal_10488, signal_4127}), .c ({signal_10766, signal_4159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3580 ( .a ({signal_7643, signal_4352}), .b ({signal_11005, signal_4192}), .c ({signal_11270, signal_4224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3581 ( .a ({signal_7488, signal_4320}), .b ({signal_10767, signal_4160}), .c ({signal_11005, signal_4192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3582 ( .a ({signal_7512, signal_4288}), .b ({signal_10489, signal_4128}), .c ({signal_10767, signal_4160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3583 ( .a ({signal_7640, signal_4353}), .b ({signal_11271, signal_4193}), .c ({signal_11558, signal_4225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3584 ( .a ({signal_7485, signal_4321}), .b ({signal_11006, signal_4161}), .c ({signal_11271, signal_4193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3585 ( .a ({signal_7509, signal_4289}), .b ({signal_10771, signal_4129}), .c ({signal_11006, signal_4161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3586 ( .a ({signal_7637, signal_4354}), .b ({signal_11007, signal_4194}), .c ({signal_11272, signal_4226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3587 ( .a ({signal_7482, signal_4322}), .b ({signal_10768, signal_4162}), .c ({signal_11007, signal_4194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3588 ( .a ({signal_7506, signal_4290}), .b ({signal_10490, signal_4130}), .c ({signal_10768, signal_4162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3629 ( .a ({signal_7479, signal_4251}), .b ({signal_10293, signal_4517}), .c ({signal_10486, signal_4123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3630 ( .a ({signal_7476, signal_4252}), .b ({signal_10491, signal_4518}), .c ({signal_10769, signal_4124}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3631 ( .a ({signal_7473, signal_4253}), .b ({signal_10492, signal_4519}), .c ({signal_10770, signal_4125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3632 ( .a ({signal_7470, signal_4254}), .b ({signal_10294, signal_4520}), .c ({signal_10487, signal_4126}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3633 ( .a ({signal_7467, signal_4255}), .b ({signal_10295, signal_4521}), .c ({signal_10488, signal_4127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3634 ( .a ({signal_7464, signal_4256}), .b ({signal_10296, signal_4522}), .c ({signal_10489, signal_4128}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3635 ( .a ({signal_7461, signal_4257}), .b ({signal_10493, signal_4523}), .c ({signal_10771, signal_4129}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3636 ( .a ({signal_7458, signal_4258}), .b ({signal_10297, signal_4524}), .c ({signal_10490, signal_4130}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3667 ( .a ({signal_10265, signal_3116}), .b ({1'b0, signal_393}), .c ({signal_10293, signal_4517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3668 ( .a ({signal_10338, signal_3115}), .b ({1'b0, signal_394}), .c ({signal_10491, signal_4518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3669 ( .a ({signal_10339, signal_3114}), .b ({1'b0, signal_4379}), .c ({signal_10492, signal_4519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3670 ( .a ({signal_10268, signal_3113}), .b ({1'b0, signal_4380}), .c ({signal_10294, signal_4520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3671 ( .a ({signal_10269, signal_3112}), .b ({1'b0, signal_4381}), .c ({signal_10295, signal_4521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3672 ( .a ({signal_10270, signal_3111}), .b ({1'b0, signal_4382}), .c ({signal_10296, signal_4522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3673 ( .a ({signal_10340, signal_3110}), .b ({1'b0, signal_4383}), .c ({signal_10493, signal_4523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_3674 ( .a ({signal_10118, signal_3109}), .b ({1'b0, signal_4384}), .c ({signal_10297, signal_4524}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5601 ( .a ({signal_8271, signal_4903}), .b ({signal_9120, signal_5806}), .clk (clk), .r (Fresh[320]), .c ({signal_9229, signal_5837}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5602 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_9119, signal_5805}), .clk (clk), .r (Fresh[321]), .c ({signal_9230, signal_5838}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5603 ( .a ({signal_8074, signal_4690}), .b ({signal_9118, signal_5804}), .clk (clk), .r (Fresh[322]), .c ({signal_9231, signal_5839}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5604 ( .a ({signal_8274, signal_4906}), .b ({signal_9117, signal_5803}), .clk (clk), .r (Fresh[323]), .c ({signal_9232, signal_5840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5605 ( .a ({signal_8276, signal_4908}), .b ({signal_9120, signal_5806}), .clk (clk), .r (Fresh[324]), .c ({signal_9233, signal_5841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5606 ( .a ({signal_8078, signal_4694}), .b ({signal_9119, signal_5805}), .clk (clk), .r (Fresh[325]), .c ({signal_9234, signal_5842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5607 ( .a ({signal_8079, signal_4695}), .b ({signal_9118, signal_5804}), .clk (clk), .r (Fresh[326]), .c ({signal_9235, signal_5843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5608 ( .a ({signal_8275, signal_4907}), .b ({signal_9117, signal_5803}), .clk (clk), .r (Fresh[327]), .c ({signal_9236, signal_5844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5609 ( .a ({signal_8278, signal_4934}), .b ({signal_9124, signal_5813}), .clk (clk), .r (Fresh[328]), .c ({signal_9237, signal_5845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5610 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_9123, signal_5812}), .clk (clk), .r (Fresh[329]), .c ({signal_9238, signal_5846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5611 ( .a ({signal_8082, signal_4728}), .b ({signal_9122, signal_5811}), .clk (clk), .r (Fresh[330]), .c ({signal_9239, signal_5847}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5612 ( .a ({signal_8281, signal_4937}), .b ({signal_9121, signal_5810}), .clk (clk), .r (Fresh[331]), .c ({signal_9240, signal_5848}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5613 ( .a ({signal_8283, signal_4939}), .b ({signal_9124, signal_5813}), .clk (clk), .r (Fresh[332]), .c ({signal_9241, signal_5849}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5614 ( .a ({signal_8086, signal_4732}), .b ({signal_9123, signal_5812}), .clk (clk), .r (Fresh[333]), .c ({signal_9242, signal_5850}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5615 ( .a ({signal_8087, signal_4733}), .b ({signal_9122, signal_5811}), .clk (clk), .r (Fresh[334]), .c ({signal_9243, signal_5851}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5616 ( .a ({signal_8282, signal_4938}), .b ({signal_9121, signal_5810}), .clk (clk), .r (Fresh[335]), .c ({signal_9244, signal_5852}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5617 ( .a ({signal_8285, signal_4965}), .b ({signal_9128, signal_5820}), .clk (clk), .r (Fresh[336]), .c ({signal_9245, signal_5853}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5618 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_9127, signal_5819}), .clk (clk), .r (Fresh[337]), .c ({signal_9246, signal_5854}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5619 ( .a ({signal_8090, signal_4766}), .b ({signal_9126, signal_5818}), .clk (clk), .r (Fresh[338]), .c ({signal_9247, signal_5855}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5620 ( .a ({signal_8288, signal_4968}), .b ({signal_9125, signal_5817}), .clk (clk), .r (Fresh[339]), .c ({signal_9248, signal_5856}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5621 ( .a ({signal_8290, signal_4970}), .b ({signal_9128, signal_5820}), .clk (clk), .r (Fresh[340]), .c ({signal_9249, signal_5857}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5622 ( .a ({signal_8094, signal_4770}), .b ({signal_9127, signal_5819}), .clk (clk), .r (Fresh[341]), .c ({signal_9250, signal_5858}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5623 ( .a ({signal_8095, signal_4771}), .b ({signal_9126, signal_5818}), .clk (clk), .r (Fresh[342]), .c ({signal_9251, signal_5859}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5624 ( .a ({signal_8289, signal_4969}), .b ({signal_9125, signal_5817}), .clk (clk), .r (Fresh[343]), .c ({signal_9252, signal_5860}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5625 ( .a ({signal_8225, signal_4972}), .b ({signal_9104, signal_5824}), .clk (clk), .r (Fresh[344]), .c ({signal_9129, signal_5861}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5626 ( .a ({signal_7610, signal_4362}), .b ({signal_9103, signal_5823}), .clk (clk), .r (Fresh[345]), .c ({signal_9130, signal_5862}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5627 ( .a ({signal_8042, signal_4774}), .b ({signal_9102, signal_5822}), .clk (clk), .r (Fresh[346]), .c ({signal_9131, signal_5863}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5628 ( .a ({signal_8228, signal_4975}), .b ({signal_9101, signal_5821}), .clk (clk), .r (Fresh[347]), .c ({signal_9132, signal_5864}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5629 ( .a ({signal_8230, signal_4977}), .b ({signal_9104, signal_5824}), .clk (clk), .r (Fresh[348]), .c ({signal_9133, signal_5865}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5630 ( .a ({signal_8046, signal_4778}), .b ({signal_9103, signal_5823}), .clk (clk), .r (Fresh[349]), .c ({signal_9134, signal_5866}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5631 ( .a ({signal_8047, signal_4779}), .b ({signal_9102, signal_5822}), .clk (clk), .r (Fresh[350]), .c ({signal_9135, signal_5867}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5632 ( .a ({signal_8229, signal_4976}), .b ({signal_9101, signal_5821}), .clk (clk), .r (Fresh[351]), .c ({signal_9136, signal_5868}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5633 ( .a ({signal_8232, signal_4979}), .b ({signal_9108, signal_5828}), .clk (clk), .r (Fresh[352]), .c ({signal_9137, signal_5869}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5634 ( .a ({signal_7823, signal_4370}), .b ({signal_9107, signal_5827}), .clk (clk), .r (Fresh[353]), .c ({signal_9138, signal_5870}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5635 ( .a ({signal_8050, signal_4782}), .b ({signal_9106, signal_5826}), .clk (clk), .r (Fresh[354]), .c ({signal_9139, signal_5871}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5636 ( .a ({signal_8235, signal_4982}), .b ({signal_9105, signal_5825}), .clk (clk), .r (Fresh[355]), .c ({signal_9140, signal_5872}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5637 ( .a ({signal_8237, signal_4984}), .b ({signal_9108, signal_5828}), .clk (clk), .r (Fresh[356]), .c ({signal_9141, signal_5873}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5638 ( .a ({signal_8054, signal_4786}), .b ({signal_9107, signal_5827}), .clk (clk), .r (Fresh[357]), .c ({signal_9142, signal_5874}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5639 ( .a ({signal_8055, signal_4787}), .b ({signal_9106, signal_5826}), .clk (clk), .r (Fresh[358]), .c ({signal_9143, signal_5875}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5640 ( .a ({signal_8236, signal_4983}), .b ({signal_9105, signal_5825}), .clk (clk), .r (Fresh[359]), .c ({signal_9144, signal_5876}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5641 ( .a ({signal_8239, signal_4986}), .b ({signal_9112, signal_5832}), .clk (clk), .r (Fresh[360]), .c ({signal_9145, signal_5877}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5642 ( .a ({signal_7529, signal_4378}), .b ({signal_9111, signal_5831}), .clk (clk), .r (Fresh[361]), .c ({signal_9146, signal_5878}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5643 ( .a ({signal_8058, signal_4790}), .b ({signal_9110, signal_5830}), .clk (clk), .r (Fresh[362]), .c ({signal_9147, signal_5879}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5644 ( .a ({signal_8242, signal_4989}), .b ({signal_9109, signal_5829}), .clk (clk), .r (Fresh[363]), .c ({signal_9148, signal_5880}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5645 ( .a ({signal_8244, signal_4991}), .b ({signal_9112, signal_5832}), .clk (clk), .r (Fresh[364]), .c ({signal_9149, signal_5881}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5646 ( .a ({signal_8062, signal_4794}), .b ({signal_9111, signal_5831}), .clk (clk), .r (Fresh[365]), .c ({signal_9150, signal_5882}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5647 ( .a ({signal_8063, signal_4795}), .b ({signal_9110, signal_5830}), .clk (clk), .r (Fresh[366]), .c ({signal_9151, signal_5883}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5648 ( .a ({signal_8243, signal_4990}), .b ({signal_9109, signal_5829}), .clk (clk), .r (Fresh[367]), .c ({signal_9152, signal_5884}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5649 ( .a ({signal_8246, signal_4993}), .b ({signal_9116, signal_5836}), .clk (clk), .r (Fresh[368]), .c ({signal_9153, signal_5885}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5650 ( .a ({signal_7637, signal_4354}), .b ({signal_9115, signal_5835}), .clk (clk), .r (Fresh[369]), .c ({signal_9154, signal_5886}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5651 ( .a ({signal_8066, signal_4798}), .b ({signal_9114, signal_5834}), .clk (clk), .r (Fresh[370]), .c ({signal_9155, signal_5887}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5652 ( .a ({signal_8249, signal_4996}), .b ({signal_9113, signal_5833}), .clk (clk), .r (Fresh[371]), .c ({signal_9156, signal_5888}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5653 ( .a ({signal_8251, signal_4998}), .b ({signal_9116, signal_5836}), .clk (clk), .r (Fresh[372]), .c ({signal_9157, signal_5889}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5654 ( .a ({signal_8070, signal_4802}), .b ({signal_9115, signal_5835}), .clk (clk), .r (Fresh[373]), .c ({signal_9158, signal_5890}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5655 ( .a ({signal_8071, signal_4803}), .b ({signal_9114, signal_5834}), .clk (clk), .r (Fresh[374]), .c ({signal_9159, signal_5891}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5656 ( .a ({signal_8250, signal_4997}), .b ({signal_9113, signal_5833}), .clk (clk), .r (Fresh[375]), .c ({signal_9160, signal_5892}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5737 ( .a ({signal_8382, signal_5099}), .b ({signal_9164, signal_5896}), .clk (clk), .r (Fresh[376]), .c ({signal_9265, signal_5973}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5738 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_9163, signal_5895}), .clk (clk), .r (Fresh[377]), .c ({signal_9266, signal_5974}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5739 ( .a ({signal_8122, signal_4848}), .b ({signal_9162, signal_5894}), .clk (clk), .r (Fresh[378]), .c ({signal_9267, signal_5975}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5740 ( .a ({signal_8385, signal_5102}), .b ({signal_9161, signal_5893}), .clk (clk), .r (Fresh[379]), .c ({signal_9268, signal_5976}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5741 ( .a ({signal_8387, signal_5104}), .b ({signal_9164, signal_5896}), .clk (clk), .r (Fresh[380]), .c ({signal_9269, signal_5977}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5742 ( .a ({signal_8126, signal_4852}), .b ({signal_9163, signal_5895}), .clk (clk), .r (Fresh[381]), .c ({signal_9270, signal_5978}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5743 ( .a ({signal_8127, signal_4853}), .b ({signal_9162, signal_5894}), .clk (clk), .r (Fresh[382]), .c ({signal_9271, signal_5979}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5744 ( .a ({signal_8386, signal_5103}), .b ({signal_9161, signal_5893}), .clk (clk), .r (Fresh[383]), .c ({signal_9272, signal_5980}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5745 ( .a ({signal_8389, signal_5106}), .b ({signal_9168, signal_5900}), .clk (clk), .r (Fresh[384]), .c ({signal_9273, signal_5981}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5746 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_9167, signal_5899}), .clk (clk), .r (Fresh[385]), .c ({signal_9274, signal_5982}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5747 ( .a ({signal_8130, signal_4856}), .b ({signal_9166, signal_5898}), .clk (clk), .r (Fresh[386]), .c ({signal_9275, signal_5983}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5748 ( .a ({signal_8392, signal_5109}), .b ({signal_9165, signal_5897}), .clk (clk), .r (Fresh[387]), .c ({signal_9276, signal_5984}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5749 ( .a ({signal_8394, signal_5111}), .b ({signal_9168, signal_5900}), .clk (clk), .r (Fresh[388]), .c ({signal_9277, signal_5985}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5750 ( .a ({signal_8134, signal_4860}), .b ({signal_9167, signal_5899}), .clk (clk), .r (Fresh[389]), .c ({signal_9278, signal_5986}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5751 ( .a ({signal_8135, signal_4861}), .b ({signal_9166, signal_5898}), .clk (clk), .r (Fresh[390]), .c ({signal_9279, signal_5987}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5752 ( .a ({signal_8393, signal_5110}), .b ({signal_9165, signal_5897}), .clk (clk), .r (Fresh[391]), .c ({signal_9280, signal_5988}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5753 ( .a ({signal_8396, signal_5113}), .b ({signal_9172, signal_5904}), .clk (clk), .r (Fresh[392]), .c ({signal_9281, signal_5989}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5754 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_9171, signal_5903}), .clk (clk), .r (Fresh[393]), .c ({signal_9282, signal_5990}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5755 ( .a ({signal_8138, signal_4864}), .b ({signal_9170, signal_5902}), .clk (clk), .r (Fresh[394]), .c ({signal_9283, signal_5991}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5756 ( .a ({signal_8399, signal_5116}), .b ({signal_9169, signal_5901}), .clk (clk), .r (Fresh[395]), .c ({signal_9284, signal_5992}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5757 ( .a ({signal_8401, signal_5118}), .b ({signal_9172, signal_5904}), .clk (clk), .r (Fresh[396]), .c ({signal_9285, signal_5993}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5758 ( .a ({signal_8142, signal_4868}), .b ({signal_9171, signal_5903}), .clk (clk), .r (Fresh[397]), .c ({signal_9286, signal_5994}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5759 ( .a ({signal_8143, signal_4869}), .b ({signal_9170, signal_5902}), .clk (clk), .r (Fresh[398]), .c ({signal_9287, signal_5995}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5760 ( .a ({signal_8400, signal_5117}), .b ({signal_9169, signal_5901}), .clk (clk), .r (Fresh[399]), .c ({signal_9288, signal_5996}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5761 ( .a ({signal_8403, signal_5120}), .b ({signal_9176, signal_5908}), .clk (clk), .r (Fresh[400]), .c ({signal_9289, signal_5997}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5762 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_9175, signal_5907}), .clk (clk), .r (Fresh[401]), .c ({signal_9290, signal_5998}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5763 ( .a ({signal_8146, signal_4872}), .b ({signal_9174, signal_5906}), .clk (clk), .r (Fresh[402]), .c ({signal_9291, signal_5999}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5764 ( .a ({signal_8406, signal_5123}), .b ({signal_9173, signal_5905}), .clk (clk), .r (Fresh[403]), .c ({signal_9292, signal_6000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5765 ( .a ({signal_8408, signal_5125}), .b ({signal_9176, signal_5908}), .clk (clk), .r (Fresh[404]), .c ({signal_9293, signal_6001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5766 ( .a ({signal_8150, signal_4876}), .b ({signal_9175, signal_5907}), .clk (clk), .r (Fresh[405]), .c ({signal_9294, signal_6002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5767 ( .a ({signal_8151, signal_4877}), .b ({signal_9174, signal_5906}), .clk (clk), .r (Fresh[406]), .c ({signal_9295, signal_6003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5768 ( .a ({signal_8407, signal_5124}), .b ({signal_9173, signal_5905}), .clk (clk), .r (Fresh[407]), .c ({signal_9296, signal_6004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5769 ( .a ({signal_8410, signal_5127}), .b ({signal_9180, signal_5912}), .clk (clk), .r (Fresh[408]), .c ({signal_9297, signal_6005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5770 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_9179, signal_5911}), .clk (clk), .r (Fresh[409]), .c ({signal_9298, signal_6006}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5771 ( .a ({signal_8154, signal_4880}), .b ({signal_9178, signal_5910}), .clk (clk), .r (Fresh[410]), .c ({signal_9299, signal_6007}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5772 ( .a ({signal_8413, signal_5130}), .b ({signal_9177, signal_5909}), .clk (clk), .r (Fresh[411]), .c ({signal_9300, signal_6008}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5773 ( .a ({signal_8415, signal_5132}), .b ({signal_9180, signal_5912}), .clk (clk), .r (Fresh[412]), .c ({signal_9301, signal_6009}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5774 ( .a ({signal_8158, signal_4884}), .b ({signal_9179, signal_5911}), .clk (clk), .r (Fresh[413]), .c ({signal_9302, signal_6010}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5775 ( .a ({signal_8159, signal_4885}), .b ({signal_9178, signal_5910}), .clk (clk), .r (Fresh[414]), .c ({signal_9303, signal_6011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5776 ( .a ({signal_8414, signal_5131}), .b ({signal_9177, signal_5909}), .clk (clk), .r (Fresh[415]), .c ({signal_9304, signal_6012}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5777 ( .a ({signal_8417, signal_5134}), .b ({signal_9184, signal_5916}), .clk (clk), .r (Fresh[416]), .c ({signal_9305, signal_6013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5778 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_9183, signal_5915}), .clk (clk), .r (Fresh[417]), .c ({signal_9306, signal_6014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5779 ( .a ({signal_8162, signal_4888}), .b ({signal_9182, signal_5914}), .clk (clk), .r (Fresh[418]), .c ({signal_9307, signal_6015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5780 ( .a ({signal_8420, signal_5137}), .b ({signal_9181, signal_5913}), .clk (clk), .r (Fresh[419]), .c ({signal_9308, signal_6016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5781 ( .a ({signal_8422, signal_5139}), .b ({signal_9184, signal_5916}), .clk (clk), .r (Fresh[420]), .c ({signal_9309, signal_6017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5782 ( .a ({signal_8166, signal_4892}), .b ({signal_9183, signal_5915}), .clk (clk), .r (Fresh[421]), .c ({signal_9310, signal_6018}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5783 ( .a ({signal_8167, signal_4893}), .b ({signal_9182, signal_5914}), .clk (clk), .r (Fresh[422]), .c ({signal_9311, signal_6019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5784 ( .a ({signal_8421, signal_5138}), .b ({signal_9181, signal_5913}), .clk (clk), .r (Fresh[423]), .c ({signal_9312, signal_6020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5785 ( .a ({signal_8424, signal_5141}), .b ({signal_9188, signal_5920}), .clk (clk), .r (Fresh[424]), .c ({signal_9313, signal_6021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5786 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_9187, signal_5919}), .clk (clk), .r (Fresh[425]), .c ({signal_9314, signal_6022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5787 ( .a ({signal_8170, signal_4896}), .b ({signal_9186, signal_5918}), .clk (clk), .r (Fresh[426]), .c ({signal_9315, signal_6023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5788 ( .a ({signal_8427, signal_5144}), .b ({signal_9185, signal_5917}), .clk (clk), .r (Fresh[427]), .c ({signal_9316, signal_6024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5789 ( .a ({signal_8429, signal_5146}), .b ({signal_9188, signal_5920}), .clk (clk), .r (Fresh[428]), .c ({signal_9317, signal_6025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5790 ( .a ({signal_8174, signal_4900}), .b ({signal_9187, signal_5919}), .clk (clk), .r (Fresh[429]), .c ({signal_9318, signal_6026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5791 ( .a ({signal_8175, signal_4901}), .b ({signal_9186, signal_5918}), .clk (clk), .r (Fresh[430]), .c ({signal_9319, signal_6027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5792 ( .a ({signal_8428, signal_5145}), .b ({signal_9185, signal_5917}), .clk (clk), .r (Fresh[431]), .c ({signal_9320, signal_6028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5793 ( .a ({signal_8073, signal_4689}), .b ({signal_9256, signal_5924}), .clk (clk), .r (Fresh[432]), .c ({signal_9469, signal_6029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5794 ( .a ({signal_8077, signal_4693}), .b ({signal_9255, signal_5923}), .clk (clk), .r (Fresh[433]), .c ({signal_9470, signal_6030}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5795 ( .a ({signal_8076, signal_4692}), .b ({signal_9254, signal_5922}), .clk (clk), .r (Fresh[434]), .c ({signal_9471, signal_6031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5796 ( .a ({signal_8272, signal_4904}), .b ({signal_9253, signal_5921}), .clk (clk), .r (Fresh[435]), .c ({signal_9472, signal_6032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5797 ( .a ({signal_8075, signal_4691}), .b ({signal_9256, signal_5924}), .clk (clk), .r (Fresh[436]), .c ({signal_9473, signal_6033}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5798 ( .a ({signal_7883, signal_4551}), .b ({signal_9255, signal_5923}), .clk (clk), .r (Fresh[437]), .c ({signal_9474, signal_6034}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5799 ( .a ({signal_7881, signal_4549}), .b ({signal_9254, signal_5922}), .clk (clk), .r (Fresh[438]), .c ({signal_9475, signal_6035}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5800 ( .a ({signal_7882, signal_4550}), .b ({signal_9253, signal_5921}), .clk (clk), .r (Fresh[439]), .c ({signal_9476, signal_6036}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5801 ( .a ({signal_8431, signal_5154}), .b ({signal_9192, signal_5928}), .clk (clk), .r (Fresh[440]), .c ({signal_9321, signal_6037}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5802 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_9191, signal_5927}), .clk (clk), .r (Fresh[441]), .c ({signal_9322, signal_6038}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5803 ( .a ({signal_8178, signal_4911}), .b ({signal_9190, signal_5926}), .clk (clk), .r (Fresh[442]), .c ({signal_9323, signal_6039}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5804 ( .a ({signal_8434, signal_5157}), .b ({signal_9189, signal_5925}), .clk (clk), .r (Fresh[443]), .c ({signal_9324, signal_6040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5805 ( .a ({signal_8436, signal_5159}), .b ({signal_9192, signal_5928}), .clk (clk), .r (Fresh[444]), .c ({signal_9325, signal_6041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5806 ( .a ({signal_8182, signal_4915}), .b ({signal_9191, signal_5927}), .clk (clk), .r (Fresh[445]), .c ({signal_9326, signal_6042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5807 ( .a ({signal_8183, signal_4916}), .b ({signal_9190, signal_5926}), .clk (clk), .r (Fresh[446]), .c ({signal_9327, signal_6043}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5808 ( .a ({signal_8435, signal_5158}), .b ({signal_9189, signal_5925}), .clk (clk), .r (Fresh[447]), .c ({signal_9328, signal_6044}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5809 ( .a ({signal_8438, signal_5161}), .b ({signal_9196, signal_5932}), .clk (clk), .r (Fresh[448]), .c ({signal_9329, signal_6045}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5810 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_9195, signal_5931}), .clk (clk), .r (Fresh[449]), .c ({signal_9330, signal_6046}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5811 ( .a ({signal_8186, signal_4919}), .b ({signal_9194, signal_5930}), .clk (clk), .r (Fresh[450]), .c ({signal_9331, signal_6047}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5812 ( .a ({signal_8441, signal_5164}), .b ({signal_9193, signal_5929}), .clk (clk), .r (Fresh[451]), .c ({signal_9332, signal_6048}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5813 ( .a ({signal_8443, signal_5166}), .b ({signal_9196, signal_5932}), .clk (clk), .r (Fresh[452]), .c ({signal_9333, signal_6049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5814 ( .a ({signal_8190, signal_4923}), .b ({signal_9195, signal_5931}), .clk (clk), .r (Fresh[453]), .c ({signal_9334, signal_6050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5815 ( .a ({signal_8191, signal_4924}), .b ({signal_9194, signal_5930}), .clk (clk), .r (Fresh[454]), .c ({signal_9335, signal_6051}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5816 ( .a ({signal_8442, signal_5165}), .b ({signal_9193, signal_5929}), .clk (clk), .r (Fresh[455]), .c ({signal_9336, signal_6052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5817 ( .a ({signal_8445, signal_5168}), .b ({signal_9200, signal_5936}), .clk (clk), .r (Fresh[456]), .c ({signal_9337, signal_6053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5818 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_9199, signal_5935}), .clk (clk), .r (Fresh[457]), .c ({signal_9338, signal_6054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5819 ( .a ({signal_8194, signal_4927}), .b ({signal_9198, signal_5934}), .clk (clk), .r (Fresh[458]), .c ({signal_9339, signal_6055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5820 ( .a ({signal_8448, signal_5171}), .b ({signal_9197, signal_5933}), .clk (clk), .r (Fresh[459]), .c ({signal_9340, signal_6056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5821 ( .a ({signal_8450, signal_5173}), .b ({signal_9200, signal_5936}), .clk (clk), .r (Fresh[460]), .c ({signal_9341, signal_6057}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5822 ( .a ({signal_8198, signal_4931}), .b ({signal_9199, signal_5935}), .clk (clk), .r (Fresh[461]), .c ({signal_9342, signal_6058}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5823 ( .a ({signal_8199, signal_4932}), .b ({signal_9198, signal_5934}), .clk (clk), .r (Fresh[462]), .c ({signal_9343, signal_6059}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5824 ( .a ({signal_8449, signal_5172}), .b ({signal_9197, signal_5933}), .clk (clk), .r (Fresh[463]), .c ({signal_9344, signal_6060}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5825 ( .a ({signal_8081, signal_4727}), .b ({signal_9260, signal_5940}), .clk (clk), .r (Fresh[464]), .c ({signal_9477, signal_6061}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5826 ( .a ({signal_8085, signal_4731}), .b ({signal_9259, signal_5939}), .clk (clk), .r (Fresh[465]), .c ({signal_9478, signal_6062}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5827 ( .a ({signal_8084, signal_4730}), .b ({signal_9258, signal_5938}), .clk (clk), .r (Fresh[466]), .c ({signal_9479, signal_6063}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5828 ( .a ({signal_8279, signal_4935}), .b ({signal_9257, signal_5937}), .clk (clk), .r (Fresh[467]), .c ({signal_9480, signal_6064}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5829 ( .a ({signal_8083, signal_4729}), .b ({signal_9260, signal_5940}), .clk (clk), .r (Fresh[468]), .c ({signal_9481, signal_6065}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5830 ( .a ({signal_7893, signal_4561}), .b ({signal_9259, signal_5939}), .clk (clk), .r (Fresh[469]), .c ({signal_9482, signal_6066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5831 ( .a ({signal_7891, signal_4559}), .b ({signal_9258, signal_5938}), .clk (clk), .r (Fresh[470]), .c ({signal_9483, signal_6067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5832 ( .a ({signal_7892, signal_4560}), .b ({signal_9257, signal_5937}), .clk (clk), .r (Fresh[471]), .c ({signal_9484, signal_6068}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5833 ( .a ({signal_8452, signal_5181}), .b ({signal_9204, signal_5944}), .clk (clk), .r (Fresh[472]), .c ({signal_9345, signal_6069}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5834 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_9203, signal_5943}), .clk (clk), .r (Fresh[473]), .c ({signal_9346, signal_6070}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5835 ( .a ({signal_8202, signal_4942}), .b ({signal_9202, signal_5942}), .clk (clk), .r (Fresh[474]), .c ({signal_9347, signal_6071}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5836 ( .a ({signal_8455, signal_5184}), .b ({signal_9201, signal_5941}), .clk (clk), .r (Fresh[475]), .c ({signal_9348, signal_6072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5837 ( .a ({signal_8457, signal_5186}), .b ({signal_9204, signal_5944}), .clk (clk), .r (Fresh[476]), .c ({signal_9349, signal_6073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5838 ( .a ({signal_8206, signal_4946}), .b ({signal_9203, signal_5943}), .clk (clk), .r (Fresh[477]), .c ({signal_9350, signal_6074}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5839 ( .a ({signal_8207, signal_4947}), .b ({signal_9202, signal_5942}), .clk (clk), .r (Fresh[478]), .c ({signal_9351, signal_6075}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5840 ( .a ({signal_8456, signal_5185}), .b ({signal_9201, signal_5941}), .clk (clk), .r (Fresh[479]), .c ({signal_9352, signal_6076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5841 ( .a ({signal_8459, signal_5188}), .b ({signal_9208, signal_5948}), .clk (clk), .r (Fresh[480]), .c ({signal_9353, signal_6077}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5842 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_9207, signal_5947}), .clk (clk), .r (Fresh[481]), .c ({signal_9354, signal_6078}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5843 ( .a ({signal_8210, signal_4950}), .b ({signal_9206, signal_5946}), .clk (clk), .r (Fresh[482]), .c ({signal_9355, signal_6079}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5844 ( .a ({signal_8462, signal_5191}), .b ({signal_9205, signal_5945}), .clk (clk), .r (Fresh[483]), .c ({signal_9356, signal_6080}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5845 ( .a ({signal_8464, signal_5193}), .b ({signal_9208, signal_5948}), .clk (clk), .r (Fresh[484]), .c ({signal_9357, signal_6081}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5846 ( .a ({signal_8214, signal_4954}), .b ({signal_9207, signal_5947}), .clk (clk), .r (Fresh[485]), .c ({signal_9358, signal_6082}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5847 ( .a ({signal_8215, signal_4955}), .b ({signal_9206, signal_5946}), .clk (clk), .r (Fresh[486]), .c ({signal_9359, signal_6083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5848 ( .a ({signal_8463, signal_5192}), .b ({signal_9205, signal_5945}), .clk (clk), .r (Fresh[487]), .c ({signal_9360, signal_6084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5849 ( .a ({signal_8466, signal_5195}), .b ({signal_9212, signal_5952}), .clk (clk), .r (Fresh[488]), .c ({signal_9361, signal_6085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5850 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_9211, signal_5951}), .clk (clk), .r (Fresh[489]), .c ({signal_9362, signal_6086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5851 ( .a ({signal_8218, signal_4958}), .b ({signal_9210, signal_5950}), .clk (clk), .r (Fresh[490]), .c ({signal_9363, signal_6087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5852 ( .a ({signal_8469, signal_5198}), .b ({signal_9209, signal_5949}), .clk (clk), .r (Fresh[491]), .c ({signal_9364, signal_6088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5853 ( .a ({signal_8471, signal_5200}), .b ({signal_9212, signal_5952}), .clk (clk), .r (Fresh[492]), .c ({signal_9365, signal_6089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5854 ( .a ({signal_8222, signal_4962}), .b ({signal_9211, signal_5951}), .clk (clk), .r (Fresh[493]), .c ({signal_9366, signal_6090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5855 ( .a ({signal_8223, signal_4963}), .b ({signal_9210, signal_5950}), .clk (clk), .r (Fresh[494]), .c ({signal_9367, signal_6091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5856 ( .a ({signal_8470, signal_5199}), .b ({signal_9209, signal_5949}), .clk (clk), .r (Fresh[495]), .c ({signal_9368, signal_6092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5857 ( .a ({signal_8089, signal_4765}), .b ({signal_9264, signal_5956}), .clk (clk), .r (Fresh[496]), .c ({signal_9485, signal_6093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5858 ( .a ({signal_8093, signal_4769}), .b ({signal_9263, signal_5955}), .clk (clk), .r (Fresh[497]), .c ({signal_9486, signal_6094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5859 ( .a ({signal_8092, signal_4768}), .b ({signal_9262, signal_5954}), .clk (clk), .r (Fresh[498]), .c ({signal_9487, signal_6095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5860 ( .a ({signal_8286, signal_4966}), .b ({signal_9261, signal_5953}), .clk (clk), .r (Fresh[499]), .c ({signal_9488, signal_6096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5861 ( .a ({signal_8091, signal_4767}), .b ({signal_9264, signal_5956}), .clk (clk), .r (Fresh[500]), .c ({signal_9489, signal_6097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5862 ( .a ({signal_7903, signal_4571}), .b ({signal_9263, signal_5955}), .clk (clk), .r (Fresh[501]), .c ({signal_9490, signal_6098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5863 ( .a ({signal_7901, signal_4569}), .b ({signal_9262, signal_5954}), .clk (clk), .r (Fresh[502]), .c ({signal_9491, signal_6099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5864 ( .a ({signal_7902, signal_4570}), .b ({signal_9261, signal_5953}), .clk (clk), .r (Fresh[503]), .c ({signal_9492, signal_6100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5865 ( .a ({signal_8041, signal_4773}), .b ({signal_9216, signal_5960}), .clk (clk), .r (Fresh[504]), .c ({signal_9369, signal_6101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5866 ( .a ({signal_8045, signal_4777}), .b ({signal_9215, signal_5959}), .clk (clk), .r (Fresh[505]), .c ({signal_9370, signal_6102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5867 ( .a ({signal_8044, signal_4776}), .b ({signal_9214, signal_5958}), .clk (clk), .r (Fresh[506]), .c ({signal_9371, signal_6103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5868 ( .a ({signal_8226, signal_4973}), .b ({signal_9213, signal_5957}), .clk (clk), .r (Fresh[507]), .c ({signal_9372, signal_6104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5869 ( .a ({signal_8043, signal_4775}), .b ({signal_9216, signal_5960}), .clk (clk), .r (Fresh[508]), .c ({signal_9373, signal_6105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5870 ( .a ({signal_7843, signal_4581}), .b ({signal_9215, signal_5959}), .clk (clk), .r (Fresh[509]), .c ({signal_9374, signal_6106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5871 ( .a ({signal_7841, signal_4579}), .b ({signal_9214, signal_5958}), .clk (clk), .r (Fresh[510]), .c ({signal_9375, signal_6107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5872 ( .a ({signal_7842, signal_4580}), .b ({signal_9213, signal_5957}), .clk (clk), .r (Fresh[511]), .c ({signal_9376, signal_6108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5873 ( .a ({signal_8049, signal_4781}), .b ({signal_9220, signal_5964}), .clk (clk), .r (Fresh[512]), .c ({signal_9377, signal_6109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5874 ( .a ({signal_8053, signal_4785}), .b ({signal_9219, signal_5963}), .clk (clk), .r (Fresh[513]), .c ({signal_9378, signal_6110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5875 ( .a ({signal_8052, signal_4784}), .b ({signal_9218, signal_5962}), .clk (clk), .r (Fresh[514]), .c ({signal_9379, signal_6111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5876 ( .a ({signal_8233, signal_4980}), .b ({signal_9217, signal_5961}), .clk (clk), .r (Fresh[515]), .c ({signal_9380, signal_6112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5877 ( .a ({signal_8051, signal_4783}), .b ({signal_9220, signal_5964}), .clk (clk), .r (Fresh[516]), .c ({signal_9381, signal_6113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5878 ( .a ({signal_7853, signal_4591}), .b ({signal_9219, signal_5963}), .clk (clk), .r (Fresh[517]), .c ({signal_9382, signal_6114}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5879 ( .a ({signal_7851, signal_4589}), .b ({signal_9218, signal_5962}), .clk (clk), .r (Fresh[518]), .c ({signal_9383, signal_6115}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5880 ( .a ({signal_7852, signal_4590}), .b ({signal_9217, signal_5961}), .clk (clk), .r (Fresh[519]), .c ({signal_9384, signal_6116}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5881 ( .a ({signal_8057, signal_4789}), .b ({signal_9224, signal_5968}), .clk (clk), .r (Fresh[520]), .c ({signal_9385, signal_6117}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5882 ( .a ({signal_8061, signal_4793}), .b ({signal_9223, signal_5967}), .clk (clk), .r (Fresh[521]), .c ({signal_9386, signal_6118}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5883 ( .a ({signal_8060, signal_4792}), .b ({signal_9222, signal_5966}), .clk (clk), .r (Fresh[522]), .c ({signal_9387, signal_6119}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5884 ( .a ({signal_8240, signal_4987}), .b ({signal_9221, signal_5965}), .clk (clk), .r (Fresh[523]), .c ({signal_9388, signal_6120}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5885 ( .a ({signal_8059, signal_4791}), .b ({signal_9224, signal_5968}), .clk (clk), .r (Fresh[524]), .c ({signal_9389, signal_6121}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5886 ( .a ({signal_7863, signal_4601}), .b ({signal_9223, signal_5967}), .clk (clk), .r (Fresh[525]), .c ({signal_9390, signal_6122}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5887 ( .a ({signal_7861, signal_4599}), .b ({signal_9222, signal_5966}), .clk (clk), .r (Fresh[526]), .c ({signal_9391, signal_6123}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5888 ( .a ({signal_7862, signal_4600}), .b ({signal_9221, signal_5965}), .clk (clk), .r (Fresh[527]), .c ({signal_9392, signal_6124}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5889 ( .a ({signal_8065, signal_4797}), .b ({signal_9228, signal_5972}), .clk (clk), .r (Fresh[528]), .c ({signal_9393, signal_6125}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5890 ( .a ({signal_8069, signal_4801}), .b ({signal_9227, signal_5971}), .clk (clk), .r (Fresh[529]), .c ({signal_9394, signal_6126}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5891 ( .a ({signal_8068, signal_4800}), .b ({signal_9226, signal_5970}), .clk (clk), .r (Fresh[530]), .c ({signal_9395, signal_6127}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5892 ( .a ({signal_8247, signal_4994}), .b ({signal_9225, signal_5969}), .clk (clk), .r (Fresh[531]), .c ({signal_9396, signal_6128}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5893 ( .a ({signal_8067, signal_4799}), .b ({signal_9228, signal_5972}), .clk (clk), .r (Fresh[532]), .c ({signal_9397, signal_6129}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5894 ( .a ({signal_7873, signal_4611}), .b ({signal_9227, signal_5971}), .clk (clk), .r (Fresh[533]), .c ({signal_9398, signal_6130}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5895 ( .a ({signal_7871, signal_4609}), .b ({signal_9226, signal_5970}), .clk (clk), .r (Fresh[534]), .c ({signal_9399, signal_6131}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5896 ( .a ({signal_7872, signal_4610}), .b ({signal_9225, signal_5969}), .clk (clk), .r (Fresh[535]), .c ({signal_9400, signal_6132}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5926 ( .a ({signal_9231, signal_5839}), .b ({signal_9233, signal_5841}), .c ({signal_9494, signal_6162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5927 ( .a ({signal_9232, signal_5840}), .b ({signal_9235, signal_5843}), .c ({signal_9495, signal_6163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5928 ( .a ({signal_9230, signal_5838}), .b ({signal_9232, signal_5840}), .c ({signal_9496, signal_6164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5942 ( .a ({signal_9239, signal_5847}), .b ({signal_9241, signal_5849}), .c ({signal_9498, signal_6178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5943 ( .a ({signal_9240, signal_5848}), .b ({signal_9243, signal_5851}), .c ({signal_9499, signal_6179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5944 ( .a ({signal_9238, signal_5846}), .b ({signal_9240, signal_5848}), .c ({signal_9500, signal_6180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5958 ( .a ({signal_9247, signal_5855}), .b ({signal_9249, signal_5857}), .c ({signal_9502, signal_6194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5959 ( .a ({signal_9248, signal_5856}), .b ({signal_9251, signal_5859}), .c ({signal_9503, signal_6195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5960 ( .a ({signal_9246, signal_5854}), .b ({signal_9248, signal_5856}), .c ({signal_9504, signal_6196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5962 ( .a ({signal_9131, signal_5863}), .b ({signal_9133, signal_5865}), .c ({signal_9454, signal_6198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5963 ( .a ({signal_9132, signal_5864}), .b ({signal_9135, signal_5867}), .c ({signal_9455, signal_6199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5964 ( .a ({signal_9130, signal_5862}), .b ({signal_9132, signal_5864}), .c ({signal_9456, signal_6200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5966 ( .a ({signal_9139, signal_5871}), .b ({signal_9141, signal_5873}), .c ({signal_9458, signal_6202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5967 ( .a ({signal_9140, signal_5872}), .b ({signal_9143, signal_5875}), .c ({signal_9459, signal_6203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5968 ( .a ({signal_9138, signal_5870}), .b ({signal_9140, signal_5872}), .c ({signal_9460, signal_6204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5970 ( .a ({signal_9147, signal_5879}), .b ({signal_9149, signal_5881}), .c ({signal_9462, signal_6206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5971 ( .a ({signal_9148, signal_5880}), .b ({signal_9151, signal_5883}), .c ({signal_9463, signal_6207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5972 ( .a ({signal_9146, signal_5878}), .b ({signal_9148, signal_5880}), .c ({signal_9464, signal_6208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5974 ( .a ({signal_9155, signal_5887}), .b ({signal_9157, signal_5889}), .c ({signal_9466, signal_6210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5975 ( .a ({signal_9156, signal_5888}), .b ({signal_9159, signal_5891}), .c ({signal_9467, signal_6211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_5976 ( .a ({signal_9154, signal_5886}), .b ({signal_9156, signal_5888}), .c ({signal_9468, signal_6212}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5977 ( .a ({signal_8121, signal_4847}), .b ({signal_9404, signal_6136}), .clk (clk), .r (Fresh[536]), .c ({signal_9505, signal_6213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5978 ( .a ({signal_8125, signal_4851}), .b ({signal_9403, signal_6135}), .clk (clk), .r (Fresh[537]), .c ({signal_9506, signal_6214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5979 ( .a ({signal_8124, signal_4850}), .b ({signal_9402, signal_6134}), .clk (clk), .r (Fresh[538]), .c ({signal_9507, signal_6215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5980 ( .a ({signal_8383, signal_5100}), .b ({signal_9401, signal_6133}), .clk (clk), .r (Fresh[539]), .c ({signal_9508, signal_6216}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5981 ( .a ({signal_8123, signal_4849}), .b ({signal_9404, signal_6136}), .clk (clk), .r (Fresh[540]), .c ({signal_9509, signal_6217}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5982 ( .a ({signal_7913, signal_4621}), .b ({signal_9403, signal_6135}), .clk (clk), .r (Fresh[541]), .c ({signal_9510, signal_6218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5983 ( .a ({signal_7911, signal_4619}), .b ({signal_9402, signal_6134}), .clk (clk), .r (Fresh[542]), .c ({signal_9511, signal_6219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5984 ( .a ({signal_7912, signal_4620}), .b ({signal_9401, signal_6133}), .clk (clk), .r (Fresh[543]), .c ({signal_9512, signal_6220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5985 ( .a ({signal_8129, signal_4855}), .b ({signal_9408, signal_6140}), .clk (clk), .r (Fresh[544]), .c ({signal_9513, signal_6221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5986 ( .a ({signal_8133, signal_4859}), .b ({signal_9407, signal_6139}), .clk (clk), .r (Fresh[545]), .c ({signal_9514, signal_6222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5987 ( .a ({signal_8132, signal_4858}), .b ({signal_9406, signal_6138}), .clk (clk), .r (Fresh[546]), .c ({signal_9515, signal_6223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5988 ( .a ({signal_8390, signal_5107}), .b ({signal_9405, signal_6137}), .clk (clk), .r (Fresh[547]), .c ({signal_9516, signal_6224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5989 ( .a ({signal_8131, signal_4857}), .b ({signal_9408, signal_6140}), .clk (clk), .r (Fresh[548]), .c ({signal_9517, signal_6225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5990 ( .a ({signal_7923, signal_4631}), .b ({signal_9407, signal_6139}), .clk (clk), .r (Fresh[549]), .c ({signal_9518, signal_6226}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5991 ( .a ({signal_7921, signal_4629}), .b ({signal_9406, signal_6138}), .clk (clk), .r (Fresh[550]), .c ({signal_9519, signal_6227}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5992 ( .a ({signal_7922, signal_4630}), .b ({signal_9405, signal_6137}), .clk (clk), .r (Fresh[551]), .c ({signal_9520, signal_6228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5993 ( .a ({signal_8137, signal_4863}), .b ({signal_9412, signal_6144}), .clk (clk), .r (Fresh[552]), .c ({signal_9521, signal_6229}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5994 ( .a ({signal_8141, signal_4867}), .b ({signal_9411, signal_6143}), .clk (clk), .r (Fresh[553]), .c ({signal_9522, signal_6230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5995 ( .a ({signal_8140, signal_4866}), .b ({signal_9410, signal_6142}), .clk (clk), .r (Fresh[554]), .c ({signal_9523, signal_6231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5996 ( .a ({signal_8397, signal_5114}), .b ({signal_9409, signal_6141}), .clk (clk), .r (Fresh[555]), .c ({signal_9524, signal_6232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5997 ( .a ({signal_8139, signal_4865}), .b ({signal_9412, signal_6144}), .clk (clk), .r (Fresh[556]), .c ({signal_9525, signal_6233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5998 ( .a ({signal_7933, signal_4641}), .b ({signal_9411, signal_6143}), .clk (clk), .r (Fresh[557]), .c ({signal_9526, signal_6234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_5999 ( .a ({signal_7931, signal_4639}), .b ({signal_9410, signal_6142}), .clk (clk), .r (Fresh[558]), .c ({signal_9527, signal_6235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6000 ( .a ({signal_7932, signal_4640}), .b ({signal_9409, signal_6141}), .clk (clk), .r (Fresh[559]), .c ({signal_9528, signal_6236}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6001 ( .a ({signal_8145, signal_4871}), .b ({signal_9416, signal_6148}), .clk (clk), .r (Fresh[560]), .c ({signal_9529, signal_6237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6002 ( .a ({signal_8149, signal_4875}), .b ({signal_9415, signal_6147}), .clk (clk), .r (Fresh[561]), .c ({signal_9530, signal_6238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6003 ( .a ({signal_8148, signal_4874}), .b ({signal_9414, signal_6146}), .clk (clk), .r (Fresh[562]), .c ({signal_9531, signal_6239}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6004 ( .a ({signal_8404, signal_5121}), .b ({signal_9413, signal_6145}), .clk (clk), .r (Fresh[563]), .c ({signal_9532, signal_6240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6005 ( .a ({signal_8147, signal_4873}), .b ({signal_9416, signal_6148}), .clk (clk), .r (Fresh[564]), .c ({signal_9533, signal_6241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6006 ( .a ({signal_7943, signal_4651}), .b ({signal_9415, signal_6147}), .clk (clk), .r (Fresh[565]), .c ({signal_9534, signal_6242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6007 ( .a ({signal_7941, signal_4649}), .b ({signal_9414, signal_6146}), .clk (clk), .r (Fresh[566]), .c ({signal_9535, signal_6243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6008 ( .a ({signal_7942, signal_4650}), .b ({signal_9413, signal_6145}), .clk (clk), .r (Fresh[567]), .c ({signal_9536, signal_6244}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6009 ( .a ({signal_8153, signal_4879}), .b ({signal_9420, signal_6152}), .clk (clk), .r (Fresh[568]), .c ({signal_9537, signal_6245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6010 ( .a ({signal_8157, signal_4883}), .b ({signal_9419, signal_6151}), .clk (clk), .r (Fresh[569]), .c ({signal_9538, signal_6246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6011 ( .a ({signal_8156, signal_4882}), .b ({signal_9418, signal_6150}), .clk (clk), .r (Fresh[570]), .c ({signal_9539, signal_6247}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6012 ( .a ({signal_8411, signal_5128}), .b ({signal_9417, signal_6149}), .clk (clk), .r (Fresh[571]), .c ({signal_9540, signal_6248}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6013 ( .a ({signal_8155, signal_4881}), .b ({signal_9420, signal_6152}), .clk (clk), .r (Fresh[572]), .c ({signal_9541, signal_6249}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6014 ( .a ({signal_7953, signal_4661}), .b ({signal_9419, signal_6151}), .clk (clk), .r (Fresh[573]), .c ({signal_9542, signal_6250}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6015 ( .a ({signal_7951, signal_4659}), .b ({signal_9418, signal_6150}), .clk (clk), .r (Fresh[574]), .c ({signal_9543, signal_6251}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6016 ( .a ({signal_7952, signal_4660}), .b ({signal_9417, signal_6149}), .clk (clk), .r (Fresh[575]), .c ({signal_9544, signal_6252}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6017 ( .a ({signal_8161, signal_4887}), .b ({signal_9424, signal_6156}), .clk (clk), .r (Fresh[576]), .c ({signal_9545, signal_6253}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6018 ( .a ({signal_8165, signal_4891}), .b ({signal_9423, signal_6155}), .clk (clk), .r (Fresh[577]), .c ({signal_9546, signal_6254}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6019 ( .a ({signal_8164, signal_4890}), .b ({signal_9422, signal_6154}), .clk (clk), .r (Fresh[578]), .c ({signal_9547, signal_6255}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6020 ( .a ({signal_8418, signal_5135}), .b ({signal_9421, signal_6153}), .clk (clk), .r (Fresh[579]), .c ({signal_9548, signal_6256}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6021 ( .a ({signal_8163, signal_4889}), .b ({signal_9424, signal_6156}), .clk (clk), .r (Fresh[580]), .c ({signal_9549, signal_6257}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6022 ( .a ({signal_7963, signal_4671}), .b ({signal_9423, signal_6155}), .clk (clk), .r (Fresh[581]), .c ({signal_9550, signal_6258}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6023 ( .a ({signal_7961, signal_4669}), .b ({signal_9422, signal_6154}), .clk (clk), .r (Fresh[582]), .c ({signal_9551, signal_6259}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6024 ( .a ({signal_7962, signal_4670}), .b ({signal_9421, signal_6153}), .clk (clk), .r (Fresh[583]), .c ({signal_9552, signal_6260}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6025 ( .a ({signal_8169, signal_4895}), .b ({signal_9428, signal_6160}), .clk (clk), .r (Fresh[584]), .c ({signal_9553, signal_6261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6026 ( .a ({signal_8173, signal_4899}), .b ({signal_9427, signal_6159}), .clk (clk), .r (Fresh[585]), .c ({signal_9554, signal_6262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6027 ( .a ({signal_8172, signal_4898}), .b ({signal_9426, signal_6158}), .clk (clk), .r (Fresh[586]), .c ({signal_9555, signal_6263}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6028 ( .a ({signal_8425, signal_5142}), .b ({signal_9425, signal_6157}), .clk (clk), .r (Fresh[587]), .c ({signal_9556, signal_6264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6029 ( .a ({signal_8171, signal_4897}), .b ({signal_9428, signal_6160}), .clk (clk), .r (Fresh[588]), .c ({signal_9557, signal_6265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6030 ( .a ({signal_7973, signal_4681}), .b ({signal_9427, signal_6159}), .clk (clk), .r (Fresh[589]), .c ({signal_9558, signal_6266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6031 ( .a ({signal_7971, signal_4679}), .b ({signal_9426, signal_6158}), .clk (clk), .r (Fresh[590]), .c ({signal_9559, signal_6267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6032 ( .a ({signal_7972, signal_4680}), .b ({signal_9425, signal_6157}), .clk (clk), .r (Fresh[591]), .c ({signal_9560, signal_6268}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6033 ( .a ({signal_8080, signal_4696}), .b ({signal_9493, signal_6161}), .clk (clk), .r (Fresh[592]), .c ({signal_9701, signal_6269}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6034 ( .a ({signal_7884, signal_4552}), .b ({signal_9493, signal_6161}), .clk (clk), .r (Fresh[593]), .c ({signal_9702, signal_6270}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6035 ( .a ({signal_8177, signal_4910}), .b ({signal_9432, signal_6168}), .clk (clk), .r (Fresh[594]), .c ({signal_9561, signal_6271}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6036 ( .a ({signal_8181, signal_4914}), .b ({signal_9431, signal_6167}), .clk (clk), .r (Fresh[595]), .c ({signal_9562, signal_6272}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6037 ( .a ({signal_8180, signal_4913}), .b ({signal_9430, signal_6166}), .clk (clk), .r (Fresh[596]), .c ({signal_9563, signal_6273}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6038 ( .a ({signal_8432, signal_5155}), .b ({signal_9429, signal_6165}), .clk (clk), .r (Fresh[597]), .c ({signal_9564, signal_6274}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6039 ( .a ({signal_8179, signal_4912}), .b ({signal_9432, signal_6168}), .clk (clk), .r (Fresh[598]), .c ({signal_9565, signal_6275}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6040 ( .a ({signal_7983, signal_4699}), .b ({signal_9431, signal_6167}), .clk (clk), .r (Fresh[599]), .c ({signal_9566, signal_6276}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6041 ( .a ({signal_7981, signal_4697}), .b ({signal_9430, signal_6166}), .clk (clk), .r (Fresh[600]), .c ({signal_9567, signal_6277}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6042 ( .a ({signal_7982, signal_4698}), .b ({signal_9429, signal_6165}), .clk (clk), .r (Fresh[601]), .c ({signal_9568, signal_6278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6043 ( .a ({signal_8185, signal_4918}), .b ({signal_9436, signal_6172}), .clk (clk), .r (Fresh[602]), .c ({signal_9569, signal_6279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6044 ( .a ({signal_8189, signal_4922}), .b ({signal_9435, signal_6171}), .clk (clk), .r (Fresh[603]), .c ({signal_9570, signal_6280}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6045 ( .a ({signal_8188, signal_4921}), .b ({signal_9434, signal_6170}), .clk (clk), .r (Fresh[604]), .c ({signal_9571, signal_6281}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6046 ( .a ({signal_8439, signal_5162}), .b ({signal_9433, signal_6169}), .clk (clk), .r (Fresh[605]), .c ({signal_9572, signal_6282}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6047 ( .a ({signal_8187, signal_4920}), .b ({signal_9436, signal_6172}), .clk (clk), .r (Fresh[606]), .c ({signal_9573, signal_6283}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6048 ( .a ({signal_7993, signal_4709}), .b ({signal_9435, signal_6171}), .clk (clk), .r (Fresh[607]), .c ({signal_9574, signal_6284}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6049 ( .a ({signal_7991, signal_4707}), .b ({signal_9434, signal_6170}), .clk (clk), .r (Fresh[608]), .c ({signal_9575, signal_6285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6050 ( .a ({signal_7992, signal_4708}), .b ({signal_9433, signal_6169}), .clk (clk), .r (Fresh[609]), .c ({signal_9576, signal_6286}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6051 ( .a ({signal_8193, signal_4926}), .b ({signal_9440, signal_6176}), .clk (clk), .r (Fresh[610]), .c ({signal_9577, signal_6287}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6052 ( .a ({signal_8197, signal_4930}), .b ({signal_9439, signal_6175}), .clk (clk), .r (Fresh[611]), .c ({signal_9578, signal_6288}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6053 ( .a ({signal_8196, signal_4929}), .b ({signal_9438, signal_6174}), .clk (clk), .r (Fresh[612]), .c ({signal_9579, signal_6289}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6054 ( .a ({signal_8446, signal_5169}), .b ({signal_9437, signal_6173}), .clk (clk), .r (Fresh[613]), .c ({signal_9580, signal_6290}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6055 ( .a ({signal_8195, signal_4928}), .b ({signal_9440, signal_6176}), .clk (clk), .r (Fresh[614]), .c ({signal_9581, signal_6291}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6056 ( .a ({signal_8003, signal_4719}), .b ({signal_9439, signal_6175}), .clk (clk), .r (Fresh[615]), .c ({signal_9582, signal_6292}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6057 ( .a ({signal_8001, signal_4717}), .b ({signal_9438, signal_6174}), .clk (clk), .r (Fresh[616]), .c ({signal_9583, signal_6293}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6058 ( .a ({signal_8002, signal_4718}), .b ({signal_9437, signal_6173}), .clk (clk), .r (Fresh[617]), .c ({signal_9584, signal_6294}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6059 ( .a ({signal_8088, signal_4734}), .b ({signal_9497, signal_6177}), .clk (clk), .r (Fresh[618]), .c ({signal_9703, signal_6295}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6060 ( .a ({signal_7894, signal_4562}), .b ({signal_9497, signal_6177}), .clk (clk), .r (Fresh[619]), .c ({signal_9704, signal_6296}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6061 ( .a ({signal_8201, signal_4941}), .b ({signal_9444, signal_6184}), .clk (clk), .r (Fresh[620]), .c ({signal_9585, signal_6297}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6062 ( .a ({signal_8205, signal_4945}), .b ({signal_9443, signal_6183}), .clk (clk), .r (Fresh[621]), .c ({signal_9586, signal_6298}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6063 ( .a ({signal_8204, signal_4944}), .b ({signal_9442, signal_6182}), .clk (clk), .r (Fresh[622]), .c ({signal_9587, signal_6299}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6064 ( .a ({signal_8453, signal_5182}), .b ({signal_9441, signal_6181}), .clk (clk), .r (Fresh[623]), .c ({signal_9588, signal_6300}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6065 ( .a ({signal_8203, signal_4943}), .b ({signal_9444, signal_6184}), .clk (clk), .r (Fresh[624]), .c ({signal_9589, signal_6301}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6066 ( .a ({signal_8013, signal_4737}), .b ({signal_9443, signal_6183}), .clk (clk), .r (Fresh[625]), .c ({signal_9590, signal_6302}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6067 ( .a ({signal_8011, signal_4735}), .b ({signal_9442, signal_6182}), .clk (clk), .r (Fresh[626]), .c ({signal_9591, signal_6303}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6068 ( .a ({signal_8012, signal_4736}), .b ({signal_9441, signal_6181}), .clk (clk), .r (Fresh[627]), .c ({signal_9592, signal_6304}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6069 ( .a ({signal_8209, signal_4949}), .b ({signal_9448, signal_6188}), .clk (clk), .r (Fresh[628]), .c ({signal_9593, signal_6305}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6070 ( .a ({signal_8213, signal_4953}), .b ({signal_9447, signal_6187}), .clk (clk), .r (Fresh[629]), .c ({signal_9594, signal_6306}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6071 ( .a ({signal_8212, signal_4952}), .b ({signal_9446, signal_6186}), .clk (clk), .r (Fresh[630]), .c ({signal_9595, signal_6307}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6072 ( .a ({signal_8460, signal_5189}), .b ({signal_9445, signal_6185}), .clk (clk), .r (Fresh[631]), .c ({signal_9596, signal_6308}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6073 ( .a ({signal_8211, signal_4951}), .b ({signal_9448, signal_6188}), .clk (clk), .r (Fresh[632]), .c ({signal_9597, signal_6309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6074 ( .a ({signal_8023, signal_4747}), .b ({signal_9447, signal_6187}), .clk (clk), .r (Fresh[633]), .c ({signal_9598, signal_6310}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6075 ( .a ({signal_8021, signal_4745}), .b ({signal_9446, signal_6186}), .clk (clk), .r (Fresh[634]), .c ({signal_9599, signal_6311}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6076 ( .a ({signal_8022, signal_4746}), .b ({signal_9445, signal_6185}), .clk (clk), .r (Fresh[635]), .c ({signal_9600, signal_6312}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6077 ( .a ({signal_8217, signal_4957}), .b ({signal_9452, signal_6192}), .clk (clk), .r (Fresh[636]), .c ({signal_9601, signal_6313}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6078 ( .a ({signal_8221, signal_4961}), .b ({signal_9451, signal_6191}), .clk (clk), .r (Fresh[637]), .c ({signal_9602, signal_6314}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6079 ( .a ({signal_8220, signal_4960}), .b ({signal_9450, signal_6190}), .clk (clk), .r (Fresh[638]), .c ({signal_9603, signal_6315}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6080 ( .a ({signal_8467, signal_5196}), .b ({signal_9449, signal_6189}), .clk (clk), .r (Fresh[639]), .c ({signal_9604, signal_6316}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6081 ( .a ({signal_8219, signal_4959}), .b ({signal_9452, signal_6192}), .clk (clk), .r (Fresh[640]), .c ({signal_9605, signal_6317}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6082 ( .a ({signal_8033, signal_4757}), .b ({signal_9451, signal_6191}), .clk (clk), .r (Fresh[641]), .c ({signal_9606, signal_6318}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6083 ( .a ({signal_8031, signal_4755}), .b ({signal_9450, signal_6190}), .clk (clk), .r (Fresh[642]), .c ({signal_9607, signal_6319}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6084 ( .a ({signal_8032, signal_4756}), .b ({signal_9449, signal_6189}), .clk (clk), .r (Fresh[643]), .c ({signal_9608, signal_6320}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6085 ( .a ({signal_8096, signal_4772}), .b ({signal_9501, signal_6193}), .clk (clk), .r (Fresh[644]), .c ({signal_9705, signal_6321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6086 ( .a ({signal_7904, signal_4572}), .b ({signal_9501, signal_6193}), .clk (clk), .r (Fresh[645]), .c ({signal_9706, signal_6322}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6087 ( .a ({signal_8048, signal_4780}), .b ({signal_9453, signal_6197}), .clk (clk), .r (Fresh[646]), .c ({signal_9609, signal_6323}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6088 ( .a ({signal_7844, signal_4582}), .b ({signal_9453, signal_6197}), .clk (clk), .r (Fresh[647]), .c ({signal_9610, signal_6324}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6089 ( .a ({signal_8056, signal_4788}), .b ({signal_9457, signal_6201}), .clk (clk), .r (Fresh[648]), .c ({signal_9611, signal_6325}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6090 ( .a ({signal_7854, signal_4592}), .b ({signal_9457, signal_6201}), .clk (clk), .r (Fresh[649]), .c ({signal_9612, signal_6326}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6091 ( .a ({signal_8064, signal_4796}), .b ({signal_9461, signal_6205}), .clk (clk), .r (Fresh[650]), .c ({signal_9613, signal_6327}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6092 ( .a ({signal_7864, signal_4602}), .b ({signal_9461, signal_6205}), .clk (clk), .r (Fresh[651]), .c ({signal_9614, signal_6328}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6093 ( .a ({signal_8072, signal_4804}), .b ({signal_9465, signal_6209}), .clk (clk), .r (Fresh[652]), .c ({signal_9615, signal_6329}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6094 ( .a ({signal_7874, signal_4612}), .b ({signal_9465, signal_6209}), .clk (clk), .r (Fresh[653]), .c ({signal_9616, signal_6330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6096 ( .a ({signal_9267, signal_5975}), .b ({signal_9269, signal_5977}), .c ({signal_9618, signal_6332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6097 ( .a ({signal_9268, signal_5976}), .b ({signal_9271, signal_5979}), .c ({signal_9619, signal_6333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6098 ( .a ({signal_9266, signal_5974}), .b ({signal_9268, signal_5976}), .c ({signal_9620, signal_6334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6100 ( .a ({signal_9275, signal_5983}), .b ({signal_9277, signal_5985}), .c ({signal_9622, signal_6336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6101 ( .a ({signal_9276, signal_5984}), .b ({signal_9279, signal_5987}), .c ({signal_9623, signal_6337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6102 ( .a ({signal_9274, signal_5982}), .b ({signal_9276, signal_5984}), .c ({signal_9624, signal_6338}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6104 ( .a ({signal_9283, signal_5991}), .b ({signal_9285, signal_5993}), .c ({signal_9626, signal_6340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6105 ( .a ({signal_9284, signal_5992}), .b ({signal_9287, signal_5995}), .c ({signal_9627, signal_6341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6106 ( .a ({signal_9282, signal_5990}), .b ({signal_9284, signal_5992}), .c ({signal_9628, signal_6342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6108 ( .a ({signal_9291, signal_5999}), .b ({signal_9293, signal_6001}), .c ({signal_9630, signal_6344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6109 ( .a ({signal_9292, signal_6000}), .b ({signal_9295, signal_6003}), .c ({signal_9631, signal_6345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6110 ( .a ({signal_9290, signal_5998}), .b ({signal_9292, signal_6000}), .c ({signal_9632, signal_6346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6112 ( .a ({signal_9299, signal_6007}), .b ({signal_9301, signal_6009}), .c ({signal_9634, signal_6348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6113 ( .a ({signal_9300, signal_6008}), .b ({signal_9303, signal_6011}), .c ({signal_9635, signal_6349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6114 ( .a ({signal_9298, signal_6006}), .b ({signal_9300, signal_6008}), .c ({signal_9636, signal_6350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6116 ( .a ({signal_9307, signal_6015}), .b ({signal_9309, signal_6017}), .c ({signal_9638, signal_6352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6117 ( .a ({signal_9308, signal_6016}), .b ({signal_9311, signal_6019}), .c ({signal_9639, signal_6353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6118 ( .a ({signal_9306, signal_6014}), .b ({signal_9308, signal_6016}), .c ({signal_9640, signal_6354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6120 ( .a ({signal_9315, signal_6023}), .b ({signal_9317, signal_6025}), .c ({signal_9642, signal_6356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6121 ( .a ({signal_9316, signal_6024}), .b ({signal_9319, signal_6027}), .c ({signal_9643, signal_6357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6122 ( .a ({signal_9314, signal_6022}), .b ({signal_9316, signal_6024}), .c ({signal_9644, signal_6358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6123 ( .a ({signal_9230, signal_5838}), .b ({signal_9469, signal_6029}), .c ({signal_9707, signal_6359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6124 ( .a ({signal_9229, signal_5837}), .b ({signal_9473, signal_6033}), .c ({signal_9708, signal_6360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6125 ( .a ({signal_9472, signal_6032}), .b ({signal_9474, signal_6034}), .c ({signal_9709, signal_6361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6126 ( .a ({signal_9470, signal_6030}), .b ({signal_9475, signal_6035}), .c ({signal_9710, signal_6362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6127 ( .a ({signal_9471, signal_6031}), .b ({signal_9475, signal_6035}), .c ({signal_9711, signal_6363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6128 ( .a ({signal_9473, signal_6033}), .b ({signal_9494, signal_6162}), .c ({signal_9712, signal_6364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6129 ( .a ({signal_9234, signal_5842}), .b ({signal_9494, signal_6162}), .c ({signal_9713, signal_6365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6130 ( .a ({signal_9474, signal_6034}), .b ({signal_9495, signal_6163}), .c ({signal_9714, signal_6366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6132 ( .a ({signal_9323, signal_6039}), .b ({signal_9325, signal_6041}), .c ({signal_9646, signal_6368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6133 ( .a ({signal_9324, signal_6040}), .b ({signal_9327, signal_6043}), .c ({signal_9647, signal_6369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6134 ( .a ({signal_9322, signal_6038}), .b ({signal_9324, signal_6040}), .c ({signal_9648, signal_6370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6136 ( .a ({signal_9331, signal_6047}), .b ({signal_9333, signal_6049}), .c ({signal_9650, signal_6372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6137 ( .a ({signal_9332, signal_6048}), .b ({signal_9335, signal_6051}), .c ({signal_9651, signal_6373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6138 ( .a ({signal_9330, signal_6046}), .b ({signal_9332, signal_6048}), .c ({signal_9652, signal_6374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6140 ( .a ({signal_9339, signal_6055}), .b ({signal_9341, signal_6057}), .c ({signal_9654, signal_6376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6141 ( .a ({signal_9340, signal_6056}), .b ({signal_9343, signal_6059}), .c ({signal_9655, signal_6377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6142 ( .a ({signal_9338, signal_6054}), .b ({signal_9340, signal_6056}), .c ({signal_9656, signal_6378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6143 ( .a ({signal_9238, signal_5846}), .b ({signal_9477, signal_6061}), .c ({signal_9715, signal_6379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6144 ( .a ({signal_9237, signal_5845}), .b ({signal_9481, signal_6065}), .c ({signal_9716, signal_6380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6145 ( .a ({signal_9480, signal_6064}), .b ({signal_9482, signal_6066}), .c ({signal_9717, signal_6381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6146 ( .a ({signal_9478, signal_6062}), .b ({signal_9483, signal_6067}), .c ({signal_9718, signal_6382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6147 ( .a ({signal_9479, signal_6063}), .b ({signal_9483, signal_6067}), .c ({signal_9719, signal_6383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6148 ( .a ({signal_9481, signal_6065}), .b ({signal_9498, signal_6178}), .c ({signal_9720, signal_6384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6149 ( .a ({signal_9242, signal_5850}), .b ({signal_9498, signal_6178}), .c ({signal_9721, signal_6385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6150 ( .a ({signal_9482, signal_6066}), .b ({signal_9499, signal_6179}), .c ({signal_9722, signal_6386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6152 ( .a ({signal_9347, signal_6071}), .b ({signal_9349, signal_6073}), .c ({signal_9658, signal_6388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6153 ( .a ({signal_9348, signal_6072}), .b ({signal_9351, signal_6075}), .c ({signal_9659, signal_6389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6154 ( .a ({signal_9346, signal_6070}), .b ({signal_9348, signal_6072}), .c ({signal_9660, signal_6390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6156 ( .a ({signal_9355, signal_6079}), .b ({signal_9357, signal_6081}), .c ({signal_9662, signal_6392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6157 ( .a ({signal_9356, signal_6080}), .b ({signal_9359, signal_6083}), .c ({signal_9663, signal_6393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6158 ( .a ({signal_9354, signal_6078}), .b ({signal_9356, signal_6080}), .c ({signal_9664, signal_6394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6160 ( .a ({signal_9363, signal_6087}), .b ({signal_9365, signal_6089}), .c ({signal_9666, signal_6396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6161 ( .a ({signal_9364, signal_6088}), .b ({signal_9367, signal_6091}), .c ({signal_9667, signal_6397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6162 ( .a ({signal_9362, signal_6086}), .b ({signal_9364, signal_6088}), .c ({signal_9668, signal_6398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6163 ( .a ({signal_9246, signal_5854}), .b ({signal_9485, signal_6093}), .c ({signal_9723, signal_6399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6164 ( .a ({signal_9245, signal_5853}), .b ({signal_9489, signal_6097}), .c ({signal_9724, signal_6400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6165 ( .a ({signal_9488, signal_6096}), .b ({signal_9490, signal_6098}), .c ({signal_9725, signal_6401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6166 ( .a ({signal_9486, signal_6094}), .b ({signal_9491, signal_6099}), .c ({signal_9726, signal_6402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6167 ( .a ({signal_9487, signal_6095}), .b ({signal_9491, signal_6099}), .c ({signal_9727, signal_6403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6168 ( .a ({signal_9489, signal_6097}), .b ({signal_9502, signal_6194}), .c ({signal_9728, signal_6404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6169 ( .a ({signal_9250, signal_5858}), .b ({signal_9502, signal_6194}), .c ({signal_9729, signal_6405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6170 ( .a ({signal_9490, signal_6098}), .b ({signal_9503, signal_6195}), .c ({signal_9730, signal_6406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6171 ( .a ({signal_9130, signal_5862}), .b ({signal_9369, signal_6101}), .c ({signal_9669, signal_6407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6172 ( .a ({signal_9129, signal_5861}), .b ({signal_9373, signal_6105}), .c ({signal_9670, signal_6408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6173 ( .a ({signal_9372, signal_6104}), .b ({signal_9374, signal_6106}), .c ({signal_9671, signal_6409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6174 ( .a ({signal_9370, signal_6102}), .b ({signal_9375, signal_6107}), .c ({signal_9672, signal_6410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6175 ( .a ({signal_9371, signal_6103}), .b ({signal_9375, signal_6107}), .c ({signal_9673, signal_6411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6176 ( .a ({signal_9373, signal_6105}), .b ({signal_9454, signal_6198}), .c ({signal_9674, signal_6412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6177 ( .a ({signal_9134, signal_5866}), .b ({signal_9454, signal_6198}), .c ({signal_9675, signal_6413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6178 ( .a ({signal_9374, signal_6106}), .b ({signal_9455, signal_6199}), .c ({signal_9676, signal_6414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6179 ( .a ({signal_9138, signal_5870}), .b ({signal_9377, signal_6109}), .c ({signal_9677, signal_6415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6180 ( .a ({signal_9137, signal_5869}), .b ({signal_9381, signal_6113}), .c ({signal_9678, signal_6416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6181 ( .a ({signal_9380, signal_6112}), .b ({signal_9382, signal_6114}), .c ({signal_9679, signal_6417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6182 ( .a ({signal_9378, signal_6110}), .b ({signal_9383, signal_6115}), .c ({signal_9680, signal_6418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6183 ( .a ({signal_9379, signal_6111}), .b ({signal_9383, signal_6115}), .c ({signal_9681, signal_6419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6184 ( .a ({signal_9381, signal_6113}), .b ({signal_9458, signal_6202}), .c ({signal_9682, signal_6420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6185 ( .a ({signal_9142, signal_5874}), .b ({signal_9458, signal_6202}), .c ({signal_9683, signal_6421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6186 ( .a ({signal_9382, signal_6114}), .b ({signal_9459, signal_6203}), .c ({signal_9684, signal_6422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6187 ( .a ({signal_9146, signal_5878}), .b ({signal_9385, signal_6117}), .c ({signal_9685, signal_6423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6188 ( .a ({signal_9145, signal_5877}), .b ({signal_9389, signal_6121}), .c ({signal_9686, signal_6424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6189 ( .a ({signal_9388, signal_6120}), .b ({signal_9390, signal_6122}), .c ({signal_9687, signal_6425}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6190 ( .a ({signal_9386, signal_6118}), .b ({signal_9391, signal_6123}), .c ({signal_9688, signal_6426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6191 ( .a ({signal_9387, signal_6119}), .b ({signal_9391, signal_6123}), .c ({signal_9689, signal_6427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6192 ( .a ({signal_9389, signal_6121}), .b ({signal_9462, signal_6206}), .c ({signal_9690, signal_6428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6193 ( .a ({signal_9150, signal_5882}), .b ({signal_9462, signal_6206}), .c ({signal_9691, signal_6429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6194 ( .a ({signal_9390, signal_6122}), .b ({signal_9463, signal_6207}), .c ({signal_9692, signal_6430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6195 ( .a ({signal_9154, signal_5886}), .b ({signal_9393, signal_6125}), .c ({signal_9693, signal_6431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6196 ( .a ({signal_9153, signal_5885}), .b ({signal_9397, signal_6129}), .c ({signal_9694, signal_6432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6197 ( .a ({signal_9396, signal_6128}), .b ({signal_9398, signal_6130}), .c ({signal_9695, signal_6433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6198 ( .a ({signal_9394, signal_6126}), .b ({signal_9399, signal_6131}), .c ({signal_9696, signal_6434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6199 ( .a ({signal_9395, signal_6127}), .b ({signal_9399, signal_6131}), .c ({signal_9697, signal_6435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6200 ( .a ({signal_9397, signal_6129}), .b ({signal_9466, signal_6210}), .c ({signal_9698, signal_6436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6201 ( .a ({signal_9158, signal_5890}), .b ({signal_9466, signal_6210}), .c ({signal_9699, signal_6437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6202 ( .a ({signal_9398, signal_6130}), .b ({signal_9467, signal_6211}), .c ({signal_9700, signal_6438}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6203 ( .a ({signal_8128, signal_4854}), .b ({signal_9617, signal_6331}), .clk (clk), .r (Fresh[654]), .c ({signal_9731, signal_6439}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6204 ( .a ({signal_7914, signal_4622}), .b ({signal_9617, signal_6331}), .clk (clk), .r (Fresh[655]), .c ({signal_9732, signal_6440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6205 ( .a ({signal_8136, signal_4862}), .b ({signal_9621, signal_6335}), .clk (clk), .r (Fresh[656]), .c ({signal_9733, signal_6441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6206 ( .a ({signal_7924, signal_4632}), .b ({signal_9621, signal_6335}), .clk (clk), .r (Fresh[657]), .c ({signal_9734, signal_6442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6207 ( .a ({signal_8144, signal_4870}), .b ({signal_9625, signal_6339}), .clk (clk), .r (Fresh[658]), .c ({signal_9735, signal_6443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6208 ( .a ({signal_7934, signal_4642}), .b ({signal_9625, signal_6339}), .clk (clk), .r (Fresh[659]), .c ({signal_9736, signal_6444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6209 ( .a ({signal_8152, signal_4878}), .b ({signal_9629, signal_6343}), .clk (clk), .r (Fresh[660]), .c ({signal_9737, signal_6445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6210 ( .a ({signal_7944, signal_4652}), .b ({signal_9629, signal_6343}), .clk (clk), .r (Fresh[661]), .c ({signal_9738, signal_6446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6211 ( .a ({signal_8160, signal_4886}), .b ({signal_9633, signal_6347}), .clk (clk), .r (Fresh[662]), .c ({signal_9739, signal_6447}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6212 ( .a ({signal_7954, signal_4662}), .b ({signal_9633, signal_6347}), .clk (clk), .r (Fresh[663]), .c ({signal_9740, signal_6448}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6213 ( .a ({signal_8168, signal_4894}), .b ({signal_9637, signal_6351}), .clk (clk), .r (Fresh[664]), .c ({signal_9741, signal_6449}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6214 ( .a ({signal_7964, signal_4672}), .b ({signal_9637, signal_6351}), .clk (clk), .r (Fresh[665]), .c ({signal_9742, signal_6450}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6215 ( .a ({signal_8176, signal_4902}), .b ({signal_9641, signal_6355}), .clk (clk), .r (Fresh[666]), .c ({signal_9743, signal_6451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6216 ( .a ({signal_7974, signal_4682}), .b ({signal_9641, signal_6355}), .clk (clk), .r (Fresh[667]), .c ({signal_9744, signal_6452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6217 ( .a ({signal_8184, signal_4917}), .b ({signal_9645, signal_6367}), .clk (clk), .r (Fresh[668]), .c ({signal_9745, signal_6453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6218 ( .a ({signal_7984, signal_4700}), .b ({signal_9645, signal_6367}), .clk (clk), .r (Fresh[669]), .c ({signal_9746, signal_6454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6219 ( .a ({signal_8192, signal_4925}), .b ({signal_9649, signal_6371}), .clk (clk), .r (Fresh[670]), .c ({signal_9747, signal_6455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6220 ( .a ({signal_7994, signal_4710}), .b ({signal_9649, signal_6371}), .clk (clk), .r (Fresh[671]), .c ({signal_9748, signal_6456}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6221 ( .a ({signal_8200, signal_4933}), .b ({signal_9653, signal_6375}), .clk (clk), .r (Fresh[672]), .c ({signal_9749, signal_6457}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6222 ( .a ({signal_8004, signal_4720}), .b ({signal_9653, signal_6375}), .clk (clk), .r (Fresh[673]), .c ({signal_9750, signal_6458}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6223 ( .a ({signal_8208, signal_4948}), .b ({signal_9657, signal_6387}), .clk (clk), .r (Fresh[674]), .c ({signal_9751, signal_6459}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6224 ( .a ({signal_8014, signal_4738}), .b ({signal_9657, signal_6387}), .clk (clk), .r (Fresh[675]), .c ({signal_9752, signal_6460}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6225 ( .a ({signal_8216, signal_4956}), .b ({signal_9661, signal_6391}), .clk (clk), .r (Fresh[676]), .c ({signal_9753, signal_6461}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6226 ( .a ({signal_8024, signal_4748}), .b ({signal_9661, signal_6391}), .clk (clk), .r (Fresh[677]), .c ({signal_9754, signal_6462}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6227 ( .a ({signal_8224, signal_4964}), .b ({signal_9665, signal_6395}), .clk (clk), .r (Fresh[678]), .c ({signal_9755, signal_6463}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_6228 ( .a ({signal_8034, signal_4758}), .b ({signal_9665, signal_6395}), .clk (clk), .r (Fresh[679]), .c ({signal_9756, signal_6464}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6229 ( .a ({signal_9266, signal_5974}), .b ({signal_9505, signal_6213}), .c ({signal_9757, signal_6465}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6230 ( .a ({signal_9265, signal_5973}), .b ({signal_9509, signal_6217}), .c ({signal_9758, signal_6466}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6231 ( .a ({signal_9508, signal_6216}), .b ({signal_9510, signal_6218}), .c ({signal_9759, signal_6467}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6232 ( .a ({signal_9506, signal_6214}), .b ({signal_9511, signal_6219}), .c ({signal_9760, signal_6468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6233 ( .a ({signal_9507, signal_6215}), .b ({signal_9511, signal_6219}), .c ({signal_9761, signal_6469}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6234 ( .a ({signal_9509, signal_6217}), .b ({signal_9618, signal_6332}), .c ({signal_9762, signal_6470}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6235 ( .a ({signal_9270, signal_5978}), .b ({signal_9618, signal_6332}), .c ({signal_9763, signal_6471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6236 ( .a ({signal_9510, signal_6218}), .b ({signal_9619, signal_6333}), .c ({signal_9764, signal_6472}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6237 ( .a ({signal_9274, signal_5982}), .b ({signal_9513, signal_6221}), .c ({signal_9765, signal_6473}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6238 ( .a ({signal_9273, signal_5981}), .b ({signal_9517, signal_6225}), .c ({signal_9766, signal_6474}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6239 ( .a ({signal_9516, signal_6224}), .b ({signal_9518, signal_6226}), .c ({signal_9767, signal_6475}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6240 ( .a ({signal_9514, signal_6222}), .b ({signal_9519, signal_6227}), .c ({signal_9768, signal_6476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6241 ( .a ({signal_9515, signal_6223}), .b ({signal_9519, signal_6227}), .c ({signal_9769, signal_6477}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6242 ( .a ({signal_9517, signal_6225}), .b ({signal_9622, signal_6336}), .c ({signal_9770, signal_6478}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6243 ( .a ({signal_9278, signal_5986}), .b ({signal_9622, signal_6336}), .c ({signal_9771, signal_6479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6244 ( .a ({signal_9518, signal_6226}), .b ({signal_9623, signal_6337}), .c ({signal_9772, signal_6480}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6245 ( .a ({signal_9282, signal_5990}), .b ({signal_9521, signal_6229}), .c ({signal_9773, signal_6481}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6246 ( .a ({signal_9281, signal_5989}), .b ({signal_9525, signal_6233}), .c ({signal_9774, signal_6482}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6247 ( .a ({signal_9524, signal_6232}), .b ({signal_9526, signal_6234}), .c ({signal_9775, signal_6483}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6248 ( .a ({signal_9522, signal_6230}), .b ({signal_9527, signal_6235}), .c ({signal_9776, signal_6484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6249 ( .a ({signal_9523, signal_6231}), .b ({signal_9527, signal_6235}), .c ({signal_9777, signal_6485}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6250 ( .a ({signal_9525, signal_6233}), .b ({signal_9626, signal_6340}), .c ({signal_9778, signal_6486}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6251 ( .a ({signal_9286, signal_5994}), .b ({signal_9626, signal_6340}), .c ({signal_9779, signal_6487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6252 ( .a ({signal_9526, signal_6234}), .b ({signal_9627, signal_6341}), .c ({signal_9780, signal_6488}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6253 ( .a ({signal_9290, signal_5998}), .b ({signal_9529, signal_6237}), .c ({signal_9781, signal_6489}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6254 ( .a ({signal_9289, signal_5997}), .b ({signal_9533, signal_6241}), .c ({signal_9782, signal_6490}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6255 ( .a ({signal_9532, signal_6240}), .b ({signal_9534, signal_6242}), .c ({signal_9783, signal_6491}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6256 ( .a ({signal_9530, signal_6238}), .b ({signal_9535, signal_6243}), .c ({signal_9784, signal_6492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6257 ( .a ({signal_9531, signal_6239}), .b ({signal_9535, signal_6243}), .c ({signal_9785, signal_6493}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6258 ( .a ({signal_9533, signal_6241}), .b ({signal_9630, signal_6344}), .c ({signal_9786, signal_6494}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6259 ( .a ({signal_9294, signal_6002}), .b ({signal_9630, signal_6344}), .c ({signal_9787, signal_6495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6260 ( .a ({signal_9534, signal_6242}), .b ({signal_9631, signal_6345}), .c ({signal_9788, signal_6496}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6261 ( .a ({signal_9298, signal_6006}), .b ({signal_9537, signal_6245}), .c ({signal_9789, signal_6497}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6262 ( .a ({signal_9297, signal_6005}), .b ({signal_9541, signal_6249}), .c ({signal_9790, signal_6498}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6263 ( .a ({signal_9540, signal_6248}), .b ({signal_9542, signal_6250}), .c ({signal_9791, signal_6499}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6264 ( .a ({signal_9538, signal_6246}), .b ({signal_9543, signal_6251}), .c ({signal_9792, signal_6500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6265 ( .a ({signal_9539, signal_6247}), .b ({signal_9543, signal_6251}), .c ({signal_9793, signal_6501}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6266 ( .a ({signal_9541, signal_6249}), .b ({signal_9634, signal_6348}), .c ({signal_9794, signal_6502}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6267 ( .a ({signal_9302, signal_6010}), .b ({signal_9634, signal_6348}), .c ({signal_9795, signal_6503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6268 ( .a ({signal_9542, signal_6250}), .b ({signal_9635, signal_6349}), .c ({signal_9796, signal_6504}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6269 ( .a ({signal_9306, signal_6014}), .b ({signal_9545, signal_6253}), .c ({signal_9797, signal_6505}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6270 ( .a ({signal_9305, signal_6013}), .b ({signal_9549, signal_6257}), .c ({signal_9798, signal_6506}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6271 ( .a ({signal_9548, signal_6256}), .b ({signal_9550, signal_6258}), .c ({signal_9799, signal_6507}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6272 ( .a ({signal_9546, signal_6254}), .b ({signal_9551, signal_6259}), .c ({signal_9800, signal_6508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6273 ( .a ({signal_9547, signal_6255}), .b ({signal_9551, signal_6259}), .c ({signal_9801, signal_6509}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6274 ( .a ({signal_9549, signal_6257}), .b ({signal_9638, signal_6352}), .c ({signal_9802, signal_6510}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6275 ( .a ({signal_9310, signal_6018}), .b ({signal_9638, signal_6352}), .c ({signal_9803, signal_6511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6276 ( .a ({signal_9550, signal_6258}), .b ({signal_9639, signal_6353}), .c ({signal_9804, signal_6512}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6277 ( .a ({signal_9314, signal_6022}), .b ({signal_9553, signal_6261}), .c ({signal_9805, signal_6513}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6278 ( .a ({signal_9313, signal_6021}), .b ({signal_9557, signal_6265}), .c ({signal_9806, signal_6514}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6279 ( .a ({signal_9556, signal_6264}), .b ({signal_9558, signal_6266}), .c ({signal_9807, signal_6515}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6280 ( .a ({signal_9554, signal_6262}), .b ({signal_9559, signal_6267}), .c ({signal_9808, signal_6516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6281 ( .a ({signal_9555, signal_6263}), .b ({signal_9559, signal_6267}), .c ({signal_9809, signal_6517}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6282 ( .a ({signal_9557, signal_6265}), .b ({signal_9642, signal_6356}), .c ({signal_9810, signal_6518}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6283 ( .a ({signal_9318, signal_6026}), .b ({signal_9642, signal_6356}), .c ({signal_9811, signal_6519}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6284 ( .a ({signal_9558, signal_6266}), .b ({signal_9643, signal_6357}), .c ({signal_9812, signal_6520}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6285 ( .a ({signal_9475, signal_6035}), .b ({signal_9702, signal_6270}), .c ({signal_9897, signal_6521}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6286 ( .a ({signal_9702, signal_6270}), .b ({signal_9710, signal_6362}), .c ({signal_9898, signal_6522}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6287 ( .a ({signal_9469, signal_6029}), .b ({signal_9708, signal_6360}), .c ({signal_9899, signal_6523}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6288 ( .a ({signal_9471, signal_6031}), .b ({signal_9701, signal_6269}), .c ({signal_9900, signal_6524}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6289 ( .a ({signal_9701, signal_6269}), .b ({signal_9709, signal_6361}), .c ({signal_9901, signal_6525}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6290 ( .a ({signal_9236, signal_5844}), .b ({signal_9707, signal_6359}), .c ({signal_9902, signal_6526}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6291 ( .a ({signal_9476, signal_6036}), .b ({signal_9709, signal_6361}), .c ({signal_9903, signal_6527}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6292 ( .a ({signal_9496, signal_6164}), .b ({signal_9708, signal_6360}), .c ({signal_9904, signal_6528}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6293 ( .a ({signal_9707, signal_6359}), .b ({signal_9714, signal_6366}), .c ({signal_9905, signal_6529}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6294 ( .a ({signal_9322, signal_6038}), .b ({signal_9561, signal_6271}), .c ({signal_9813, signal_6530}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6295 ( .a ({signal_9321, signal_6037}), .b ({signal_9565, signal_6275}), .c ({signal_9814, signal_6531}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6296 ( .a ({signal_9564, signal_6274}), .b ({signal_9566, signal_6276}), .c ({signal_9815, signal_6532}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6297 ( .a ({signal_9562, signal_6272}), .b ({signal_9567, signal_6277}), .c ({signal_9816, signal_6533}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6298 ( .a ({signal_9563, signal_6273}), .b ({signal_9567, signal_6277}), .c ({signal_9817, signal_6534}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6299 ( .a ({signal_9565, signal_6275}), .b ({signal_9646, signal_6368}), .c ({signal_9818, signal_6535}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6300 ( .a ({signal_9326, signal_6042}), .b ({signal_9646, signal_6368}), .c ({signal_9819, signal_6536}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6301 ( .a ({signal_9566, signal_6276}), .b ({signal_9647, signal_6369}), .c ({signal_9820, signal_6537}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6302 ( .a ({signal_9330, signal_6046}), .b ({signal_9569, signal_6279}), .c ({signal_9821, signal_6538}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6303 ( .a ({signal_9329, signal_6045}), .b ({signal_9573, signal_6283}), .c ({signal_9822, signal_6539}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6304 ( .a ({signal_9572, signal_6282}), .b ({signal_9574, signal_6284}), .c ({signal_9823, signal_6540}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6305 ( .a ({signal_9570, signal_6280}), .b ({signal_9575, signal_6285}), .c ({signal_9824, signal_6541}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6306 ( .a ({signal_9571, signal_6281}), .b ({signal_9575, signal_6285}), .c ({signal_9825, signal_6542}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6307 ( .a ({signal_9573, signal_6283}), .b ({signal_9650, signal_6372}), .c ({signal_9826, signal_6543}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6308 ( .a ({signal_9334, signal_6050}), .b ({signal_9650, signal_6372}), .c ({signal_9827, signal_6544}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6309 ( .a ({signal_9574, signal_6284}), .b ({signal_9651, signal_6373}), .c ({signal_9828, signal_6545}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6310 ( .a ({signal_9338, signal_6054}), .b ({signal_9577, signal_6287}), .c ({signal_9829, signal_6546}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6311 ( .a ({signal_9337, signal_6053}), .b ({signal_9581, signal_6291}), .c ({signal_9830, signal_6547}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6312 ( .a ({signal_9580, signal_6290}), .b ({signal_9582, signal_6292}), .c ({signal_9831, signal_6548}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6313 ( .a ({signal_9578, signal_6288}), .b ({signal_9583, signal_6293}), .c ({signal_9832, signal_6549}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6314 ( .a ({signal_9579, signal_6289}), .b ({signal_9583, signal_6293}), .c ({signal_9833, signal_6550}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6315 ( .a ({signal_9581, signal_6291}), .b ({signal_9654, signal_6376}), .c ({signal_9834, signal_6551}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6316 ( .a ({signal_9342, signal_6058}), .b ({signal_9654, signal_6376}), .c ({signal_9835, signal_6552}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6317 ( .a ({signal_9582, signal_6292}), .b ({signal_9655, signal_6377}), .c ({signal_9836, signal_6553}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6318 ( .a ({signal_9483, signal_6067}), .b ({signal_9704, signal_6296}), .c ({signal_9906, signal_6554}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6319 ( .a ({signal_9704, signal_6296}), .b ({signal_9718, signal_6382}), .c ({signal_9907, signal_6555}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6320 ( .a ({signal_9477, signal_6061}), .b ({signal_9716, signal_6380}), .c ({signal_9908, signal_6556}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6321 ( .a ({signal_9479, signal_6063}), .b ({signal_9703, signal_6295}), .c ({signal_9909, signal_6557}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6322 ( .a ({signal_9703, signal_6295}), .b ({signal_9717, signal_6381}), .c ({signal_9910, signal_6558}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6323 ( .a ({signal_9244, signal_5852}), .b ({signal_9715, signal_6379}), .c ({signal_9911, signal_6559}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6324 ( .a ({signal_9484, signal_6068}), .b ({signal_9717, signal_6381}), .c ({signal_9912, signal_6560}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6325 ( .a ({signal_9500, signal_6180}), .b ({signal_9716, signal_6380}), .c ({signal_9913, signal_6561}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6326 ( .a ({signal_9715, signal_6379}), .b ({signal_9722, signal_6386}), .c ({signal_9914, signal_6562}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6327 ( .a ({signal_9346, signal_6070}), .b ({signal_9585, signal_6297}), .c ({signal_9837, signal_6563}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6328 ( .a ({signal_9345, signal_6069}), .b ({signal_9589, signal_6301}), .c ({signal_9838, signal_6564}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6329 ( .a ({signal_9588, signal_6300}), .b ({signal_9590, signal_6302}), .c ({signal_9839, signal_6565}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6330 ( .a ({signal_9586, signal_6298}), .b ({signal_9591, signal_6303}), .c ({signal_9840, signal_6566}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6331 ( .a ({signal_9587, signal_6299}), .b ({signal_9591, signal_6303}), .c ({signal_9841, signal_6567}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6332 ( .a ({signal_9589, signal_6301}), .b ({signal_9658, signal_6388}), .c ({signal_9842, signal_6568}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6333 ( .a ({signal_9350, signal_6074}), .b ({signal_9658, signal_6388}), .c ({signal_9843, signal_6569}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6334 ( .a ({signal_9590, signal_6302}), .b ({signal_9659, signal_6389}), .c ({signal_9844, signal_6570}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6335 ( .a ({signal_9354, signal_6078}), .b ({signal_9593, signal_6305}), .c ({signal_9845, signal_6571}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6336 ( .a ({signal_9353, signal_6077}), .b ({signal_9597, signal_6309}), .c ({signal_9846, signal_6572}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6337 ( .a ({signal_9596, signal_6308}), .b ({signal_9598, signal_6310}), .c ({signal_9847, signal_6573}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6338 ( .a ({signal_9594, signal_6306}), .b ({signal_9599, signal_6311}), .c ({signal_9848, signal_6574}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6339 ( .a ({signal_9595, signal_6307}), .b ({signal_9599, signal_6311}), .c ({signal_9849, signal_6575}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6340 ( .a ({signal_9597, signal_6309}), .b ({signal_9662, signal_6392}), .c ({signal_9850, signal_6576}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6341 ( .a ({signal_9358, signal_6082}), .b ({signal_9662, signal_6392}), .c ({signal_9851, signal_6577}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6342 ( .a ({signal_9598, signal_6310}), .b ({signal_9663, signal_6393}), .c ({signal_9852, signal_6578}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6343 ( .a ({signal_9362, signal_6086}), .b ({signal_9601, signal_6313}), .c ({signal_9853, signal_6579}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6344 ( .a ({signal_9361, signal_6085}), .b ({signal_9605, signal_6317}), .c ({signal_9854, signal_6580}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6345 ( .a ({signal_9604, signal_6316}), .b ({signal_9606, signal_6318}), .c ({signal_9855, signal_6581}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6346 ( .a ({signal_9602, signal_6314}), .b ({signal_9607, signal_6319}), .c ({signal_9856, signal_6582}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6347 ( .a ({signal_9603, signal_6315}), .b ({signal_9607, signal_6319}), .c ({signal_9857, signal_6583}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6348 ( .a ({signal_9605, signal_6317}), .b ({signal_9666, signal_6396}), .c ({signal_9858, signal_6584}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6349 ( .a ({signal_9366, signal_6090}), .b ({signal_9666, signal_6396}), .c ({signal_9859, signal_6585}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6350 ( .a ({signal_9606, signal_6318}), .b ({signal_9667, signal_6397}), .c ({signal_9860, signal_6586}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6351 ( .a ({signal_9491, signal_6099}), .b ({signal_9706, signal_6322}), .c ({signal_9915, signal_6587}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6352 ( .a ({signal_9706, signal_6322}), .b ({signal_9726, signal_6402}), .c ({signal_9916, signal_6588}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6353 ( .a ({signal_9485, signal_6093}), .b ({signal_9724, signal_6400}), .c ({signal_9917, signal_6589}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6354 ( .a ({signal_9487, signal_6095}), .b ({signal_9705, signal_6321}), .c ({signal_9918, signal_6590}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6355 ( .a ({signal_9705, signal_6321}), .b ({signal_9725, signal_6401}), .c ({signal_9919, signal_6591}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6356 ( .a ({signal_9252, signal_5860}), .b ({signal_9723, signal_6399}), .c ({signal_9920, signal_6592}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6357 ( .a ({signal_9492, signal_6100}), .b ({signal_9725, signal_6401}), .c ({signal_9921, signal_6593}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6358 ( .a ({signal_9504, signal_6196}), .b ({signal_9724, signal_6400}), .c ({signal_9922, signal_6594}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6359 ( .a ({signal_9723, signal_6399}), .b ({signal_9730, signal_6406}), .c ({signal_9923, signal_6595}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6360 ( .a ({signal_9375, signal_6107}), .b ({signal_9610, signal_6324}), .c ({signal_9861, signal_6596}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6361 ( .a ({signal_9610, signal_6324}), .b ({signal_9672, signal_6410}), .c ({signal_9862, signal_6597}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6362 ( .a ({signal_9369, signal_6101}), .b ({signal_9670, signal_6408}), .c ({signal_9863, signal_6598}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6363 ( .a ({signal_9371, signal_6103}), .b ({signal_9609, signal_6323}), .c ({signal_9864, signal_6599}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6364 ( .a ({signal_9609, signal_6323}), .b ({signal_9671, signal_6409}), .c ({signal_9865, signal_6600}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6365 ( .a ({signal_9136, signal_5868}), .b ({signal_9669, signal_6407}), .c ({signal_9866, signal_6601}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6366 ( .a ({signal_9376, signal_6108}), .b ({signal_9671, signal_6409}), .c ({signal_9867, signal_6602}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6367 ( .a ({signal_9456, signal_6200}), .b ({signal_9670, signal_6408}), .c ({signal_9868, signal_6603}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6368 ( .a ({signal_9669, signal_6407}), .b ({signal_9676, signal_6414}), .c ({signal_9869, signal_6604}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6369 ( .a ({signal_9383, signal_6115}), .b ({signal_9612, signal_6326}), .c ({signal_9870, signal_6605}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6370 ( .a ({signal_9612, signal_6326}), .b ({signal_9680, signal_6418}), .c ({signal_9871, signal_6606}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6371 ( .a ({signal_9377, signal_6109}), .b ({signal_9678, signal_6416}), .c ({signal_9872, signal_6607}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6372 ( .a ({signal_9379, signal_6111}), .b ({signal_9611, signal_6325}), .c ({signal_9873, signal_6608}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6373 ( .a ({signal_9611, signal_6325}), .b ({signal_9679, signal_6417}), .c ({signal_9874, signal_6609}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6374 ( .a ({signal_9144, signal_5876}), .b ({signal_9677, signal_6415}), .c ({signal_9875, signal_6610}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6375 ( .a ({signal_9384, signal_6116}), .b ({signal_9679, signal_6417}), .c ({signal_9876, signal_6611}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6376 ( .a ({signal_9460, signal_6204}), .b ({signal_9678, signal_6416}), .c ({signal_9877, signal_6612}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6377 ( .a ({signal_9677, signal_6415}), .b ({signal_9684, signal_6422}), .c ({signal_9878, signal_6613}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6378 ( .a ({signal_9391, signal_6123}), .b ({signal_9614, signal_6328}), .c ({signal_9879, signal_6614}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6379 ( .a ({signal_9614, signal_6328}), .b ({signal_9688, signal_6426}), .c ({signal_9880, signal_6615}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6380 ( .a ({signal_9385, signal_6117}), .b ({signal_9686, signal_6424}), .c ({signal_9881, signal_6616}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6381 ( .a ({signal_9387, signal_6119}), .b ({signal_9613, signal_6327}), .c ({signal_9882, signal_6617}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6382 ( .a ({signal_9613, signal_6327}), .b ({signal_9687, signal_6425}), .c ({signal_9883, signal_6618}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6383 ( .a ({signal_9152, signal_5884}), .b ({signal_9685, signal_6423}), .c ({signal_9884, signal_6619}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6384 ( .a ({signal_9392, signal_6124}), .b ({signal_9687, signal_6425}), .c ({signal_9885, signal_6620}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6385 ( .a ({signal_9464, signal_6208}), .b ({signal_9686, signal_6424}), .c ({signal_9886, signal_6621}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6386 ( .a ({signal_9685, signal_6423}), .b ({signal_9692, signal_6430}), .c ({signal_9887, signal_6622}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6387 ( .a ({signal_9399, signal_6131}), .b ({signal_9616, signal_6330}), .c ({signal_9888, signal_6623}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6388 ( .a ({signal_9616, signal_6330}), .b ({signal_9696, signal_6434}), .c ({signal_9889, signal_6624}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6389 ( .a ({signal_9393, signal_6125}), .b ({signal_9694, signal_6432}), .c ({signal_9890, signal_6625}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6390 ( .a ({signal_9395, signal_6127}), .b ({signal_9615, signal_6329}), .c ({signal_9891, signal_6626}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6391 ( .a ({signal_9615, signal_6329}), .b ({signal_9695, signal_6433}), .c ({signal_9892, signal_6627}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6392 ( .a ({signal_9160, signal_5892}), .b ({signal_9693, signal_6431}), .c ({signal_9893, signal_6628}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6393 ( .a ({signal_9400, signal_6132}), .b ({signal_9695, signal_6433}), .c ({signal_9894, signal_6629}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6394 ( .a ({signal_9468, signal_6212}), .b ({signal_9694, signal_6432}), .c ({signal_9895, signal_6630}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6395 ( .a ({signal_9693, signal_6431}), .b ({signal_9700, signal_6438}), .c ({signal_9896, signal_6631}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6396 ( .a ({signal_9511, signal_6219}), .b ({signal_9732, signal_6440}), .c ({signal_9924, signal_6632}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6397 ( .a ({signal_9732, signal_6440}), .b ({signal_9760, signal_6468}), .c ({signal_9925, signal_6633}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6398 ( .a ({signal_9505, signal_6213}), .b ({signal_9758, signal_6466}), .c ({signal_9926, signal_6634}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6399 ( .a ({signal_9507, signal_6215}), .b ({signal_9731, signal_6439}), .c ({signal_9927, signal_6635}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6400 ( .a ({signal_9731, signal_6439}), .b ({signal_9759, signal_6467}), .c ({signal_9928, signal_6636}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6401 ( .a ({signal_9272, signal_5980}), .b ({signal_9757, signal_6465}), .c ({signal_9929, signal_6637}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6402 ( .a ({signal_9512, signal_6220}), .b ({signal_9759, signal_6467}), .c ({signal_9930, signal_6638}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6403 ( .a ({signal_9620, signal_6334}), .b ({signal_9758, signal_6466}), .c ({signal_9931, signal_6639}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6404 ( .a ({signal_9757, signal_6465}), .b ({signal_9764, signal_6472}), .c ({signal_9932, signal_6640}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6405 ( .a ({signal_9519, signal_6227}), .b ({signal_9734, signal_6442}), .c ({signal_9933, signal_6641}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6406 ( .a ({signal_9734, signal_6442}), .b ({signal_9768, signal_6476}), .c ({signal_9934, signal_6642}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6407 ( .a ({signal_9513, signal_6221}), .b ({signal_9766, signal_6474}), .c ({signal_9935, signal_6643}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6408 ( .a ({signal_9515, signal_6223}), .b ({signal_9733, signal_6441}), .c ({signal_9936, signal_6644}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6409 ( .a ({signal_9733, signal_6441}), .b ({signal_9767, signal_6475}), .c ({signal_9937, signal_6645}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6410 ( .a ({signal_9280, signal_5988}), .b ({signal_9765, signal_6473}), .c ({signal_9938, signal_6646}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6411 ( .a ({signal_9520, signal_6228}), .b ({signal_9767, signal_6475}), .c ({signal_9939, signal_6647}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6412 ( .a ({signal_9624, signal_6338}), .b ({signal_9766, signal_6474}), .c ({signal_9940, signal_6648}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6413 ( .a ({signal_9765, signal_6473}), .b ({signal_9772, signal_6480}), .c ({signal_9941, signal_6649}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6414 ( .a ({signal_9527, signal_6235}), .b ({signal_9736, signal_6444}), .c ({signal_9942, signal_6650}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6415 ( .a ({signal_9736, signal_6444}), .b ({signal_9776, signal_6484}), .c ({signal_9943, signal_6651}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6416 ( .a ({signal_9521, signal_6229}), .b ({signal_9774, signal_6482}), .c ({signal_9944, signal_6652}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6417 ( .a ({signal_9523, signal_6231}), .b ({signal_9735, signal_6443}), .c ({signal_9945, signal_6653}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6418 ( .a ({signal_9735, signal_6443}), .b ({signal_9775, signal_6483}), .c ({signal_9946, signal_6654}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6419 ( .a ({signal_9288, signal_5996}), .b ({signal_9773, signal_6481}), .c ({signal_9947, signal_6655}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6420 ( .a ({signal_9528, signal_6236}), .b ({signal_9775, signal_6483}), .c ({signal_9948, signal_6656}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6421 ( .a ({signal_9628, signal_6342}), .b ({signal_9774, signal_6482}), .c ({signal_9949, signal_6657}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6422 ( .a ({signal_9773, signal_6481}), .b ({signal_9780, signal_6488}), .c ({signal_9950, signal_6658}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6423 ( .a ({signal_9535, signal_6243}), .b ({signal_9738, signal_6446}), .c ({signal_9951, signal_6659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6424 ( .a ({signal_9738, signal_6446}), .b ({signal_9784, signal_6492}), .c ({signal_9952, signal_6660}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6425 ( .a ({signal_9529, signal_6237}), .b ({signal_9782, signal_6490}), .c ({signal_9953, signal_6661}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6426 ( .a ({signal_9531, signal_6239}), .b ({signal_9737, signal_6445}), .c ({signal_9954, signal_6662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6427 ( .a ({signal_9737, signal_6445}), .b ({signal_9783, signal_6491}), .c ({signal_9955, signal_6663}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6428 ( .a ({signal_9296, signal_6004}), .b ({signal_9781, signal_6489}), .c ({signal_9956, signal_6664}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6429 ( .a ({signal_9536, signal_6244}), .b ({signal_9783, signal_6491}), .c ({signal_9957, signal_6665}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6430 ( .a ({signal_9632, signal_6346}), .b ({signal_9782, signal_6490}), .c ({signal_9958, signal_6666}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6431 ( .a ({signal_9781, signal_6489}), .b ({signal_9788, signal_6496}), .c ({signal_9959, signal_6667}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6432 ( .a ({signal_9543, signal_6251}), .b ({signal_9740, signal_6448}), .c ({signal_9960, signal_6668}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6433 ( .a ({signal_9740, signal_6448}), .b ({signal_9792, signal_6500}), .c ({signal_9961, signal_6669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6434 ( .a ({signal_9537, signal_6245}), .b ({signal_9790, signal_6498}), .c ({signal_9962, signal_6670}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6435 ( .a ({signal_9539, signal_6247}), .b ({signal_9739, signal_6447}), .c ({signal_9963, signal_6671}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6436 ( .a ({signal_9739, signal_6447}), .b ({signal_9791, signal_6499}), .c ({signal_9964, signal_6672}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6437 ( .a ({signal_9304, signal_6012}), .b ({signal_9789, signal_6497}), .c ({signal_9965, signal_6673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6438 ( .a ({signal_9544, signal_6252}), .b ({signal_9791, signal_6499}), .c ({signal_9966, signal_6674}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6439 ( .a ({signal_9636, signal_6350}), .b ({signal_9790, signal_6498}), .c ({signal_9967, signal_6675}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6440 ( .a ({signal_9789, signal_6497}), .b ({signal_9796, signal_6504}), .c ({signal_9968, signal_6676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6441 ( .a ({signal_9551, signal_6259}), .b ({signal_9742, signal_6450}), .c ({signal_9969, signal_6677}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6442 ( .a ({signal_9742, signal_6450}), .b ({signal_9800, signal_6508}), .c ({signal_9970, signal_6678}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6443 ( .a ({signal_9545, signal_6253}), .b ({signal_9798, signal_6506}), .c ({signal_9971, signal_6679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6444 ( .a ({signal_9547, signal_6255}), .b ({signal_9741, signal_6449}), .c ({signal_9972, signal_6680}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6445 ( .a ({signal_9741, signal_6449}), .b ({signal_9799, signal_6507}), .c ({signal_9973, signal_6681}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6446 ( .a ({signal_9312, signal_6020}), .b ({signal_9797, signal_6505}), .c ({signal_9974, signal_6682}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6447 ( .a ({signal_9552, signal_6260}), .b ({signal_9799, signal_6507}), .c ({signal_9975, signal_6683}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6448 ( .a ({signal_9640, signal_6354}), .b ({signal_9798, signal_6506}), .c ({signal_9976, signal_6684}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6449 ( .a ({signal_9797, signal_6505}), .b ({signal_9804, signal_6512}), .c ({signal_9977, signal_6685}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6450 ( .a ({signal_9559, signal_6267}), .b ({signal_9744, signal_6452}), .c ({signal_9978, signal_6686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6451 ( .a ({signal_9744, signal_6452}), .b ({signal_9808, signal_6516}), .c ({signal_9979, signal_6687}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6452 ( .a ({signal_9553, signal_6261}), .b ({signal_9806, signal_6514}), .c ({signal_9980, signal_6688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6453 ( .a ({signal_9555, signal_6263}), .b ({signal_9743, signal_6451}), .c ({signal_9981, signal_6689}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6454 ( .a ({signal_9743, signal_6451}), .b ({signal_9807, signal_6515}), .c ({signal_9982, signal_6690}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6455 ( .a ({signal_9320, signal_6028}), .b ({signal_9805, signal_6513}), .c ({signal_9983, signal_6691}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6456 ( .a ({signal_9560, signal_6268}), .b ({signal_9807, signal_6515}), .c ({signal_9984, signal_6692}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6457 ( .a ({signal_9644, signal_6358}), .b ({signal_9806, signal_6514}), .c ({signal_9985, signal_6693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6458 ( .a ({signal_9805, signal_6513}), .b ({signal_9812, signal_6520}), .c ({signal_9986, signal_6694}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6459 ( .a ({signal_9231, signal_5839}), .b ({signal_9897, signal_6521}), .c ({signal_10085, signal_6695}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6460 ( .a ({signal_9233, signal_5841}), .b ({signal_9897, signal_6521}), .c ({signal_10086, signal_6696}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6461 ( .a ({signal_9494, signal_6162}), .b ({signal_9897, signal_6521}), .c ({signal_10087, signal_6697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6462 ( .a ({signal_9494, signal_6162}), .b ({signal_9899, signal_6523}), .c ({signal_10088, signal_6698}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6463 ( .a ({signal_9712, signal_6364}), .b ({signal_9900, signal_6524}), .c ({signal_10089, signal_6699}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6464 ( .a ({signal_9898, signal_6522}), .b ({signal_9901, signal_6525}), .c ({signal_10090, signal_6700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6465 ( .a ({signal_9899, signal_6523}), .b ({signal_9900, signal_6524}), .c ({signal_10091, signal_6701}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6466 ( .a ({signal_9495, signal_6163}), .b ({signal_9901, signal_6525}), .c ({signal_10092, signal_6702}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6467 ( .a ({signal_9711, signal_6363}), .b ({signal_9902, signal_6526}), .c ({signal_10093, signal_6703}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6468 ( .a ({signal_9713, signal_6365}), .b ({signal_9902, signal_6526}), .c ({signal_10094, signal_6704}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6469 ( .a ({signal_9898, signal_6522}), .b ({signal_9905, signal_6529}), .c ({signal_10095, signal_6705}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6470 ( .a ({signal_9567, signal_6277}), .b ({signal_9746, signal_6454}), .c ({signal_9987, signal_6706}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6471 ( .a ({signal_9746, signal_6454}), .b ({signal_9816, signal_6533}), .c ({signal_9988, signal_6707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6472 ( .a ({signal_9561, signal_6271}), .b ({signal_9814, signal_6531}), .c ({signal_9989, signal_6708}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6473 ( .a ({signal_9563, signal_6273}), .b ({signal_9745, signal_6453}), .c ({signal_9990, signal_6709}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6474 ( .a ({signal_9745, signal_6453}), .b ({signal_9815, signal_6532}), .c ({signal_9991, signal_6710}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6475 ( .a ({signal_9328, signal_6044}), .b ({signal_9813, signal_6530}), .c ({signal_9992, signal_6711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6476 ( .a ({signal_9568, signal_6278}), .b ({signal_9815, signal_6532}), .c ({signal_9993, signal_6712}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6477 ( .a ({signal_9648, signal_6370}), .b ({signal_9814, signal_6531}), .c ({signal_9994, signal_6713}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6478 ( .a ({signal_9813, signal_6530}), .b ({signal_9820, signal_6537}), .c ({signal_9995, signal_6714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6479 ( .a ({signal_9575, signal_6285}), .b ({signal_9748, signal_6456}), .c ({signal_9996, signal_6715}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6480 ( .a ({signal_9748, signal_6456}), .b ({signal_9824, signal_6541}), .c ({signal_9997, signal_6716}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6481 ( .a ({signal_9569, signal_6279}), .b ({signal_9822, signal_6539}), .c ({signal_9998, signal_6717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6482 ( .a ({signal_9571, signal_6281}), .b ({signal_9747, signal_6455}), .c ({signal_9999, signal_6718}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6483 ( .a ({signal_9747, signal_6455}), .b ({signal_9823, signal_6540}), .c ({signal_10000, signal_6719}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6484 ( .a ({signal_9336, signal_6052}), .b ({signal_9821, signal_6538}), .c ({signal_10001, signal_6720}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6485 ( .a ({signal_9576, signal_6286}), .b ({signal_9823, signal_6540}), .c ({signal_10002, signal_6721}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6486 ( .a ({signal_9652, signal_6374}), .b ({signal_9822, signal_6539}), .c ({signal_10003, signal_6722}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6487 ( .a ({signal_9821, signal_6538}), .b ({signal_9828, signal_6545}), .c ({signal_10004, signal_6723}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6488 ( .a ({signal_9583, signal_6293}), .b ({signal_9750, signal_6458}), .c ({signal_10005, signal_6724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6489 ( .a ({signal_9750, signal_6458}), .b ({signal_9832, signal_6549}), .c ({signal_10006, signal_6725}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6490 ( .a ({signal_9577, signal_6287}), .b ({signal_9830, signal_6547}), .c ({signal_10007, signal_6726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6491 ( .a ({signal_9579, signal_6289}), .b ({signal_9749, signal_6457}), .c ({signal_10008, signal_6727}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6492 ( .a ({signal_9749, signal_6457}), .b ({signal_9831, signal_6548}), .c ({signal_10009, signal_6728}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6493 ( .a ({signal_9344, signal_6060}), .b ({signal_9829, signal_6546}), .c ({signal_10010, signal_6729}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6494 ( .a ({signal_9584, signal_6294}), .b ({signal_9831, signal_6548}), .c ({signal_10011, signal_6730}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6495 ( .a ({signal_9656, signal_6378}), .b ({signal_9830, signal_6547}), .c ({signal_10012, signal_6731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6496 ( .a ({signal_9829, signal_6546}), .b ({signal_9836, signal_6553}), .c ({signal_10013, signal_6732}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6497 ( .a ({signal_9239, signal_5847}), .b ({signal_9906, signal_6554}), .c ({signal_10096, signal_6733}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6498 ( .a ({signal_9241, signal_5849}), .b ({signal_9906, signal_6554}), .c ({signal_10097, signal_6734}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6499 ( .a ({signal_9498, signal_6178}), .b ({signal_9906, signal_6554}), .c ({signal_10098, signal_6735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6500 ( .a ({signal_9498, signal_6178}), .b ({signal_9908, signal_6556}), .c ({signal_10099, signal_6736}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6501 ( .a ({signal_9720, signal_6384}), .b ({signal_9909, signal_6557}), .c ({signal_10100, signal_6737}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6502 ( .a ({signal_9907, signal_6555}), .b ({signal_9910, signal_6558}), .c ({signal_10101, signal_6738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6503 ( .a ({signal_9908, signal_6556}), .b ({signal_9909, signal_6557}), .c ({signal_10102, signal_6739}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6504 ( .a ({signal_9499, signal_6179}), .b ({signal_9910, signal_6558}), .c ({signal_10103, signal_6740}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6505 ( .a ({signal_9719, signal_6383}), .b ({signal_9911, signal_6559}), .c ({signal_10104, signal_6741}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6506 ( .a ({signal_9721, signal_6385}), .b ({signal_9911, signal_6559}), .c ({signal_10105, signal_6742}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6507 ( .a ({signal_9907, signal_6555}), .b ({signal_9914, signal_6562}), .c ({signal_10106, signal_6743}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6508 ( .a ({signal_9591, signal_6303}), .b ({signal_9752, signal_6460}), .c ({signal_10014, signal_6744}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6509 ( .a ({signal_9752, signal_6460}), .b ({signal_9840, signal_6566}), .c ({signal_10015, signal_6745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6510 ( .a ({signal_9585, signal_6297}), .b ({signal_9838, signal_6564}), .c ({signal_10016, signal_6746}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6511 ( .a ({signal_9587, signal_6299}), .b ({signal_9751, signal_6459}), .c ({signal_10017, signal_6747}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6512 ( .a ({signal_9751, signal_6459}), .b ({signal_9839, signal_6565}), .c ({signal_10018, signal_6748}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6513 ( .a ({signal_9352, signal_6076}), .b ({signal_9837, signal_6563}), .c ({signal_10019, signal_6749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6514 ( .a ({signal_9592, signal_6304}), .b ({signal_9839, signal_6565}), .c ({signal_10020, signal_6750}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6515 ( .a ({signal_9660, signal_6390}), .b ({signal_9838, signal_6564}), .c ({signal_10021, signal_6751}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6516 ( .a ({signal_9837, signal_6563}), .b ({signal_9844, signal_6570}), .c ({signal_10022, signal_6752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6517 ( .a ({signal_9599, signal_6311}), .b ({signal_9754, signal_6462}), .c ({signal_10023, signal_6753}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6518 ( .a ({signal_9754, signal_6462}), .b ({signal_9848, signal_6574}), .c ({signal_10024, signal_6754}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6519 ( .a ({signal_9593, signal_6305}), .b ({signal_9846, signal_6572}), .c ({signal_10025, signal_6755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6520 ( .a ({signal_9595, signal_6307}), .b ({signal_9753, signal_6461}), .c ({signal_10026, signal_6756}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6521 ( .a ({signal_9753, signal_6461}), .b ({signal_9847, signal_6573}), .c ({signal_10027, signal_6757}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6522 ( .a ({signal_9360, signal_6084}), .b ({signal_9845, signal_6571}), .c ({signal_10028, signal_6758}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6523 ( .a ({signal_9600, signal_6312}), .b ({signal_9847, signal_6573}), .c ({signal_10029, signal_6759}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6524 ( .a ({signal_9664, signal_6394}), .b ({signal_9846, signal_6572}), .c ({signal_10030, signal_6760}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6525 ( .a ({signal_9845, signal_6571}), .b ({signal_9852, signal_6578}), .c ({signal_10031, signal_6761}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6526 ( .a ({signal_9607, signal_6319}), .b ({signal_9756, signal_6464}), .c ({signal_10032, signal_6762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6527 ( .a ({signal_9756, signal_6464}), .b ({signal_9856, signal_6582}), .c ({signal_10033, signal_6763}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6528 ( .a ({signal_9601, signal_6313}), .b ({signal_9854, signal_6580}), .c ({signal_10034, signal_6764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6529 ( .a ({signal_9603, signal_6315}), .b ({signal_9755, signal_6463}), .c ({signal_10035, signal_6765}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6530 ( .a ({signal_9755, signal_6463}), .b ({signal_9855, signal_6581}), .c ({signal_10036, signal_6766}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6531 ( .a ({signal_9368, signal_6092}), .b ({signal_9853, signal_6579}), .c ({signal_10037, signal_6767}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6532 ( .a ({signal_9608, signal_6320}), .b ({signal_9855, signal_6581}), .c ({signal_10038, signal_6768}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6533 ( .a ({signal_9668, signal_6398}), .b ({signal_9854, signal_6580}), .c ({signal_10039, signal_6769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6534 ( .a ({signal_9853, signal_6579}), .b ({signal_9860, signal_6586}), .c ({signal_10040, signal_6770}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6535 ( .a ({signal_9247, signal_5855}), .b ({signal_9915, signal_6587}), .c ({signal_10107, signal_6771}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6536 ( .a ({signal_9249, signal_5857}), .b ({signal_9915, signal_6587}), .c ({signal_10108, signal_6772}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6537 ( .a ({signal_9502, signal_6194}), .b ({signal_9915, signal_6587}), .c ({signal_10109, signal_6773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6538 ( .a ({signal_9502, signal_6194}), .b ({signal_9917, signal_6589}), .c ({signal_10110, signal_6774}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6539 ( .a ({signal_9728, signal_6404}), .b ({signal_9918, signal_6590}), .c ({signal_10111, signal_6775}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6540 ( .a ({signal_9916, signal_6588}), .b ({signal_9919, signal_6591}), .c ({signal_10112, signal_6776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6541 ( .a ({signal_9917, signal_6589}), .b ({signal_9918, signal_6590}), .c ({signal_10113, signal_6777}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6542 ( .a ({signal_9503, signal_6195}), .b ({signal_9919, signal_6591}), .c ({signal_10114, signal_6778}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6543 ( .a ({signal_9727, signal_6403}), .b ({signal_9920, signal_6592}), .c ({signal_10115, signal_6779}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6544 ( .a ({signal_9729, signal_6405}), .b ({signal_9920, signal_6592}), .c ({signal_10116, signal_6780}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6545 ( .a ({signal_9916, signal_6588}), .b ({signal_9923, signal_6595}), .c ({signal_10117, signal_6781}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6546 ( .a ({signal_9131, signal_5863}), .b ({signal_9861, signal_6596}), .c ({signal_10041, signal_6782}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6547 ( .a ({signal_9133, signal_5865}), .b ({signal_9861, signal_6596}), .c ({signal_10042, signal_6783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6548 ( .a ({signal_9454, signal_6198}), .b ({signal_9861, signal_6596}), .c ({signal_10043, signal_6784}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6549 ( .a ({signal_9454, signal_6198}), .b ({signal_9863, signal_6598}), .c ({signal_10044, signal_6785}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6550 ( .a ({signal_9674, signal_6412}), .b ({signal_9864, signal_6599}), .c ({signal_10045, signal_6786}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6551 ( .a ({signal_9862, signal_6597}), .b ({signal_9865, signal_6600}), .c ({signal_10046, signal_6787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6552 ( .a ({signal_9863, signal_6598}), .b ({signal_9864, signal_6599}), .c ({signal_10047, signal_6788}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6553 ( .a ({signal_9455, signal_6199}), .b ({signal_9865, signal_6600}), .c ({signal_10048, signal_6789}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6554 ( .a ({signal_9673, signal_6411}), .b ({signal_9866, signal_6601}), .c ({signal_10049, signal_6790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6555 ( .a ({signal_9675, signal_6413}), .b ({signal_9866, signal_6601}), .c ({signal_10050, signal_6791}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6556 ( .a ({signal_9862, signal_6597}), .b ({signal_9869, signal_6604}), .c ({signal_10051, signal_6792}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6557 ( .a ({signal_9139, signal_5871}), .b ({signal_9870, signal_6605}), .c ({signal_10052, signal_6793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6558 ( .a ({signal_9141, signal_5873}), .b ({signal_9870, signal_6605}), .c ({signal_10053, signal_6794}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6559 ( .a ({signal_9458, signal_6202}), .b ({signal_9870, signal_6605}), .c ({signal_10054, signal_6795}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6560 ( .a ({signal_9458, signal_6202}), .b ({signal_9872, signal_6607}), .c ({signal_10055, signal_6796}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6561 ( .a ({signal_9682, signal_6420}), .b ({signal_9873, signal_6608}), .c ({signal_10056, signal_6797}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6562 ( .a ({signal_9871, signal_6606}), .b ({signal_9874, signal_6609}), .c ({signal_10057, signal_6798}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6563 ( .a ({signal_9872, signal_6607}), .b ({signal_9873, signal_6608}), .c ({signal_10058, signal_6799}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6564 ( .a ({signal_9459, signal_6203}), .b ({signal_9874, signal_6609}), .c ({signal_10059, signal_6800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6565 ( .a ({signal_9681, signal_6419}), .b ({signal_9875, signal_6610}), .c ({signal_10060, signal_6801}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6566 ( .a ({signal_9683, signal_6421}), .b ({signal_9875, signal_6610}), .c ({signal_10061, signal_6802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6567 ( .a ({signal_9871, signal_6606}), .b ({signal_9878, signal_6613}), .c ({signal_10062, signal_6803}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6568 ( .a ({signal_9147, signal_5879}), .b ({signal_9879, signal_6614}), .c ({signal_10063, signal_6804}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6569 ( .a ({signal_9149, signal_5881}), .b ({signal_9879, signal_6614}), .c ({signal_10064, signal_6805}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6570 ( .a ({signal_9462, signal_6206}), .b ({signal_9879, signal_6614}), .c ({signal_10065, signal_6806}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6571 ( .a ({signal_9462, signal_6206}), .b ({signal_9881, signal_6616}), .c ({signal_10066, signal_6807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6572 ( .a ({signal_9690, signal_6428}), .b ({signal_9882, signal_6617}), .c ({signal_10067, signal_6808}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6573 ( .a ({signal_9880, signal_6615}), .b ({signal_9883, signal_6618}), .c ({signal_10068, signal_6809}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6574 ( .a ({signal_9881, signal_6616}), .b ({signal_9882, signal_6617}), .c ({signal_10069, signal_6810}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6575 ( .a ({signal_9463, signal_6207}), .b ({signal_9883, signal_6618}), .c ({signal_10070, signal_6811}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6576 ( .a ({signal_9689, signal_6427}), .b ({signal_9884, signal_6619}), .c ({signal_10071, signal_6812}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6577 ( .a ({signal_9691, signal_6429}), .b ({signal_9884, signal_6619}), .c ({signal_10072, signal_6813}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6578 ( .a ({signal_9880, signal_6615}), .b ({signal_9887, signal_6622}), .c ({signal_10073, signal_6814}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6579 ( .a ({signal_9155, signal_5887}), .b ({signal_9888, signal_6623}), .c ({signal_10074, signal_6815}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6580 ( .a ({signal_9157, signal_5889}), .b ({signal_9888, signal_6623}), .c ({signal_10075, signal_6816}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6581 ( .a ({signal_9466, signal_6210}), .b ({signal_9888, signal_6623}), .c ({signal_10076, signal_6817}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6582 ( .a ({signal_9466, signal_6210}), .b ({signal_9890, signal_6625}), .c ({signal_10077, signal_6818}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6583 ( .a ({signal_9698, signal_6436}), .b ({signal_9891, signal_6626}), .c ({signal_10078, signal_6819}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6584 ( .a ({signal_9889, signal_6624}), .b ({signal_9892, signal_6627}), .c ({signal_10079, signal_6820}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6585 ( .a ({signal_9890, signal_6625}), .b ({signal_9891, signal_6626}), .c ({signal_10080, signal_6821}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6586 ( .a ({signal_9467, signal_6211}), .b ({signal_9892, signal_6627}), .c ({signal_10081, signal_6822}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6587 ( .a ({signal_9697, signal_6435}), .b ({signal_9893, signal_6628}), .c ({signal_10082, signal_6823}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6588 ( .a ({signal_9699, signal_6437}), .b ({signal_9893, signal_6628}), .c ({signal_10083, signal_6824}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6589 ( .a ({signal_9889, signal_6624}), .b ({signal_9896, signal_6631}), .c ({signal_10084, signal_6825}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6590 ( .a ({signal_10095, signal_6705}), .b ({signal_10298, signal_3938}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6591 ( .a ({signal_10106, signal_6743}), .b ({signal_10299, signal_3906}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6592 ( .a ({signal_10117, signal_6781}), .b ({signal_10300, signal_3874}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6593 ( .a ({signal_10051, signal_6792}), .b ({signal_10118, signal_3109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6594 ( .a ({signal_9267, signal_5975}), .b ({signal_9924, signal_6632}), .c ({signal_10119, signal_6826}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6595 ( .a ({signal_9269, signal_5977}), .b ({signal_9924, signal_6632}), .c ({signal_10120, signal_6827}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6596 ( .a ({signal_9618, signal_6332}), .b ({signal_9924, signal_6632}), .c ({signal_10121, signal_6828}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6597 ( .a ({signal_9618, signal_6332}), .b ({signal_9926, signal_6634}), .c ({signal_10122, signal_6829}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6598 ( .a ({signal_9762, signal_6470}), .b ({signal_9927, signal_6635}), .c ({signal_10123, signal_6830}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6599 ( .a ({signal_9925, signal_6633}), .b ({signal_9928, signal_6636}), .c ({signal_10124, signal_6831}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6600 ( .a ({signal_9926, signal_6634}), .b ({signal_9927, signal_6635}), .c ({signal_10125, signal_6832}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6601 ( .a ({signal_9619, signal_6333}), .b ({signal_9928, signal_6636}), .c ({signal_10126, signal_6833}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6602 ( .a ({signal_9761, signal_6469}), .b ({signal_9929, signal_6637}), .c ({signal_10127, signal_6834}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6603 ( .a ({signal_9763, signal_6471}), .b ({signal_9929, signal_6637}), .c ({signal_10128, signal_6835}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6604 ( .a ({signal_9925, signal_6633}), .b ({signal_9932, signal_6640}), .c ({signal_10129, signal_6836}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6605 ( .a ({signal_9275, signal_5983}), .b ({signal_9933, signal_6641}), .c ({signal_10130, signal_6837}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6606 ( .a ({signal_9277, signal_5985}), .b ({signal_9933, signal_6641}), .c ({signal_10131, signal_6838}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6607 ( .a ({signal_9622, signal_6336}), .b ({signal_9933, signal_6641}), .c ({signal_10132, signal_6839}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6608 ( .a ({signal_9622, signal_6336}), .b ({signal_9935, signal_6643}), .c ({signal_10133, signal_6840}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6609 ( .a ({signal_9770, signal_6478}), .b ({signal_9936, signal_6644}), .c ({signal_10134, signal_6841}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6610 ( .a ({signal_9934, signal_6642}), .b ({signal_9937, signal_6645}), .c ({signal_10135, signal_6842}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6611 ( .a ({signal_9935, signal_6643}), .b ({signal_9936, signal_6644}), .c ({signal_10136, signal_6843}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6612 ( .a ({signal_9623, signal_6337}), .b ({signal_9937, signal_6645}), .c ({signal_10137, signal_6844}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6613 ( .a ({signal_9769, signal_6477}), .b ({signal_9938, signal_6646}), .c ({signal_10138, signal_6845}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6614 ( .a ({signal_9771, signal_6479}), .b ({signal_9938, signal_6646}), .c ({signal_10139, signal_6846}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6615 ( .a ({signal_9934, signal_6642}), .b ({signal_9941, signal_6649}), .c ({signal_10140, signal_6847}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6616 ( .a ({signal_9283, signal_5991}), .b ({signal_9942, signal_6650}), .c ({signal_10141, signal_6848}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6617 ( .a ({signal_9285, signal_5993}), .b ({signal_9942, signal_6650}), .c ({signal_10142, signal_6849}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6618 ( .a ({signal_9626, signal_6340}), .b ({signal_9942, signal_6650}), .c ({signal_10143, signal_6850}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6619 ( .a ({signal_9626, signal_6340}), .b ({signal_9944, signal_6652}), .c ({signal_10144, signal_6851}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6620 ( .a ({signal_9778, signal_6486}), .b ({signal_9945, signal_6653}), .c ({signal_10145, signal_6852}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6621 ( .a ({signal_9943, signal_6651}), .b ({signal_9946, signal_6654}), .c ({signal_10146, signal_6853}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6622 ( .a ({signal_9944, signal_6652}), .b ({signal_9945, signal_6653}), .c ({signal_10147, signal_6854}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6623 ( .a ({signal_9627, signal_6341}), .b ({signal_9946, signal_6654}), .c ({signal_10148, signal_6855}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6624 ( .a ({signal_9777, signal_6485}), .b ({signal_9947, signal_6655}), .c ({signal_10149, signal_6856}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6625 ( .a ({signal_9779, signal_6487}), .b ({signal_9947, signal_6655}), .c ({signal_10150, signal_6857}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6626 ( .a ({signal_9943, signal_6651}), .b ({signal_9950, signal_6658}), .c ({signal_10151, signal_6858}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6627 ( .a ({signal_9291, signal_5999}), .b ({signal_9951, signal_6659}), .c ({signal_10152, signal_6859}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6628 ( .a ({signal_9293, signal_6001}), .b ({signal_9951, signal_6659}), .c ({signal_10153, signal_6860}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6629 ( .a ({signal_9630, signal_6344}), .b ({signal_9951, signal_6659}), .c ({signal_10154, signal_6861}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6630 ( .a ({signal_9630, signal_6344}), .b ({signal_9953, signal_6661}), .c ({signal_10155, signal_6862}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6631 ( .a ({signal_9786, signal_6494}), .b ({signal_9954, signal_6662}), .c ({signal_10156, signal_6863}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6632 ( .a ({signal_9952, signal_6660}), .b ({signal_9955, signal_6663}), .c ({signal_10157, signal_6864}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6633 ( .a ({signal_9953, signal_6661}), .b ({signal_9954, signal_6662}), .c ({signal_10158, signal_6865}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6634 ( .a ({signal_9631, signal_6345}), .b ({signal_9955, signal_6663}), .c ({signal_10159, signal_6866}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6635 ( .a ({signal_9785, signal_6493}), .b ({signal_9956, signal_6664}), .c ({signal_10160, signal_6867}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6636 ( .a ({signal_9787, signal_6495}), .b ({signal_9956, signal_6664}), .c ({signal_10161, signal_6868}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6637 ( .a ({signal_9952, signal_6660}), .b ({signal_9959, signal_6667}), .c ({signal_10162, signal_6869}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6638 ( .a ({signal_9299, signal_6007}), .b ({signal_9960, signal_6668}), .c ({signal_10163, signal_6870}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6639 ( .a ({signal_9301, signal_6009}), .b ({signal_9960, signal_6668}), .c ({signal_10164, signal_6871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6640 ( .a ({signal_9634, signal_6348}), .b ({signal_9960, signal_6668}), .c ({signal_10165, signal_6872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6641 ( .a ({signal_9634, signal_6348}), .b ({signal_9962, signal_6670}), .c ({signal_10166, signal_6873}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6642 ( .a ({signal_9794, signal_6502}), .b ({signal_9963, signal_6671}), .c ({signal_10167, signal_6874}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6643 ( .a ({signal_9961, signal_6669}), .b ({signal_9964, signal_6672}), .c ({signal_10168, signal_6875}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6644 ( .a ({signal_9962, signal_6670}), .b ({signal_9963, signal_6671}), .c ({signal_10169, signal_6876}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6645 ( .a ({signal_9635, signal_6349}), .b ({signal_9964, signal_6672}), .c ({signal_10170, signal_6877}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6646 ( .a ({signal_9793, signal_6501}), .b ({signal_9965, signal_6673}), .c ({signal_10171, signal_6878}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6647 ( .a ({signal_9795, signal_6503}), .b ({signal_9965, signal_6673}), .c ({signal_10172, signal_6879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6648 ( .a ({signal_9961, signal_6669}), .b ({signal_9968, signal_6676}), .c ({signal_10173, signal_6880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6649 ( .a ({signal_9307, signal_6015}), .b ({signal_9969, signal_6677}), .c ({signal_10174, signal_6881}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6650 ( .a ({signal_9309, signal_6017}), .b ({signal_9969, signal_6677}), .c ({signal_10175, signal_6882}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6651 ( .a ({signal_9638, signal_6352}), .b ({signal_9969, signal_6677}), .c ({signal_10176, signal_6883}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6652 ( .a ({signal_9638, signal_6352}), .b ({signal_9971, signal_6679}), .c ({signal_10177, signal_6884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6653 ( .a ({signal_9802, signal_6510}), .b ({signal_9972, signal_6680}), .c ({signal_10178, signal_6885}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6654 ( .a ({signal_9970, signal_6678}), .b ({signal_9973, signal_6681}), .c ({signal_10179, signal_6886}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6655 ( .a ({signal_9971, signal_6679}), .b ({signal_9972, signal_6680}), .c ({signal_10180, signal_6887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6656 ( .a ({signal_9639, signal_6353}), .b ({signal_9973, signal_6681}), .c ({signal_10181, signal_6888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6657 ( .a ({signal_9801, signal_6509}), .b ({signal_9974, signal_6682}), .c ({signal_10182, signal_6889}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6658 ( .a ({signal_9803, signal_6511}), .b ({signal_9974, signal_6682}), .c ({signal_10183, signal_6890}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6659 ( .a ({signal_9970, signal_6678}), .b ({signal_9977, signal_6685}), .c ({signal_10184, signal_6891}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6660 ( .a ({signal_9315, signal_6023}), .b ({signal_9978, signal_6686}), .c ({signal_10185, signal_6892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6661 ( .a ({signal_9317, signal_6025}), .b ({signal_9978, signal_6686}), .c ({signal_10186, signal_6893}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6662 ( .a ({signal_9642, signal_6356}), .b ({signal_9978, signal_6686}), .c ({signal_10187, signal_6894}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6663 ( .a ({signal_9642, signal_6356}), .b ({signal_9980, signal_6688}), .c ({signal_10188, signal_6895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6664 ( .a ({signal_9810, signal_6518}), .b ({signal_9981, signal_6689}), .c ({signal_10189, signal_6896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6665 ( .a ({signal_9979, signal_6687}), .b ({signal_9982, signal_6690}), .c ({signal_10190, signal_6897}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6666 ( .a ({signal_9980, signal_6688}), .b ({signal_9981, signal_6689}), .c ({signal_10191, signal_6898}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6667 ( .a ({signal_9643, signal_6357}), .b ({signal_9982, signal_6690}), .c ({signal_10192, signal_6899}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6668 ( .a ({signal_9809, signal_6517}), .b ({signal_9983, signal_6691}), .c ({signal_10193, signal_6900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6669 ( .a ({signal_9811, signal_6519}), .b ({signal_9983, signal_6691}), .c ({signal_10194, signal_6901}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6670 ( .a ({signal_9979, signal_6687}), .b ({signal_9986, signal_6694}), .c ({signal_10195, signal_6902}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6671 ( .a ({signal_9898, signal_6522}), .b ({signal_10089, signal_6699}), .c ({signal_10301, signal_4460}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6672 ( .a ({signal_10086, signal_6696}), .b ({signal_10091, signal_6701}), .c ({signal_10302, signal_6903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6673 ( .a ({signal_9903, signal_6527}), .b ({signal_10093, signal_6703}), .c ({signal_10303, signal_6904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6674 ( .a ({signal_9898, signal_6522}), .b ({signal_10088, signal_6698}), .c ({signal_10304, signal_4455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6675 ( .a ({signal_9904, signal_6528}), .b ({signal_10087, signal_6697}), .c ({signal_10305, signal_3935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6676 ( .a ({signal_10090, signal_6700}), .b ({signal_10094, signal_6704}), .c ({signal_10306, signal_3936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6677 ( .a ({signal_10085, signal_6695}), .b ({signal_10092, signal_6702}), .c ({signal_10307, signal_6905}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6678 ( .a ({signal_9323, signal_6039}), .b ({signal_9987, signal_6706}), .c ({signal_10196, signal_6906}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6679 ( .a ({signal_9325, signal_6041}), .b ({signal_9987, signal_6706}), .c ({signal_10197, signal_6907}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6680 ( .a ({signal_9646, signal_6368}), .b ({signal_9987, signal_6706}), .c ({signal_10198, signal_6908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6681 ( .a ({signal_9646, signal_6368}), .b ({signal_9989, signal_6708}), .c ({signal_10199, signal_6909}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6682 ( .a ({signal_9818, signal_6535}), .b ({signal_9990, signal_6709}), .c ({signal_10200, signal_6910}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6683 ( .a ({signal_9988, signal_6707}), .b ({signal_9991, signal_6710}), .c ({signal_10201, signal_6911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6684 ( .a ({signal_9989, signal_6708}), .b ({signal_9990, signal_6709}), .c ({signal_10202, signal_6912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6685 ( .a ({signal_9647, signal_6369}), .b ({signal_9991, signal_6710}), .c ({signal_10203, signal_6913}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6686 ( .a ({signal_9817, signal_6534}), .b ({signal_9992, signal_6711}), .c ({signal_10204, signal_6914}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6687 ( .a ({signal_9819, signal_6536}), .b ({signal_9992, signal_6711}), .c ({signal_10205, signal_6915}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6688 ( .a ({signal_9988, signal_6707}), .b ({signal_9995, signal_6714}), .c ({signal_10206, signal_6916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6689 ( .a ({signal_9331, signal_6047}), .b ({signal_9996, signal_6715}), .c ({signal_10207, signal_6917}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6690 ( .a ({signal_9333, signal_6049}), .b ({signal_9996, signal_6715}), .c ({signal_10208, signal_6918}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6691 ( .a ({signal_9650, signal_6372}), .b ({signal_9996, signal_6715}), .c ({signal_10209, signal_6919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6692 ( .a ({signal_9650, signal_6372}), .b ({signal_9998, signal_6717}), .c ({signal_10210, signal_6920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6693 ( .a ({signal_9826, signal_6543}), .b ({signal_9999, signal_6718}), .c ({signal_10211, signal_6921}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6694 ( .a ({signal_9997, signal_6716}), .b ({signal_10000, signal_6719}), .c ({signal_10212, signal_6922}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6695 ( .a ({signal_9998, signal_6717}), .b ({signal_9999, signal_6718}), .c ({signal_10213, signal_6923}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6696 ( .a ({signal_9651, signal_6373}), .b ({signal_10000, signal_6719}), .c ({signal_10214, signal_6924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6697 ( .a ({signal_9825, signal_6542}), .b ({signal_10001, signal_6720}), .c ({signal_10215, signal_6925}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6698 ( .a ({signal_9827, signal_6544}), .b ({signal_10001, signal_6720}), .c ({signal_10216, signal_6926}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6699 ( .a ({signal_9997, signal_6716}), .b ({signal_10004, signal_6723}), .c ({signal_10217, signal_6927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6700 ( .a ({signal_9339, signal_6055}), .b ({signal_10005, signal_6724}), .c ({signal_10218, signal_6928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6701 ( .a ({signal_9341, signal_6057}), .b ({signal_10005, signal_6724}), .c ({signal_10219, signal_6929}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6702 ( .a ({signal_9654, signal_6376}), .b ({signal_10005, signal_6724}), .c ({signal_10220, signal_6930}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6703 ( .a ({signal_9654, signal_6376}), .b ({signal_10007, signal_6726}), .c ({signal_10221, signal_6931}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6704 ( .a ({signal_9834, signal_6551}), .b ({signal_10008, signal_6727}), .c ({signal_10222, signal_6932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6705 ( .a ({signal_10006, signal_6725}), .b ({signal_10009, signal_6728}), .c ({signal_10223, signal_6933}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6706 ( .a ({signal_10007, signal_6726}), .b ({signal_10008, signal_6727}), .c ({signal_10224, signal_6934}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6707 ( .a ({signal_9655, signal_6377}), .b ({signal_10009, signal_6728}), .c ({signal_10225, signal_6935}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6708 ( .a ({signal_9833, signal_6550}), .b ({signal_10010, signal_6729}), .c ({signal_10226, signal_6936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6709 ( .a ({signal_9835, signal_6552}), .b ({signal_10010, signal_6729}), .c ({signal_10227, signal_6937}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6710 ( .a ({signal_10006, signal_6725}), .b ({signal_10013, signal_6732}), .c ({signal_10228, signal_6938}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6711 ( .a ({signal_9907, signal_6555}), .b ({signal_10100, signal_6737}), .c ({signal_10308, signal_4428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6712 ( .a ({signal_10097, signal_6734}), .b ({signal_10102, signal_6739}), .c ({signal_10309, signal_6939}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6713 ( .a ({signal_9912, signal_6560}), .b ({signal_10104, signal_6741}), .c ({signal_10310, signal_6940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6714 ( .a ({signal_9907, signal_6555}), .b ({signal_10099, signal_6736}), .c ({signal_10311, signal_4423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6715 ( .a ({signal_9913, signal_6561}), .b ({signal_10098, signal_6735}), .c ({signal_10312, signal_3903}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6716 ( .a ({signal_10101, signal_6738}), .b ({signal_10105, signal_6742}), .c ({signal_10313, signal_3904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6717 ( .a ({signal_10096, signal_6733}), .b ({signal_10103, signal_6740}), .c ({signal_10314, signal_6941}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6718 ( .a ({signal_9347, signal_6071}), .b ({signal_10014, signal_6744}), .c ({signal_10229, signal_6942}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6719 ( .a ({signal_9349, signal_6073}), .b ({signal_10014, signal_6744}), .c ({signal_10230, signal_6943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6720 ( .a ({signal_9658, signal_6388}), .b ({signal_10014, signal_6744}), .c ({signal_10231, signal_6944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6721 ( .a ({signal_9658, signal_6388}), .b ({signal_10016, signal_6746}), .c ({signal_10232, signal_6945}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6722 ( .a ({signal_9842, signal_6568}), .b ({signal_10017, signal_6747}), .c ({signal_10233, signal_6946}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6723 ( .a ({signal_10015, signal_6745}), .b ({signal_10018, signal_6748}), .c ({signal_10234, signal_6947}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6724 ( .a ({signal_10016, signal_6746}), .b ({signal_10017, signal_6747}), .c ({signal_10235, signal_6948}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6725 ( .a ({signal_9659, signal_6389}), .b ({signal_10018, signal_6748}), .c ({signal_10236, signal_6949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6726 ( .a ({signal_9841, signal_6567}), .b ({signal_10019, signal_6749}), .c ({signal_10237, signal_6950}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6727 ( .a ({signal_9843, signal_6569}), .b ({signal_10019, signal_6749}), .c ({signal_10238, signal_6951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6728 ( .a ({signal_10015, signal_6745}), .b ({signal_10022, signal_6752}), .c ({signal_10239, signal_6952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6729 ( .a ({signal_9355, signal_6079}), .b ({signal_10023, signal_6753}), .c ({signal_10240, signal_6953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6730 ( .a ({signal_9357, signal_6081}), .b ({signal_10023, signal_6753}), .c ({signal_10241, signal_6954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6731 ( .a ({signal_9662, signal_6392}), .b ({signal_10023, signal_6753}), .c ({signal_10242, signal_6955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6732 ( .a ({signal_9662, signal_6392}), .b ({signal_10025, signal_6755}), .c ({signal_10243, signal_6956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6733 ( .a ({signal_9850, signal_6576}), .b ({signal_10026, signal_6756}), .c ({signal_10244, signal_6957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6734 ( .a ({signal_10024, signal_6754}), .b ({signal_10027, signal_6757}), .c ({signal_10245, signal_6958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6735 ( .a ({signal_10025, signal_6755}), .b ({signal_10026, signal_6756}), .c ({signal_10246, signal_6959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6736 ( .a ({signal_9663, signal_6393}), .b ({signal_10027, signal_6757}), .c ({signal_10247, signal_6960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6737 ( .a ({signal_9849, signal_6575}), .b ({signal_10028, signal_6758}), .c ({signal_10248, signal_6961}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6738 ( .a ({signal_9851, signal_6577}), .b ({signal_10028, signal_6758}), .c ({signal_10249, signal_6962}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6739 ( .a ({signal_10024, signal_6754}), .b ({signal_10031, signal_6761}), .c ({signal_10250, signal_6963}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6740 ( .a ({signal_9363, signal_6087}), .b ({signal_10032, signal_6762}), .c ({signal_10251, signal_6964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6741 ( .a ({signal_9365, signal_6089}), .b ({signal_10032, signal_6762}), .c ({signal_10252, signal_6965}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6742 ( .a ({signal_9666, signal_6396}), .b ({signal_10032, signal_6762}), .c ({signal_10253, signal_6966}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6743 ( .a ({signal_9666, signal_6396}), .b ({signal_10034, signal_6764}), .c ({signal_10254, signal_6967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6744 ( .a ({signal_9858, signal_6584}), .b ({signal_10035, signal_6765}), .c ({signal_10255, signal_6968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6745 ( .a ({signal_10033, signal_6763}), .b ({signal_10036, signal_6766}), .c ({signal_10256, signal_6969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6746 ( .a ({signal_10034, signal_6764}), .b ({signal_10035, signal_6765}), .c ({signal_10257, signal_6970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6747 ( .a ({signal_9667, signal_6397}), .b ({signal_10036, signal_6766}), .c ({signal_10258, signal_6971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6748 ( .a ({signal_9857, signal_6583}), .b ({signal_10037, signal_6767}), .c ({signal_10259, signal_6972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6749 ( .a ({signal_9859, signal_6585}), .b ({signal_10037, signal_6767}), .c ({signal_10260, signal_6973}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6750 ( .a ({signal_10033, signal_6763}), .b ({signal_10040, signal_6770}), .c ({signal_10261, signal_6974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6751 ( .a ({signal_9916, signal_6588}), .b ({signal_10111, signal_6775}), .c ({signal_10315, signal_4396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6752 ( .a ({signal_10108, signal_6772}), .b ({signal_10113, signal_6777}), .c ({signal_10316, signal_6975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6753 ( .a ({signal_9921, signal_6593}), .b ({signal_10115, signal_6779}), .c ({signal_10317, signal_6976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6754 ( .a ({signal_9916, signal_6588}), .b ({signal_10110, signal_6774}), .c ({signal_10318, signal_4391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6755 ( .a ({signal_9922, signal_6594}), .b ({signal_10109, signal_6773}), .c ({signal_10319, signal_3871}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6756 ( .a ({signal_10112, signal_6776}), .b ({signal_10116, signal_6780}), .c ({signal_10320, signal_3872}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6757 ( .a ({signal_10107, signal_6771}), .b ({signal_10114, signal_6778}), .c ({signal_10321, signal_6977}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6758 ( .a ({signal_7571, signal_4266}), .b ({signal_10062, signal_6803}), .c ({signal_10262, signal_6978}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6759 ( .a ({signal_7544, signal_4274}), .b ({signal_10073, signal_6814}), .c ({signal_10263, signal_6979}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6760 ( .a ({signal_7826, signal_4282}), .b ({signal_10084, signal_6825}), .c ({signal_10264, signal_6980}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6761 ( .a ({signal_9862, signal_6597}), .b ({signal_10045, signal_6786}), .c ({signal_10265, signal_3116}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6762 ( .a ({signal_10042, signal_6783}), .b ({signal_10047, signal_6788}), .c ({signal_10266, signal_6981}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6763 ( .a ({signal_9867, signal_6602}), .b ({signal_10049, signal_6790}), .c ({signal_10267, signal_6982}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6764 ( .a ({signal_9862, signal_6597}), .b ({signal_10044, signal_6785}), .c ({signal_10268, signal_3113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6765 ( .a ({signal_9868, signal_6603}), .b ({signal_10043, signal_6784}), .c ({signal_10269, signal_3112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6766 ( .a ({signal_10046, signal_6787}), .b ({signal_10050, signal_6791}), .c ({signal_10270, signal_3111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6767 ( .a ({signal_10041, signal_6782}), .b ({signal_10048, signal_6789}), .c ({signal_10271, signal_6983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6768 ( .a ({signal_9871, signal_6606}), .b ({signal_10056, signal_6797}), .c ({signal_10272, signal_6984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6769 ( .a ({signal_10053, signal_6794}), .b ({signal_10058, signal_6799}), .c ({signal_10273, signal_6985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6770 ( .a ({signal_9876, signal_6611}), .b ({signal_10060, signal_6801}), .c ({signal_10274, signal_6986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6771 ( .a ({signal_9871, signal_6606}), .b ({signal_10055, signal_6796}), .c ({signal_10275, signal_6987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6772 ( .a ({signal_9877, signal_6612}), .b ({signal_10054, signal_6795}), .c ({signal_10276, signal_6988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6773 ( .a ({signal_10057, signal_6798}), .b ({signal_10061, signal_6802}), .c ({signal_10277, signal_6989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6774 ( .a ({signal_10052, signal_6793}), .b ({signal_10059, signal_6800}), .c ({signal_10278, signal_6990}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6775 ( .a ({signal_9880, signal_6615}), .b ({signal_10067, signal_6808}), .c ({signal_10279, signal_6991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6776 ( .a ({signal_10064, signal_6805}), .b ({signal_10069, signal_6810}), .c ({signal_10280, signal_6992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6777 ( .a ({signal_9885, signal_6620}), .b ({signal_10071, signal_6812}), .c ({signal_10281, signal_6993}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6778 ( .a ({signal_9880, signal_6615}), .b ({signal_10066, signal_6807}), .c ({signal_10282, signal_6994}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6779 ( .a ({signal_9886, signal_6621}), .b ({signal_10065, signal_6806}), .c ({signal_10283, signal_6995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6780 ( .a ({signal_10068, signal_6809}), .b ({signal_10072, signal_6813}), .c ({signal_10284, signal_6996}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6781 ( .a ({signal_10063, signal_6804}), .b ({signal_10070, signal_6811}), .c ({signal_10285, signal_6997}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6782 ( .a ({signal_9889, signal_6624}), .b ({signal_10078, signal_6819}), .c ({signal_10286, signal_6998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6783 ( .a ({signal_10075, signal_6816}), .b ({signal_10080, signal_6821}), .c ({signal_10287, signal_6999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6784 ( .a ({signal_9894, signal_6629}), .b ({signal_10082, signal_6823}), .c ({signal_10288, signal_7000}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6785 ( .a ({signal_9889, signal_6624}), .b ({signal_10077, signal_6818}), .c ({signal_10289, signal_7001}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6786 ( .a ({signal_9895, signal_6630}), .b ({signal_10076, signal_6817}), .c ({signal_10290, signal_7002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6787 ( .a ({signal_10079, signal_6820}), .b ({signal_10083, signal_6824}), .c ({signal_10291, signal_7003}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6788 ( .a ({signal_10074, signal_6815}), .b ({signal_10081, signal_6822}), .c ({signal_10292, signal_7004}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6789 ( .a ({signal_10129, signal_6836}), .b ({signal_10322, signal_3898}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6790 ( .a ({signal_10140, signal_6847}), .b ({signal_10323, signal_3922}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6791 ( .a ({signal_10151, signal_6858}), .b ({signal_10324, signal_3946}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6792 ( .a ({signal_10162, signal_6869}), .b ({signal_10325, signal_3970}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6793 ( .a ({signal_10173, signal_6880}), .b ({signal_10326, signal_3994}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6794 ( .a ({signal_10184, signal_6891}), .b ({signal_10327, signal_3890}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6795 ( .a ({signal_10195, signal_6902}), .b ({signal_10328, signal_3914}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6796 ( .a ({signal_10302, signal_6903}), .b ({signal_10494, signal_4453}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6797 ( .a ({signal_10303, signal_6904}), .b ({signal_10495, signal_4454}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6798 ( .a ({signal_10307, signal_6905}), .b ({signal_10496, signal_4458}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6799 ( .a ({signal_10206, signal_6916}), .b ({signal_10329, signal_3962}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6800 ( .a ({signal_10217, signal_6927}), .b ({signal_10330, signal_3986}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6801 ( .a ({signal_10228, signal_6938}), .b ({signal_10331, signal_3882}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6802 ( .a ({signal_10309, signal_6939}), .b ({signal_10497, signal_4421}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6803 ( .a ({signal_10310, signal_6940}), .b ({signal_10498, signal_4422}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6804 ( .a ({signal_10314, signal_6941}), .b ({signal_10499, signal_4426}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6805 ( .a ({signal_10239, signal_6952}), .b ({signal_10332, signal_3930}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6806 ( .a ({signal_10250, signal_6963}), .b ({signal_10333, signal_3954}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6807 ( .a ({signal_10261, signal_6974}), .b ({signal_10334, signal_3978}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6808 ( .a ({signal_10316, signal_6975}), .b ({signal_10500, signal_4389}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6809 ( .a ({signal_10317, signal_6976}), .b ({signal_10501, signal_4390}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6810 ( .a ({signal_10321, signal_6977}), .b ({signal_10502, signal_4394}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6811 ( .a ({signal_10262, signal_6978}), .b ({signal_10335, signal_4138}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6812 ( .a ({signal_10263, signal_6979}), .b ({signal_10336, signal_4146}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6813 ( .a ({signal_10264, signal_6980}), .b ({signal_10337, signal_4154}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6814 ( .a ({signal_10266, signal_6981}), .b ({signal_10338, signal_3115}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6815 ( .a ({signal_10267, signal_6982}), .b ({signal_10339, signal_3114}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6816 ( .a ({signal_10271, signal_6983}), .b ({signal_10340, signal_3110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6817 ( .a ({signal_9925, signal_6633}), .b ({signal_10123, signal_6830}), .c ({signal_10341, signal_4420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6818 ( .a ({signal_10120, signal_6827}), .b ({signal_10125, signal_6832}), .c ({signal_10342, signal_7005}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6819 ( .a ({signal_9930, signal_6638}), .b ({signal_10127, signal_6834}), .c ({signal_10343, signal_7006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6820 ( .a ({signal_9925, signal_6633}), .b ({signal_10122, signal_6829}), .c ({signal_10344, signal_4415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6821 ( .a ({signal_9931, signal_6639}), .b ({signal_10121, signal_6828}), .c ({signal_10345, signal_3895}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6822 ( .a ({signal_10124, signal_6831}), .b ({signal_10128, signal_6835}), .c ({signal_10346, signal_3896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6823 ( .a ({signal_10119, signal_6826}), .b ({signal_10126, signal_6833}), .c ({signal_10347, signal_7007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6824 ( .a ({signal_9934, signal_6642}), .b ({signal_10134, signal_6841}), .c ({signal_10348, signal_4444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6825 ( .a ({signal_10131, signal_6838}), .b ({signal_10136, signal_6843}), .c ({signal_10349, signal_7008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6826 ( .a ({signal_9939, signal_6647}), .b ({signal_10138, signal_6845}), .c ({signal_10350, signal_7009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6827 ( .a ({signal_9934, signal_6642}), .b ({signal_10133, signal_6840}), .c ({signal_10351, signal_4439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6828 ( .a ({signal_9940, signal_6648}), .b ({signal_10132, signal_6839}), .c ({signal_10352, signal_3919}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6829 ( .a ({signal_10135, signal_6842}), .b ({signal_10139, signal_6846}), .c ({signal_10353, signal_3920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6830 ( .a ({signal_10130, signal_6837}), .b ({signal_10137, signal_6844}), .c ({signal_10354, signal_7010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6831 ( .a ({signal_9943, signal_6651}), .b ({signal_10145, signal_6852}), .c ({signal_10355, signal_4468}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6832 ( .a ({signal_10142, signal_6849}), .b ({signal_10147, signal_6854}), .c ({signal_10356, signal_7011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6833 ( .a ({signal_9948, signal_6656}), .b ({signal_10149, signal_6856}), .c ({signal_10357, signal_7012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6834 ( .a ({signal_9943, signal_6651}), .b ({signal_10144, signal_6851}), .c ({signal_10358, signal_4463}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6835 ( .a ({signal_9949, signal_6657}), .b ({signal_10143, signal_6850}), .c ({signal_10359, signal_3943}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6836 ( .a ({signal_10146, signal_6853}), .b ({signal_10150, signal_6857}), .c ({signal_10360, signal_3944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6837 ( .a ({signal_10141, signal_6848}), .b ({signal_10148, signal_6855}), .c ({signal_10361, signal_7013}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6838 ( .a ({signal_9952, signal_6660}), .b ({signal_10156, signal_6863}), .c ({signal_10362, signal_4492}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6839 ( .a ({signal_10153, signal_6860}), .b ({signal_10158, signal_6865}), .c ({signal_10363, signal_7014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6840 ( .a ({signal_9957, signal_6665}), .b ({signal_10160, signal_6867}), .c ({signal_10364, signal_7015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6841 ( .a ({signal_9952, signal_6660}), .b ({signal_10155, signal_6862}), .c ({signal_10365, signal_4487}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6842 ( .a ({signal_9958, signal_6666}), .b ({signal_10154, signal_6861}), .c ({signal_10366, signal_3967}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6843 ( .a ({signal_10157, signal_6864}), .b ({signal_10161, signal_6868}), .c ({signal_10367, signal_3968}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6844 ( .a ({signal_10152, signal_6859}), .b ({signal_10159, signal_6866}), .c ({signal_10368, signal_7016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6845 ( .a ({signal_9961, signal_6669}), .b ({signal_10167, signal_6874}), .c ({signal_10369, signal_4516}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6846 ( .a ({signal_10164, signal_6871}), .b ({signal_10169, signal_6876}), .c ({signal_10370, signal_7017}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6847 ( .a ({signal_9966, signal_6674}), .b ({signal_10171, signal_6878}), .c ({signal_10371, signal_7018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6848 ( .a ({signal_9961, signal_6669}), .b ({signal_10166, signal_6873}), .c ({signal_10372, signal_4511}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6849 ( .a ({signal_9967, signal_6675}), .b ({signal_10165, signal_6872}), .c ({signal_10373, signal_3991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6850 ( .a ({signal_10168, signal_6875}), .b ({signal_10172, signal_6879}), .c ({signal_10374, signal_3992}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6851 ( .a ({signal_10163, signal_6870}), .b ({signal_10170, signal_6877}), .c ({signal_10375, signal_7019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6852 ( .a ({signal_9970, signal_6678}), .b ({signal_10178, signal_6885}), .c ({signal_10376, signal_4412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6853 ( .a ({signal_10175, signal_6882}), .b ({signal_10180, signal_6887}), .c ({signal_10377, signal_7020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6854 ( .a ({signal_9975, signal_6683}), .b ({signal_10182, signal_6889}), .c ({signal_10378, signal_7021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6855 ( .a ({signal_9970, signal_6678}), .b ({signal_10177, signal_6884}), .c ({signal_10379, signal_4407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6856 ( .a ({signal_9976, signal_6684}), .b ({signal_10176, signal_6883}), .c ({signal_10380, signal_3887}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6857 ( .a ({signal_10179, signal_6886}), .b ({signal_10183, signal_6890}), .c ({signal_10381, signal_3888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6858 ( .a ({signal_10174, signal_6881}), .b ({signal_10181, signal_6888}), .c ({signal_10382, signal_7022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6859 ( .a ({signal_9979, signal_6687}), .b ({signal_10189, signal_6896}), .c ({signal_10383, signal_4436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6860 ( .a ({signal_10186, signal_6893}), .b ({signal_10191, signal_6898}), .c ({signal_10384, signal_7023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6861 ( .a ({signal_9984, signal_6692}), .b ({signal_10193, signal_6900}), .c ({signal_10385, signal_7024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6862 ( .a ({signal_9979, signal_6687}), .b ({signal_10188, signal_6895}), .c ({signal_10386, signal_4431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6863 ( .a ({signal_9985, signal_6693}), .b ({signal_10187, signal_6894}), .c ({signal_10387, signal_3911}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6864 ( .a ({signal_10190, signal_6897}), .b ({signal_10194, signal_6901}), .c ({signal_10388, signal_3912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6865 ( .a ({signal_10185, signal_6892}), .b ({signal_10192, signal_6899}), .c ({signal_10389, signal_7025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6866 ( .a ({signal_9988, signal_6707}), .b ({signal_10200, signal_6910}), .c ({signal_10390, signal_4484}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6867 ( .a ({signal_10197, signal_6907}), .b ({signal_10202, signal_6912}), .c ({signal_10391, signal_7026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6868 ( .a ({signal_9993, signal_6712}), .b ({signal_10204, signal_6914}), .c ({signal_10392, signal_7027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6869 ( .a ({signal_9988, signal_6707}), .b ({signal_10199, signal_6909}), .c ({signal_10393, signal_4479}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6870 ( .a ({signal_9994, signal_6713}), .b ({signal_10198, signal_6908}), .c ({signal_10394, signal_3959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6871 ( .a ({signal_10201, signal_6911}), .b ({signal_10205, signal_6915}), .c ({signal_10395, signal_3960}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6872 ( .a ({signal_10196, signal_6906}), .b ({signal_10203, signal_6913}), .c ({signal_10396, signal_7028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6873 ( .a ({signal_9997, signal_6716}), .b ({signal_10211, signal_6921}), .c ({signal_10397, signal_4508}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6874 ( .a ({signal_10208, signal_6918}), .b ({signal_10213, signal_6923}), .c ({signal_10398, signal_7029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6875 ( .a ({signal_10002, signal_6721}), .b ({signal_10215, signal_6925}), .c ({signal_10399, signal_7030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6876 ( .a ({signal_9997, signal_6716}), .b ({signal_10210, signal_6920}), .c ({signal_10400, signal_4503}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6877 ( .a ({signal_10003, signal_6722}), .b ({signal_10209, signal_6919}), .c ({signal_10401, signal_3983}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6878 ( .a ({signal_10212, signal_6922}), .b ({signal_10216, signal_6926}), .c ({signal_10402, signal_3984}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6879 ( .a ({signal_10207, signal_6917}), .b ({signal_10214, signal_6924}), .c ({signal_10403, signal_7031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6880 ( .a ({signal_10006, signal_6725}), .b ({signal_10222, signal_6932}), .c ({signal_10404, signal_4404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6881 ( .a ({signal_10219, signal_6929}), .b ({signal_10224, signal_6934}), .c ({signal_10405, signal_7032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6882 ( .a ({signal_10011, signal_6730}), .b ({signal_10226, signal_6936}), .c ({signal_10406, signal_7033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6883 ( .a ({signal_10006, signal_6725}), .b ({signal_10221, signal_6931}), .c ({signal_10407, signal_4399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6884 ( .a ({signal_10012, signal_6731}), .b ({signal_10220, signal_6930}), .c ({signal_10408, signal_3879}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6885 ( .a ({signal_10223, signal_6933}), .b ({signal_10227, signal_6937}), .c ({signal_10409, signal_3880}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6886 ( .a ({signal_10218, signal_6928}), .b ({signal_10225, signal_6935}), .c ({signal_10410, signal_7034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6887 ( .a ({signal_10015, signal_6745}), .b ({signal_10233, signal_6946}), .c ({signal_10411, signal_4452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6888 ( .a ({signal_10230, signal_6943}), .b ({signal_10235, signal_6948}), .c ({signal_10412, signal_7035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6889 ( .a ({signal_10020, signal_6750}), .b ({signal_10237, signal_6950}), .c ({signal_10413, signal_7036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6890 ( .a ({signal_10015, signal_6745}), .b ({signal_10232, signal_6945}), .c ({signal_10414, signal_4447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6891 ( .a ({signal_10021, signal_6751}), .b ({signal_10231, signal_6944}), .c ({signal_10415, signal_3927}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6892 ( .a ({signal_10234, signal_6947}), .b ({signal_10238, signal_6951}), .c ({signal_10416, signal_3928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6893 ( .a ({signal_10229, signal_6942}), .b ({signal_10236, signal_6949}), .c ({signal_10417, signal_7037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6894 ( .a ({signal_10024, signal_6754}), .b ({signal_10244, signal_6957}), .c ({signal_10418, signal_4476}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6895 ( .a ({signal_10241, signal_6954}), .b ({signal_10246, signal_6959}), .c ({signal_10419, signal_7038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6896 ( .a ({signal_10029, signal_6759}), .b ({signal_10248, signal_6961}), .c ({signal_10420, signal_7039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6897 ( .a ({signal_10024, signal_6754}), .b ({signal_10243, signal_6956}), .c ({signal_10421, signal_4471}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6898 ( .a ({signal_10030, signal_6760}), .b ({signal_10242, signal_6955}), .c ({signal_10422, signal_3951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6899 ( .a ({signal_10245, signal_6958}), .b ({signal_10249, signal_6962}), .c ({signal_10423, signal_3952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6900 ( .a ({signal_10240, signal_6953}), .b ({signal_10247, signal_6960}), .c ({signal_10424, signal_7040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6901 ( .a ({signal_10033, signal_6763}), .b ({signal_10255, signal_6968}), .c ({signal_10425, signal_4500}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6902 ( .a ({signal_10252, signal_6965}), .b ({signal_10257, signal_6970}), .c ({signal_10426, signal_7041}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6903 ( .a ({signal_10038, signal_6768}), .b ({signal_10259, signal_6972}), .c ({signal_10427, signal_7042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6904 ( .a ({signal_10033, signal_6763}), .b ({signal_10254, signal_6967}), .c ({signal_10428, signal_4495}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6905 ( .a ({signal_10039, signal_6769}), .b ({signal_10253, signal_6966}), .c ({signal_10429, signal_3975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6906 ( .a ({signal_10256, signal_6969}), .b ({signal_10260, signal_6973}), .c ({signal_10430, signal_3976}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6907 ( .a ({signal_10251, signal_6964}), .b ({signal_10258, signal_6971}), .c ({signal_10431, signal_7043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6908 ( .a ({signal_10228, signal_6938}), .b ({signal_10315, signal_4396}), .c ({signal_10503, signal_7044}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6909 ( .a ({signal_10315, signal_4396}), .b ({signal_10319, signal_3871}), .c ({signal_10504, signal_7045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6910 ( .a ({signal_10315, signal_4396}), .b ({signal_10320, signal_3872}), .c ({signal_10505, signal_7046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6911 ( .a ({signal_10117, signal_6781}), .b ({signal_10315, signal_4396}), .c ({signal_10506, signal_7047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6912 ( .a ({signal_10195, signal_6902}), .b ({signal_10308, signal_4428}), .c ({signal_10507, signal_7048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6913 ( .a ({signal_10308, signal_4428}), .b ({signal_10312, signal_3903}), .c ({signal_10508, signal_7049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6914 ( .a ({signal_10308, signal_4428}), .b ({signal_10313, signal_3904}), .c ({signal_10509, signal_7050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6915 ( .a ({signal_10106, signal_6743}), .b ({signal_10308, signal_4428}), .c ({signal_10510, signal_7051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6916 ( .a ({signal_10151, signal_6858}), .b ({signal_10301, signal_4460}), .c ({signal_10511, signal_7052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6917 ( .a ({signal_10301, signal_4460}), .b ({signal_10305, signal_3935}), .c ({signal_10512, signal_7053}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6918 ( .a ({signal_10301, signal_4460}), .b ({signal_10306, signal_3936}), .c ({signal_10513, signal_7054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6919 ( .a ({signal_10095, signal_6705}), .b ({signal_10301, signal_4460}), .c ({signal_10514, signal_7055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6920 ( .a ({signal_7772, signal_4306}), .b ({signal_10263, signal_6979}), .c ({signal_10432, signal_7056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6921 ( .a ({signal_7835, signal_4279}), .b ({signal_10290, signal_7002}), .c ({signal_10433, signal_4151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6922 ( .a ({signal_7832, signal_4280}), .b ({signal_10291, signal_7003}), .c ({signal_10434, signal_4152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6923 ( .a ({signal_7829, signal_4281}), .b ({signal_10292, signal_7004}), .c ({signal_10435, signal_7057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6924 ( .a ({signal_7799, signal_4298}), .b ({signal_10262, signal_6978}), .c ({signal_10436, signal_7058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6925 ( .a ({signal_7592, signal_4259}), .b ({signal_10272, signal_6984}), .c ({signal_10437, signal_4131}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6926 ( .a ({signal_7589, signal_4260}), .b ({signal_10273, signal_6985}), .c ({signal_10438, signal_7059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6927 ( .a ({signal_7586, signal_4261}), .b ({signal_10274, signal_6986}), .c ({signal_10439, signal_7060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6928 ( .a ({signal_7583, signal_4262}), .b ({signal_10275, signal_6987}), .c ({signal_10440, signal_4134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6929 ( .a ({signal_7580, signal_4263}), .b ({signal_10276, signal_6988}), .c ({signal_10441, signal_4135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6930 ( .a ({signal_7577, signal_4264}), .b ({signal_10277, signal_6989}), .c ({signal_10442, signal_4136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6931 ( .a ({signal_7574, signal_4265}), .b ({signal_10278, signal_6990}), .c ({signal_10443, signal_7061}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6932 ( .a ({signal_7568, signal_4267}), .b ({signal_10279, signal_6991}), .c ({signal_10444, signal_4139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6933 ( .a ({signal_7565, signal_4268}), .b ({signal_10280, signal_6992}), .c ({signal_10445, signal_7062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6934 ( .a ({signal_7559, signal_4269}), .b ({signal_10281, signal_6993}), .c ({signal_10446, signal_7063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6935 ( .a ({signal_7556, signal_4270}), .b ({signal_10282, signal_6994}), .c ({signal_10447, signal_4142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6936 ( .a ({signal_7553, signal_4271}), .b ({signal_10283, signal_6995}), .c ({signal_10448, signal_4143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6937 ( .a ({signal_7550, signal_4272}), .b ({signal_10284, signal_6996}), .c ({signal_10449, signal_4144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6938 ( .a ({signal_7547, signal_4273}), .b ({signal_10285, signal_6997}), .c ({signal_10450, signal_7064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6939 ( .a ({signal_7541, signal_4275}), .b ({signal_10286, signal_6998}), .c ({signal_10451, signal_4147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6940 ( .a ({signal_7538, signal_4276}), .b ({signal_10287, signal_6999}), .c ({signal_10452, signal_7065}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6941 ( .a ({signal_7535, signal_4277}), .b ({signal_10288, signal_7000}), .c ({signal_10453, signal_7066}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6942 ( .a ({signal_7532, signal_4278}), .b ({signal_10289, signal_7001}), .c ({signal_10454, signal_4150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6943 ( .a ({signal_7745, signal_4314}), .b ({signal_10264, signal_6980}), .c ({signal_10455, signal_7067}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6944 ( .a ({signal_10342, signal_7005}), .b ({signal_10515, signal_4413}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6945 ( .a ({signal_10343, signal_7006}), .b ({signal_10516, signal_4414}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6946 ( .a ({signal_10347, signal_7007}), .b ({signal_10517, signal_4418}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6947 ( .a ({signal_10349, signal_7008}), .b ({signal_10518, signal_4437}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6948 ( .a ({signal_10350, signal_7009}), .b ({signal_10519, signal_4438}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6949 ( .a ({signal_10354, signal_7010}), .b ({signal_10520, signal_4442}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6950 ( .a ({signal_10356, signal_7011}), .b ({signal_10521, signal_4461}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6951 ( .a ({signal_10357, signal_7012}), .b ({signal_10522, signal_4462}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6952 ( .a ({signal_10361, signal_7013}), .b ({signal_10523, signal_4466}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6953 ( .a ({signal_10363, signal_7014}), .b ({signal_10524, signal_4485}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6954 ( .a ({signal_10364, signal_7015}), .b ({signal_10525, signal_4486}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6955 ( .a ({signal_10368, signal_7016}), .b ({signal_10526, signal_4490}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6956 ( .a ({signal_10370, signal_7017}), .b ({signal_10527, signal_4509}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6957 ( .a ({signal_10371, signal_7018}), .b ({signal_10528, signal_4510}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6958 ( .a ({signal_10375, signal_7019}), .b ({signal_10529, signal_4514}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6959 ( .a ({signal_10377, signal_7020}), .b ({signal_10530, signal_4405}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6960 ( .a ({signal_10378, signal_7021}), .b ({signal_10531, signal_4406}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6961 ( .a ({signal_10382, signal_7022}), .b ({signal_10532, signal_4410}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6962 ( .a ({signal_10384, signal_7023}), .b ({signal_10533, signal_4429}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6963 ( .a ({signal_10385, signal_7024}), .b ({signal_10534, signal_4430}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6964 ( .a ({signal_10389, signal_7025}), .b ({signal_10535, signal_4434}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6965 ( .a ({signal_10391, signal_7026}), .b ({signal_10536, signal_4477}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6966 ( .a ({signal_10392, signal_7027}), .b ({signal_10537, signal_4478}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6967 ( .a ({signal_10396, signal_7028}), .b ({signal_10538, signal_4482}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6968 ( .a ({signal_10398, signal_7029}), .b ({signal_10539, signal_4501}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6969 ( .a ({signal_10399, signal_7030}), .b ({signal_10540, signal_4502}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6970 ( .a ({signal_10403, signal_7031}), .b ({signal_10541, signal_4506}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6971 ( .a ({signal_10405, signal_7032}), .b ({signal_10542, signal_4397}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6972 ( .a ({signal_10406, signal_7033}), .b ({signal_10543, signal_4398}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6973 ( .a ({signal_10410, signal_7034}), .b ({signal_10544, signal_4402}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6974 ( .a ({signal_10412, signal_7035}), .b ({signal_10545, signal_4445}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6975 ( .a ({signal_10413, signal_7036}), .b ({signal_10546, signal_4446}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6976 ( .a ({signal_10417, signal_7037}), .b ({signal_10547, signal_4450}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6977 ( .a ({signal_10419, signal_7038}), .b ({signal_10548, signal_4469}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6978 ( .a ({signal_10420, signal_7039}), .b ({signal_10549, signal_4470}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6979 ( .a ({signal_10424, signal_7040}), .b ({signal_10550, signal_4474}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6980 ( .a ({signal_10426, signal_7041}), .b ({signal_10551, signal_4493}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6981 ( .a ({signal_10427, signal_7042}), .b ({signal_10552, signal_4494}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6982 ( .a ({signal_10431, signal_7043}), .b ({signal_10553, signal_4498}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6983 ( .a ({signal_10432, signal_7056}), .b ({signal_10554, signal_4178}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6984 ( .a ({signal_10435, signal_7057}), .b ({signal_10555, signal_4153}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6985 ( .a ({signal_10436, signal_7058}), .b ({signal_10556, signal_4170}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6986 ( .a ({signal_10438, signal_7059}), .b ({signal_10557, signal_4132}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6987 ( .a ({signal_10439, signal_7060}), .b ({signal_10558, signal_4133}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6988 ( .a ({signal_10443, signal_7061}), .b ({signal_10559, signal_4137}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6989 ( .a ({signal_10445, signal_7062}), .b ({signal_10560, signal_4140}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6990 ( .a ({signal_10446, signal_7063}), .b ({signal_10561, signal_4141}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6991 ( .a ({signal_10450, signal_7064}), .b ({signal_10562, signal_4145}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6992 ( .a ({signal_10452, signal_7065}), .b ({signal_10563, signal_4148}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6993 ( .a ({signal_10453, signal_7066}), .b ({signal_10564, signal_4149}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_6994 ( .a ({signal_10455, signal_7067}), .b ({signal_10565, signal_4186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6995 ( .a ({signal_10316, signal_6975}), .b ({signal_10404, signal_4404}), .c ({signal_10566, signal_7068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6996 ( .a ({signal_10317, signal_6976}), .b ({signal_10405, signal_7032}), .c ({signal_10567, signal_7069}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6997 ( .a ({signal_10318, signal_4391}), .b ({signal_10406, signal_7033}), .c ({signal_10568, signal_7070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6998 ( .a ({signal_10407, signal_4399}), .b ({signal_10504, signal_7045}), .c ({signal_10772, signal_7071}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_6999 ( .a ({signal_10408, signal_3879}), .b ({signal_10505, signal_7046}), .c ({signal_10773, signal_7072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7000 ( .a ({signal_10321, signal_6977}), .b ({signal_10409, signal_3880}), .c ({signal_10569, signal_7073}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7001 ( .a ({signal_10129, signal_6836}), .b ({signal_10503, signal_7044}), .c ({signal_10774, signal_7074}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7002 ( .a ({signal_10376, signal_4412}), .b ({signal_10405, signal_7032}), .c ({signal_10570, signal_7075}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7003 ( .a ({signal_10377, signal_7020}), .b ({signal_10406, signal_7033}), .c ({signal_10571, signal_7076}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7004 ( .a ({signal_10378, signal_7021}), .b ({signal_10407, signal_4399}), .c ({signal_10572, signal_7077}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7005 ( .a ({signal_10410, signal_7034}), .b ({signal_10506, signal_7047}), .c ({signal_10775, signal_7078}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7006 ( .a ({signal_10381, signal_3888}), .b ({signal_10410, signal_7034}), .c ({signal_10573, signal_7079}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7007 ( .a ({signal_10184, signal_6891}), .b ({signal_10404, signal_4404}), .c ({signal_10574, signal_7080}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7008 ( .a ({signal_10129, signal_6836}), .b ({signal_10376, signal_4412}), .c ({signal_10575, signal_7081}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7009 ( .a ({signal_10341, signal_4420}), .b ({signal_10377, signal_7020}), .c ({signal_10576, signal_7082}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7010 ( .a ({signal_10315, signal_4396}), .b ({signal_10342, signal_7005}), .c ({signal_10577, signal_7083}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7011 ( .a ({signal_10342, signal_7005}), .b ({signal_10378, signal_7021}), .c ({signal_10578, signal_7084}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7012 ( .a ({signal_10316, signal_6975}), .b ({signal_10343, signal_7006}), .c ({signal_10579, signal_7085}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7013 ( .a ({signal_10343, signal_7006}), .b ({signal_10379, signal_4407}), .c ({signal_10580, signal_7086}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7014 ( .a ({signal_10317, signal_6976}), .b ({signal_10344, signal_4415}), .c ({signal_10581, signal_7087}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7015 ( .a ({signal_10346, signal_3896}), .b ({signal_10382, signal_7022}), .c ({signal_10582, signal_7088}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7016 ( .a ({signal_10320, signal_3872}), .b ({signal_10347, signal_7007}), .c ({signal_10583, signal_7089}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7017 ( .a ({signal_10117, signal_6781}), .b ({signal_10341, signal_4420}), .c ({signal_10584, signal_7090}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7018 ( .a ({signal_10404, signal_4404}), .b ({signal_10408, signal_3879}), .c ({signal_10585, signal_7091}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7019 ( .a ({signal_10404, signal_4404}), .b ({signal_10409, signal_3880}), .c ({signal_10586, signal_7092}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7020 ( .a ({signal_10228, signal_6938}), .b ({signal_10404, signal_4404}), .c ({signal_10587, signal_7093}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7021 ( .a ({signal_10376, signal_4412}), .b ({signal_10380, signal_3887}), .c ({signal_10588, signal_7094}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7022 ( .a ({signal_10376, signal_4412}), .b ({signal_10381, signal_3888}), .c ({signal_10589, signal_7095}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7023 ( .a ({signal_10184, signal_6891}), .b ({signal_10376, signal_4412}), .c ({signal_10590, signal_7096}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7024 ( .a ({signal_10341, signal_4420}), .b ({signal_10345, signal_3895}), .c ({signal_10591, signal_7097}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7025 ( .a ({signal_10341, signal_4420}), .b ({signal_10346, signal_3896}), .c ({signal_10592, signal_7098}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7026 ( .a ({signal_10129, signal_6836}), .b ({signal_10341, signal_4420}), .c ({signal_10593, signal_7099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7027 ( .a ({signal_10309, signal_6939}), .b ({signal_10383, signal_4436}), .c ({signal_10594, signal_7100}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7028 ( .a ({signal_10310, signal_6940}), .b ({signal_10384, signal_7023}), .c ({signal_10595, signal_7101}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7029 ( .a ({signal_10311, signal_4423}), .b ({signal_10385, signal_7024}), .c ({signal_10596, signal_7102}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7030 ( .a ({signal_10386, signal_4431}), .b ({signal_10508, signal_7049}), .c ({signal_10776, signal_7103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7031 ( .a ({signal_10387, signal_3911}), .b ({signal_10509, signal_7050}), .c ({signal_10777, signal_7104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7032 ( .a ({signal_10314, signal_6941}), .b ({signal_10388, signal_3912}), .c ({signal_10597, signal_7105}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7033 ( .a ({signal_10239, signal_6952}), .b ({signal_10507, signal_7048}), .c ({signal_10778, signal_7106}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7034 ( .a ({signal_10348, signal_4444}), .b ({signal_10384, signal_7023}), .c ({signal_10598, signal_7107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7035 ( .a ({signal_10349, signal_7008}), .b ({signal_10385, signal_7024}), .c ({signal_10599, signal_7108}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7036 ( .a ({signal_10350, signal_7009}), .b ({signal_10386, signal_4431}), .c ({signal_10600, signal_7109}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7037 ( .a ({signal_10389, signal_7025}), .b ({signal_10510, signal_7051}), .c ({signal_10779, signal_7110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7038 ( .a ({signal_10353, signal_3920}), .b ({signal_10389, signal_7025}), .c ({signal_10601, signal_7111}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7039 ( .a ({signal_10140, signal_6847}), .b ({signal_10383, signal_4436}), .c ({signal_10602, signal_7112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7040 ( .a ({signal_10239, signal_6952}), .b ({signal_10348, signal_4444}), .c ({signal_10603, signal_7113}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7041 ( .a ({signal_10349, signal_7008}), .b ({signal_10411, signal_4452}), .c ({signal_10604, signal_7114}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7042 ( .a ({signal_10308, signal_4428}), .b ({signal_10412, signal_7035}), .c ({signal_10605, signal_7115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7043 ( .a ({signal_10350, signal_7009}), .b ({signal_10412, signal_7035}), .c ({signal_10606, signal_7116}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7044 ( .a ({signal_10309, signal_6939}), .b ({signal_10413, signal_7036}), .c ({signal_10607, signal_7117}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7045 ( .a ({signal_10351, signal_4439}), .b ({signal_10413, signal_7036}), .c ({signal_10608, signal_7118}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7046 ( .a ({signal_10310, signal_6940}), .b ({signal_10414, signal_4447}), .c ({signal_10609, signal_7119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7047 ( .a ({signal_10354, signal_7010}), .b ({signal_10416, signal_3928}), .c ({signal_10610, signal_7120}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7048 ( .a ({signal_10313, signal_3904}), .b ({signal_10417, signal_7037}), .c ({signal_10611, signal_7121}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7049 ( .a ({signal_10106, signal_6743}), .b ({signal_10411, signal_4452}), .c ({signal_10612, signal_7122}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7050 ( .a ({signal_10383, signal_4436}), .b ({signal_10387, signal_3911}), .c ({signal_10613, signal_7123}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7051 ( .a ({signal_10383, signal_4436}), .b ({signal_10388, signal_3912}), .c ({signal_10614, signal_7124}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7052 ( .a ({signal_10195, signal_6902}), .b ({signal_10383, signal_4436}), .c ({signal_10615, signal_7125}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7053 ( .a ({signal_10348, signal_4444}), .b ({signal_10352, signal_3919}), .c ({signal_10616, signal_7126}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7054 ( .a ({signal_10348, signal_4444}), .b ({signal_10353, signal_3920}), .c ({signal_10617, signal_7127}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7055 ( .a ({signal_10140, signal_6847}), .b ({signal_10348, signal_4444}), .c ({signal_10618, signal_7128}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7056 ( .a ({signal_10411, signal_4452}), .b ({signal_10415, signal_3927}), .c ({signal_10619, signal_7129}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7057 ( .a ({signal_10411, signal_4452}), .b ({signal_10416, signal_3928}), .c ({signal_10620, signal_7130}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7058 ( .a ({signal_10239, signal_6952}), .b ({signal_10411, signal_4452}), .c ({signal_10621, signal_7131}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7059 ( .a ({signal_10302, signal_6903}), .b ({signal_10355, signal_4468}), .c ({signal_10622, signal_7132}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7060 ( .a ({signal_10303, signal_6904}), .b ({signal_10356, signal_7011}), .c ({signal_10623, signal_7133}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7061 ( .a ({signal_10304, signal_4455}), .b ({signal_10357, signal_7012}), .c ({signal_10624, signal_7134}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7062 ( .a ({signal_10358, signal_4463}), .b ({signal_10512, signal_7053}), .c ({signal_10780, signal_7135}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7063 ( .a ({signal_10359, signal_3943}), .b ({signal_10513, signal_7054}), .c ({signal_10781, signal_7136}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7064 ( .a ({signal_10307, signal_6905}), .b ({signal_10360, signal_3944}), .c ({signal_10625, signal_7137}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7065 ( .a ({signal_10206, signal_6916}), .b ({signal_10511, signal_7052}), .c ({signal_10782, signal_7138}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7066 ( .a ({signal_10356, signal_7011}), .b ({signal_10418, signal_4476}), .c ({signal_10626, signal_7139}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7067 ( .a ({signal_10357, signal_7012}), .b ({signal_10419, signal_7038}), .c ({signal_10627, signal_7140}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7068 ( .a ({signal_10358, signal_4463}), .b ({signal_10420, signal_7039}), .c ({signal_10628, signal_7141}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7069 ( .a ({signal_10361, signal_7013}), .b ({signal_10514, signal_7055}), .c ({signal_10783, signal_7142}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7070 ( .a ({signal_10361, signal_7013}), .b ({signal_10423, signal_3952}), .c ({signal_10629, signal_7143}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7071 ( .a ({signal_10250, signal_6963}), .b ({signal_10355, signal_4468}), .c ({signal_10630, signal_7144}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7072 ( .a ({signal_10206, signal_6916}), .b ({signal_10418, signal_4476}), .c ({signal_10631, signal_7145}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7073 ( .a ({signal_10390, signal_4484}), .b ({signal_10419, signal_7038}), .c ({signal_10632, signal_7146}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7074 ( .a ({signal_10301, signal_4460}), .b ({signal_10391, signal_7026}), .c ({signal_10633, signal_7147}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7075 ( .a ({signal_10391, signal_7026}), .b ({signal_10420, signal_7039}), .c ({signal_10634, signal_7148}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7076 ( .a ({signal_10302, signal_6903}), .b ({signal_10392, signal_7027}), .c ({signal_10635, signal_7149}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7077 ( .a ({signal_10392, signal_7027}), .b ({signal_10421, signal_4471}), .c ({signal_10636, signal_7150}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7078 ( .a ({signal_10303, signal_6904}), .b ({signal_10393, signal_4479}), .c ({signal_10637, signal_7151}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7079 ( .a ({signal_10395, signal_3960}), .b ({signal_10424, signal_7040}), .c ({signal_10638, signal_7152}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7080 ( .a ({signal_10306, signal_3936}), .b ({signal_10396, signal_7028}), .c ({signal_10639, signal_7153}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7081 ( .a ({signal_10095, signal_6705}), .b ({signal_10390, signal_4484}), .c ({signal_10640, signal_7154}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7082 ( .a ({signal_10355, signal_4468}), .b ({signal_10359, signal_3943}), .c ({signal_10641, signal_7155}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7083 ( .a ({signal_10355, signal_4468}), .b ({signal_10360, signal_3944}), .c ({signal_10642, signal_7156}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7084 ( .a ({signal_10151, signal_6858}), .b ({signal_10355, signal_4468}), .c ({signal_10643, signal_7157}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7085 ( .a ({signal_10418, signal_4476}), .b ({signal_10422, signal_3951}), .c ({signal_10644, signal_7158}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7086 ( .a ({signal_10418, signal_4476}), .b ({signal_10423, signal_3952}), .c ({signal_10645, signal_7159}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7087 ( .a ({signal_10250, signal_6963}), .b ({signal_10418, signal_4476}), .c ({signal_10646, signal_7160}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7088 ( .a ({signal_10390, signal_4484}), .b ({signal_10394, signal_3959}), .c ({signal_10647, signal_7161}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7089 ( .a ({signal_10390, signal_4484}), .b ({signal_10395, signal_3960}), .c ({signal_10648, signal_7162}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7090 ( .a ({signal_10206, signal_6916}), .b ({signal_10390, signal_4484}), .c ({signal_10649, signal_7163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7091 ( .a ({signal_10363, signal_7014}), .b ({signal_10425, signal_4500}), .c ({signal_10650, signal_7164}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7092 ( .a ({signal_10364, signal_7015}), .b ({signal_10426, signal_7041}), .c ({signal_10651, signal_7165}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7093 ( .a ({signal_10365, signal_4487}), .b ({signal_10427, signal_7042}), .c ({signal_10652, signal_7166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7094 ( .a ({signal_10368, signal_7016}), .b ({signal_10430, signal_3976}), .c ({signal_10653, signal_7167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7095 ( .a ({signal_10397, signal_4508}), .b ({signal_10426, signal_7041}), .c ({signal_10654, signal_7168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7096 ( .a ({signal_10398, signal_7029}), .b ({signal_10427, signal_7042}), .c ({signal_10655, signal_7169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7097 ( .a ({signal_10399, signal_7030}), .b ({signal_10428, signal_4495}), .c ({signal_10656, signal_7170}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7098 ( .a ({signal_10402, signal_3984}), .b ({signal_10431, signal_7043}), .c ({signal_10657, signal_7171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7099 ( .a ({signal_10217, signal_6927}), .b ({signal_10425, signal_4500}), .c ({signal_10658, signal_7172}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7100 ( .a ({signal_10173, signal_6880}), .b ({signal_10397, signal_4508}), .c ({signal_10659, signal_7173}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7101 ( .a ({signal_10369, signal_4516}), .b ({signal_10398, signal_7029}), .c ({signal_10660, signal_7174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7102 ( .a ({signal_10362, signal_4492}), .b ({signal_10370, signal_7017}), .c ({signal_10661, signal_7175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7103 ( .a ({signal_10370, signal_7017}), .b ({signal_10399, signal_7030}), .c ({signal_10662, signal_7176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7104 ( .a ({signal_10363, signal_7014}), .b ({signal_10371, signal_7018}), .c ({signal_10663, signal_7177}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7105 ( .a ({signal_10371, signal_7018}), .b ({signal_10400, signal_4503}), .c ({signal_10664, signal_7178}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7106 ( .a ({signal_10364, signal_7015}), .b ({signal_10372, signal_4511}), .c ({signal_10665, signal_7179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7107 ( .a ({signal_10374, signal_3992}), .b ({signal_10403, signal_7031}), .c ({signal_10666, signal_7180}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7108 ( .a ({signal_10367, signal_3968}), .b ({signal_10375, signal_7019}), .c ({signal_10667, signal_7181}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7109 ( .a ({signal_10261, signal_6974}), .b ({signal_10362, signal_4492}), .c ({signal_10668, signal_7182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7110 ( .a ({signal_10162, signal_6869}), .b ({signal_10369, signal_4516}), .c ({signal_10669, signal_7183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7111 ( .a ({signal_10362, signal_4492}), .b ({signal_10366, signal_3967}), .c ({signal_10670, signal_7184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7112 ( .a ({signal_10362, signal_4492}), .b ({signal_10367, signal_3968}), .c ({signal_10671, signal_7185}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7113 ( .a ({signal_10162, signal_6869}), .b ({signal_10362, signal_4492}), .c ({signal_10672, signal_7186}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7114 ( .a ({signal_10425, signal_4500}), .b ({signal_10429, signal_3975}), .c ({signal_10673, signal_7187}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7115 ( .a ({signal_10425, signal_4500}), .b ({signal_10430, signal_3976}), .c ({signal_10674, signal_7188}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7116 ( .a ({signal_10261, signal_6974}), .b ({signal_10425, signal_4500}), .c ({signal_10675, signal_7189}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7117 ( .a ({signal_10397, signal_4508}), .b ({signal_10401, signal_3983}), .c ({signal_10676, signal_7190}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7118 ( .a ({signal_10397, signal_4508}), .b ({signal_10402, signal_3984}), .c ({signal_10677, signal_7191}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7119 ( .a ({signal_10217, signal_6927}), .b ({signal_10397, signal_4508}), .c ({signal_10678, signal_7192}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7120 ( .a ({signal_10369, signal_4516}), .b ({signal_10373, signal_3991}), .c ({signal_10679, signal_7193}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7121 ( .a ({signal_10369, signal_4516}), .b ({signal_10374, signal_3992}), .c ({signal_10680, signal_7194}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7122 ( .a ({signal_10173, signal_6880}), .b ({signal_10369, signal_4516}), .c ({signal_10681, signal_7195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7123 ( .a ({signal_7775, signal_4305}), .b ({signal_10450, signal_7064}), .c ({signal_10682, signal_7196}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7124 ( .a ({signal_7691, signal_4338}), .b ({signal_10432, signal_7056}), .c ({signal_10683, signal_7197}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7125 ( .a ({signal_7769, signal_4307}), .b ({signal_10451, signal_4147}), .c ({signal_10684, signal_4179}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7126 ( .a ({signal_7766, signal_4308}), .b ({signal_10452, signal_7065}), .c ({signal_10685, signal_7198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7127 ( .a ({signal_7760, signal_4309}), .b ({signal_10453, signal_7066}), .c ({signal_10686, signal_7199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7128 ( .a ({signal_7757, signal_4310}), .b ({signal_10454, signal_4150}), .c ({signal_10687, signal_4182}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7129 ( .a ({signal_7754, signal_4311}), .b ({signal_10433, signal_4151}), .c ({signal_10688, signal_4183}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7130 ( .a ({signal_7751, signal_4312}), .b ({signal_10434, signal_4152}), .c ({signal_10689, signal_4184}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7131 ( .a ({signal_7820, signal_4291}), .b ({signal_10437, signal_4131}), .c ({signal_10690, signal_4163}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7132 ( .a ({signal_7817, signal_4292}), .b ({signal_10438, signal_7059}), .c ({signal_10691, signal_7200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7133 ( .a ({signal_7814, signal_4293}), .b ({signal_10439, signal_7060}), .c ({signal_10692, signal_7201}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7134 ( .a ({signal_7811, signal_4294}), .b ({signal_10440, signal_4134}), .c ({signal_10693, signal_4166}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7135 ( .a ({signal_7748, signal_4313}), .b ({signal_10435, signal_7057}), .c ({signal_10694, signal_7202}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7136 ( .a ({signal_7808, signal_4295}), .b ({signal_10441, signal_4135}), .c ({signal_10695, signal_4167}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7137 ( .a ({signal_7805, signal_4296}), .b ({signal_10442, signal_4136}), .c ({signal_10696, signal_4168}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7138 ( .a ({signal_7802, signal_4297}), .b ({signal_10443, signal_7061}), .c ({signal_10697, signal_7203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7139 ( .a ({signal_7715, signal_4330}), .b ({signal_10436, signal_7058}), .c ({signal_10698, signal_7204}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7140 ( .a ({signal_7793, signal_4299}), .b ({signal_10444, signal_4139}), .c ({signal_10699, signal_4171}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7141 ( .a ({signal_7790, signal_4300}), .b ({signal_10445, signal_7062}), .c ({signal_10700, signal_7205}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7142 ( .a ({signal_7787, signal_4301}), .b ({signal_10446, signal_7063}), .c ({signal_10701, signal_7206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7143 ( .a ({signal_7784, signal_4302}), .b ({signal_10447, signal_4142}), .c ({signal_10702, signal_4174}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7144 ( .a ({signal_7781, signal_4303}), .b ({signal_10448, signal_4143}), .c ({signal_10703, signal_4175}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7145 ( .a ({signal_7778, signal_4304}), .b ({signal_10449, signal_4144}), .c ({signal_10704, signal_4176}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7146 ( .a ({signal_7664, signal_4346}), .b ({signal_10455, signal_7067}), .c ({signal_10705, signal_7207}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7147 ( .a ({signal_10682, signal_7196}), .b ({signal_10784, signal_4177}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7148 ( .a ({signal_10683, signal_7197}), .b ({signal_10785, signal_4210}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7149 ( .a ({signal_10685, signal_7198}), .b ({signal_10786, signal_4180}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7150 ( .a ({signal_10686, signal_7199}), .b ({signal_10787, signal_4181}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7151 ( .a ({signal_10691, signal_7200}), .b ({signal_10788, signal_4164}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7152 ( .a ({signal_10692, signal_7201}), .b ({signal_10789, signal_4165}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7153 ( .a ({signal_10694, signal_7202}), .b ({signal_10790, signal_4185}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7154 ( .a ({signal_10697, signal_7203}), .b ({signal_10791, signal_4169}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7155 ( .a ({signal_10698, signal_7204}), .b ({signal_10792, signal_4202}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7156 ( .a ({signal_10700, signal_7205}), .b ({signal_10793, signal_4172}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7157 ( .a ({signal_10701, signal_7206}), .b ({signal_10794, signal_4173}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7158 ( .a ({signal_10705, signal_7207}), .b ({signal_10795, signal_4218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7159 ( .a ({signal_10228, signal_6938}), .b ({signal_10584, signal_7090}), .c ({signal_10796, signal_7208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7160 ( .a ({signal_10376, signal_4412}), .b ({signal_10577, signal_7083}), .c ({signal_10797, signal_7209}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7161 ( .a ({signal_10377, signal_7020}), .b ({signal_10579, signal_7085}), .c ({signal_10798, signal_7210}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7162 ( .a ({signal_10378, signal_7021}), .b ({signal_10581, signal_7087}), .c ({signal_10799, signal_7211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7163 ( .a ({signal_10341, signal_4420}), .b ({signal_10570, signal_7075}), .c ({signal_10800, signal_7212}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7164 ( .a ({signal_10342, signal_7005}), .b ({signal_10571, signal_7076}), .c ({signal_10801, signal_7213}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7165 ( .a ({signal_10381, signal_3888}), .b ({signal_10583, signal_7089}), .c ({signal_10802, signal_7214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7166 ( .a ({signal_10343, signal_7006}), .b ({signal_10572, signal_7077}), .c ({signal_10803, signal_7215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7167 ( .a ({signal_10346, signal_3896}), .b ({signal_10573, signal_7079}), .c ({signal_10804, signal_7216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7168 ( .a ({signal_10774, signal_7074}), .b ({signal_10574, signal_7080}), .c ({signal_11008, signal_7217}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7169 ( .a ({signal_10315, signal_4396}), .b ({signal_10576, signal_7082}), .c ({signal_10805, signal_7218}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7170 ( .a ({signal_10316, signal_6975}), .b ({signal_10578, signal_7084}), .c ({signal_10806, signal_7219}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7171 ( .a ({signal_10317, signal_6976}), .b ({signal_10580, signal_7086}), .c ({signal_10807, signal_7220}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7172 ( .a ({signal_10379, signal_4407}), .b ({signal_10585, signal_7091}), .c ({signal_10808, signal_7221}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7173 ( .a ({signal_10321, signal_6977}), .b ({signal_10593, signal_7099}), .c ({signal_10809, signal_7222}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7174 ( .a ({signal_10380, signal_3887}), .b ({signal_10586, signal_7092}), .c ({signal_10810, signal_7223}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7175 ( .a ({signal_10320, signal_3872}), .b ({signal_10582, signal_7088}), .c ({signal_10811, signal_7224}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7176 ( .a ({signal_10382, signal_7022}), .b ({signal_10587, signal_7093}), .c ({signal_10812, signal_7225}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7177 ( .a ({signal_10347, signal_7007}), .b ({signal_10590, signal_7096}), .c ({signal_10813, signal_7226}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7178 ( .a ({signal_10117, signal_6781}), .b ({signal_10575, signal_7081}), .c ({signal_10814, signal_7227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7179 ( .a ({signal_10404, signal_4404}), .b ({signal_10577, signal_7083}), .c ({signal_10815, signal_7228}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7180 ( .a ({signal_10405, signal_7032}), .b ({signal_10579, signal_7085}), .c ({signal_10816, signal_7229}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7181 ( .a ({signal_10406, signal_7033}), .b ({signal_10581, signal_7087}), .c ({signal_10817, signal_7230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7182 ( .a ({signal_10344, signal_4415}), .b ({signal_10588, signal_7094}), .c ({signal_10818, signal_7231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7183 ( .a ({signal_10318, signal_4391}), .b ({signal_10591, signal_7097}), .c ({signal_10819, signal_7232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7184 ( .a ({signal_10345, signal_3895}), .b ({signal_10589, signal_7095}), .c ({signal_10820, signal_7233}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7185 ( .a ({signal_10319, signal_3871}), .b ({signal_10592, signal_7098}), .c ({signal_10821, signal_7234}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7186 ( .a ({signal_10409, signal_3880}), .b ({signal_10583, signal_7089}), .c ({signal_10822, signal_7235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7187 ( .a ({signal_10503, signal_7044}), .b ({signal_10584, signal_7090}), .c ({signal_10823, signal_7236}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7188 ( .a ({signal_10195, signal_6902}), .b ({signal_10612, signal_7122}), .c ({signal_10824, signal_7237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7189 ( .a ({signal_10348, signal_4444}), .b ({signal_10605, signal_7115}), .c ({signal_10825, signal_7238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7190 ( .a ({signal_10349, signal_7008}), .b ({signal_10607, signal_7117}), .c ({signal_10826, signal_7239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7191 ( .a ({signal_10350, signal_7009}), .b ({signal_10609, signal_7119}), .c ({signal_10827, signal_7240}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7192 ( .a ({signal_10411, signal_4452}), .b ({signal_10598, signal_7107}), .c ({signal_10828, signal_7241}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7193 ( .a ({signal_10412, signal_7035}), .b ({signal_10599, signal_7108}), .c ({signal_10829, signal_7242}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7194 ( .a ({signal_10353, signal_3920}), .b ({signal_10611, signal_7121}), .c ({signal_10830, signal_7243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7195 ( .a ({signal_10413, signal_7036}), .b ({signal_10600, signal_7109}), .c ({signal_10831, signal_7244}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7196 ( .a ({signal_10416, signal_3928}), .b ({signal_10601, signal_7111}), .c ({signal_10832, signal_7245}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7197 ( .a ({signal_10778, signal_7106}), .b ({signal_10602, signal_7112}), .c ({signal_11009, signal_7246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7198 ( .a ({signal_10308, signal_4428}), .b ({signal_10604, signal_7114}), .c ({signal_10833, signal_7247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7199 ( .a ({signal_10309, signal_6939}), .b ({signal_10606, signal_7116}), .c ({signal_10834, signal_7248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7200 ( .a ({signal_10310, signal_6940}), .b ({signal_10608, signal_7118}), .c ({signal_10835, signal_7249}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7201 ( .a ({signal_10351, signal_4439}), .b ({signal_10613, signal_7123}), .c ({signal_10836, signal_7250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7202 ( .a ({signal_10314, signal_6941}), .b ({signal_10621, signal_7131}), .c ({signal_10837, signal_7251}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7203 ( .a ({signal_10352, signal_3919}), .b ({signal_10614, signal_7124}), .c ({signal_10838, signal_7252}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7204 ( .a ({signal_10313, signal_3904}), .b ({signal_10610, signal_7120}), .c ({signal_10839, signal_7253}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7205 ( .a ({signal_10354, signal_7010}), .b ({signal_10615, signal_7125}), .c ({signal_10840, signal_7254}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7206 ( .a ({signal_10417, signal_7037}), .b ({signal_10618, signal_7128}), .c ({signal_10841, signal_7255}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7207 ( .a ({signal_10106, signal_6743}), .b ({signal_10603, signal_7113}), .c ({signal_10842, signal_7256}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7208 ( .a ({signal_10383, signal_4436}), .b ({signal_10605, signal_7115}), .c ({signal_10843, signal_7257}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7209 ( .a ({signal_10384, signal_7023}), .b ({signal_10607, signal_7117}), .c ({signal_10844, signal_7258}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7210 ( .a ({signal_10385, signal_7024}), .b ({signal_10609, signal_7119}), .c ({signal_10845, signal_7259}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7211 ( .a ({signal_10414, signal_4447}), .b ({signal_10616, signal_7126}), .c ({signal_10846, signal_7260}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7212 ( .a ({signal_10311, signal_4423}), .b ({signal_10619, signal_7129}), .c ({signal_10847, signal_7261}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7213 ( .a ({signal_10415, signal_3927}), .b ({signal_10617, signal_7127}), .c ({signal_10848, signal_7262}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7214 ( .a ({signal_10312, signal_3903}), .b ({signal_10620, signal_7130}), .c ({signal_10849, signal_7263}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7215 ( .a ({signal_10388, signal_3912}), .b ({signal_10611, signal_7121}), .c ({signal_10850, signal_7264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7216 ( .a ({signal_10507, signal_7048}), .b ({signal_10612, signal_7122}), .c ({signal_10851, signal_7265}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7217 ( .a ({signal_10151, signal_6858}), .b ({signal_10640, signal_7154}), .c ({signal_10852, signal_7266}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7218 ( .a ({signal_10418, signal_4476}), .b ({signal_10633, signal_7147}), .c ({signal_10853, signal_7267}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7219 ( .a ({signal_10419, signal_7038}), .b ({signal_10635, signal_7149}), .c ({signal_10854, signal_7268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7220 ( .a ({signal_10420, signal_7039}), .b ({signal_10637, signal_7151}), .c ({signal_10855, signal_7269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7221 ( .a ({signal_10390, signal_4484}), .b ({signal_10626, signal_7139}), .c ({signal_10856, signal_7270}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7222 ( .a ({signal_10391, signal_7026}), .b ({signal_10627, signal_7140}), .c ({signal_10857, signal_7271}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7223 ( .a ({signal_10423, signal_3952}), .b ({signal_10639, signal_7153}), .c ({signal_10858, signal_7272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7224 ( .a ({signal_10392, signal_7027}), .b ({signal_10628, signal_7141}), .c ({signal_10859, signal_7273}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7225 ( .a ({signal_10395, signal_3960}), .b ({signal_10629, signal_7143}), .c ({signal_10860, signal_7274}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7226 ( .a ({signal_10782, signal_7138}), .b ({signal_10630, signal_7144}), .c ({signal_11010, signal_7275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7227 ( .a ({signal_10301, signal_4460}), .b ({signal_10632, signal_7146}), .c ({signal_10861, signal_7276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7228 ( .a ({signal_10302, signal_6903}), .b ({signal_10634, signal_7148}), .c ({signal_10862, signal_7277}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7229 ( .a ({signal_10303, signal_6904}), .b ({signal_10636, signal_7150}), .c ({signal_10863, signal_7278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7230 ( .a ({signal_10421, signal_4471}), .b ({signal_10641, signal_7155}), .c ({signal_10864, signal_7279}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7231 ( .a ({signal_10307, signal_6905}), .b ({signal_10649, signal_7163}), .c ({signal_10865, signal_7280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7232 ( .a ({signal_10422, signal_3951}), .b ({signal_10642, signal_7156}), .c ({signal_10866, signal_7281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7233 ( .a ({signal_10306, signal_3936}), .b ({signal_10638, signal_7152}), .c ({signal_10867, signal_7282}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7234 ( .a ({signal_10424, signal_7040}), .b ({signal_10643, signal_7157}), .c ({signal_10868, signal_7283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7235 ( .a ({signal_10396, signal_7028}), .b ({signal_10646, signal_7160}), .c ({signal_10869, signal_7284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7236 ( .a ({signal_10095, signal_6705}), .b ({signal_10631, signal_7145}), .c ({signal_10870, signal_7285}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7237 ( .a ({signal_10355, signal_4468}), .b ({signal_10633, signal_7147}), .c ({signal_10871, signal_7286}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7238 ( .a ({signal_10356, signal_7011}), .b ({signal_10635, signal_7149}), .c ({signal_10872, signal_7287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7239 ( .a ({signal_10357, signal_7012}), .b ({signal_10637, signal_7151}), .c ({signal_10873, signal_7288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7240 ( .a ({signal_10393, signal_4479}), .b ({signal_10644, signal_7158}), .c ({signal_10874, signal_7289}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7241 ( .a ({signal_10304, signal_4455}), .b ({signal_10647, signal_7161}), .c ({signal_10875, signal_7290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7242 ( .a ({signal_10394, signal_3959}), .b ({signal_10645, signal_7159}), .c ({signal_10876, signal_7291}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7243 ( .a ({signal_10305, signal_3935}), .b ({signal_10648, signal_7162}), .c ({signal_10877, signal_7292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7244 ( .a ({signal_10360, signal_3944}), .b ({signal_10639, signal_7153}), .c ({signal_10878, signal_7293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7245 ( .a ({signal_10511, signal_7052}), .b ({signal_10640, signal_7154}), .c ({signal_10879, signal_7294}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7246 ( .a ({signal_10261, signal_6974}), .b ({signal_10669, signal_7183}), .c ({signal_10880, signal_7295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7247 ( .a ({signal_10397, signal_4508}), .b ({signal_10661, signal_7175}), .c ({signal_10881, signal_7296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7248 ( .a ({signal_10398, signal_7029}), .b ({signal_10663, signal_7177}), .c ({signal_10882, signal_7297}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7249 ( .a ({signal_10399, signal_7030}), .b ({signal_10665, signal_7179}), .c ({signal_10883, signal_7298}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7250 ( .a ({signal_10369, signal_4516}), .b ({signal_10654, signal_7168}), .c ({signal_10884, signal_7299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7251 ( .a ({signal_10370, signal_7017}), .b ({signal_10655, signal_7169}), .c ({signal_10885, signal_7300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7252 ( .a ({signal_10402, signal_3984}), .b ({signal_10667, signal_7181}), .c ({signal_10886, signal_7301}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7253 ( .a ({signal_10371, signal_7018}), .b ({signal_10656, signal_7170}), .c ({signal_10887, signal_7302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7254 ( .a ({signal_10428, signal_4495}), .b ({signal_10670, signal_7184}), .c ({signal_10888, signal_7303}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7255 ( .a ({signal_10429, signal_3975}), .b ({signal_10671, signal_7185}), .c ({signal_10889, signal_7304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7256 ( .a ({signal_10374, signal_3992}), .b ({signal_10657, signal_7171}), .c ({signal_10890, signal_7305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7257 ( .a ({signal_10173, signal_6880}), .b ({signal_10668, signal_7182}), .c ({signal_10891, signal_7306}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7258 ( .a ({signal_10362, signal_4492}), .b ({signal_10660, signal_7174}), .c ({signal_10892, signal_7307}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7259 ( .a ({signal_10363, signal_7014}), .b ({signal_10662, signal_7176}), .c ({signal_10893, signal_7308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7260 ( .a ({signal_10364, signal_7015}), .b ({signal_10664, signal_7178}), .c ({signal_10894, signal_7309}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7261 ( .a ({signal_10400, signal_4503}), .b ({signal_10673, signal_7187}), .c ({signal_10895, signal_7310}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7262 ( .a ({signal_10431, signal_7043}), .b ({signal_10672, signal_7186}), .c ({signal_10896, signal_7311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7263 ( .a ({signal_10368, signal_7016}), .b ({signal_10681, signal_7195}), .c ({signal_10897, signal_7312}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7264 ( .a ({signal_10401, signal_3983}), .b ({signal_10674, signal_7188}), .c ({signal_10898, signal_7313}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7265 ( .a ({signal_10367, signal_3968}), .b ({signal_10666, signal_7180}), .c ({signal_10899, signal_7314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7266 ( .a ({signal_10403, signal_7031}), .b ({signal_10675, signal_7189}), .c ({signal_10900, signal_7315}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7267 ( .a ({signal_10375, signal_7019}), .b ({signal_10678, signal_7192}), .c ({signal_10901, signal_7316}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7268 ( .a ({signal_10162, signal_6869}), .b ({signal_10659, signal_7173}), .c ({signal_10902, signal_7317}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7269 ( .a ({signal_10425, signal_4500}), .b ({signal_10661, signal_7175}), .c ({signal_10903, signal_7318}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7270 ( .a ({signal_10426, signal_7041}), .b ({signal_10663, signal_7177}), .c ({signal_10904, signal_7319}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7271 ( .a ({signal_10427, signal_7042}), .b ({signal_10665, signal_7179}), .c ({signal_10905, signal_7320}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7272 ( .a ({signal_10372, signal_4511}), .b ({signal_10676, signal_7190}), .c ({signal_10906, signal_7321}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7273 ( .a ({signal_10365, signal_4487}), .b ({signal_10679, signal_7193}), .c ({signal_10907, signal_7322}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7274 ( .a ({signal_10373, signal_3991}), .b ({signal_10677, signal_7191}), .c ({signal_10908, signal_7323}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7275 ( .a ({signal_10366, signal_3967}), .b ({signal_10680, signal_7194}), .c ({signal_10909, signal_7324}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7276 ( .a ({signal_10430, signal_3976}), .b ({signal_10667, signal_7181}), .c ({signal_10910, signal_7325}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7277 ( .a ({signal_10668, signal_7182}), .b ({signal_10669, signal_7183}), .c ({signal_10911, signal_7326}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7278 ( .a ({signal_7823, signal_4370}), .b ({signal_10683, signal_7197}), .c ({signal_10912, signal_7327}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7279 ( .a ({signal_7694, signal_4337}), .b ({signal_10682, signal_7196}), .c ({signal_10913, signal_7328}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7280 ( .a ({signal_7685, signal_4339}), .b ({signal_10684, signal_4179}), .c ({signal_10914, signal_4211}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7281 ( .a ({signal_7682, signal_4340}), .b ({signal_10685, signal_7198}), .c ({signal_10915, signal_7329}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7282 ( .a ({signal_7679, signal_4341}), .b ({signal_10686, signal_7199}), .c ({signal_10916, signal_7330}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7283 ( .a ({signal_7676, signal_4342}), .b ({signal_10687, signal_4182}), .c ({signal_10917, signal_4214}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7284 ( .a ({signal_7673, signal_4343}), .b ({signal_10688, signal_4183}), .c ({signal_10918, signal_4215}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7285 ( .a ({signal_7670, signal_4344}), .b ({signal_10689, signal_4184}), .c ({signal_10919, signal_4216}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7286 ( .a ({signal_7739, signal_4323}), .b ({signal_10690, signal_4163}), .c ({signal_10920, signal_4195}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7287 ( .a ({signal_7736, signal_4324}), .b ({signal_10691, signal_7200}), .c ({signal_10921, signal_7331}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7288 ( .a ({signal_7733, signal_4325}), .b ({signal_10692, signal_7201}), .c ({signal_10922, signal_7332}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7289 ( .a ({signal_7730, signal_4326}), .b ({signal_10693, signal_4166}), .c ({signal_10923, signal_4198}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7290 ( .a ({signal_7667, signal_4345}), .b ({signal_10694, signal_7202}), .c ({signal_10924, signal_7333}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7291 ( .a ({signal_7727, signal_4327}), .b ({signal_10695, signal_4167}), .c ({signal_10925, signal_4199}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7292 ( .a ({signal_7724, signal_4328}), .b ({signal_10696, signal_4168}), .c ({signal_10926, signal_4200}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7293 ( .a ({signal_7718, signal_4329}), .b ({signal_10697, signal_7203}), .c ({signal_10927, signal_7334}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7294 ( .a ({signal_7610, signal_4362}), .b ({signal_10698, signal_7204}), .c ({signal_10928, signal_7335}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7295 ( .a ({signal_7712, signal_4331}), .b ({signal_10699, signal_4171}), .c ({signal_10929, signal_4203}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7296 ( .a ({signal_7709, signal_4332}), .b ({signal_10700, signal_7205}), .c ({signal_10930, signal_7336}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7297 ( .a ({signal_7706, signal_4333}), .b ({signal_10701, signal_7206}), .c ({signal_10931, signal_7337}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7298 ( .a ({signal_7703, signal_4334}), .b ({signal_10702, signal_4174}), .c ({signal_10932, signal_4206}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7299 ( .a ({signal_7700, signal_4335}), .b ({signal_10703, signal_4175}), .c ({signal_10933, signal_4207}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7300 ( .a ({signal_7697, signal_4336}), .b ({signal_10704, signal_4176}), .c ({signal_10934, signal_4208}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7301 ( .a ({signal_7529, signal_4378}), .b ({signal_10705, signal_7207}), .c ({signal_10935, signal_7338}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7302 ( .a ({signal_11008, signal_7217}), .b ({signal_11273, signal_4002}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7303 ( .a ({signal_11009, signal_7246}), .b ({signal_11274, signal_4034}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7304 ( .a ({signal_11010, signal_7275}), .b ({signal_11275, signal_4066}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7305 ( .a ({signal_10912, signal_7327}), .b ({signal_11011, signal_4242}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7306 ( .a ({signal_10913, signal_7328}), .b ({signal_11012, signal_4209}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7307 ( .a ({signal_10915, signal_7329}), .b ({signal_11013, signal_4212}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7308 ( .a ({signal_10916, signal_7330}), .b ({signal_11014, signal_4213}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7309 ( .a ({signal_10921, signal_7331}), .b ({signal_11015, signal_4196}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7310 ( .a ({signal_10922, signal_7332}), .b ({signal_11016, signal_4197}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7311 ( .a ({signal_10924, signal_7333}), .b ({signal_11017, signal_4217}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7312 ( .a ({signal_10927, signal_7334}), .b ({signal_11018, signal_4201}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7313 ( .a ({signal_10928, signal_7335}), .b ({signal_11019, signal_4234}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7314 ( .a ({signal_10930, signal_7336}), .b ({signal_11020, signal_4204}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7315 ( .a ({signal_10931, signal_7337}), .b ({signal_11021, signal_4205}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7316 ( .a ({signal_10935, signal_7338}), .b ({signal_11022, signal_4250}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7317 ( .a ({signal_10809, signal_7222}), .b ({signal_10813, signal_7226}), .c ({signal_11023, signal_7339}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7318 ( .a ({signal_10575, signal_7081}), .b ({signal_10796, signal_7208}), .c ({signal_11024, signal_7340}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7319 ( .a ({signal_10566, signal_7068}), .b ({signal_10797, signal_7209}), .c ({signal_11025, signal_4019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7320 ( .a ({signal_10567, signal_7069}), .b ({signal_10798, signal_7210}), .c ({signal_11026, signal_7341}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7321 ( .a ({signal_10568, signal_7070}), .b ({signal_10799, signal_7211}), .c ({signal_11027, signal_7342}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7322 ( .a ({signal_10379, signal_4407}), .b ({signal_10819, signal_7232}), .c ({signal_11028, signal_7343}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7323 ( .a ({signal_10380, signal_3887}), .b ({signal_10821, signal_7234}), .c ({signal_11029, signal_7344}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7324 ( .a ({signal_10566, signal_7068}), .b ({signal_10800, signal_7212}), .c ({signal_11030, signal_3995}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7325 ( .a ({signal_10567, signal_7069}), .b ({signal_10801, signal_7213}), .c ({signal_11031, signal_7345}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7326 ( .a ({signal_10569, signal_7073}), .b ({signal_10802, signal_7214}), .c ({signal_11032, signal_4024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7327 ( .a ({signal_10568, signal_7070}), .b ({signal_10803, signal_7215}), .c ({signal_11033, signal_7346}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7328 ( .a ({signal_10344, signal_4415}), .b ({signal_10808, signal_7221}), .c ({signal_11034, signal_7347}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7329 ( .a ({signal_10345, signal_3895}), .b ({signal_10810, signal_7223}), .c ({signal_11035, signal_7348}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7330 ( .a ({signal_10569, signal_7073}), .b ({signal_10804, signal_7216}), .c ({signal_11036, signal_4000}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7331 ( .a ({signal_10347, signal_7007}), .b ({signal_10812, signal_7225}), .c ({signal_11037, signal_7349}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7332 ( .a ({signal_10570, signal_7075}), .b ({signal_10805, signal_7218}), .c ({signal_11038, signal_4003}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7333 ( .a ({signal_10571, signal_7076}), .b ({signal_10806, signal_7219}), .c ({signal_11039, signal_7350}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7334 ( .a ({signal_10572, signal_7077}), .b ({signal_10807, signal_7220}), .c ({signal_11040, signal_7351}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7335 ( .a ({signal_10318, signal_4391}), .b ({signal_10818, signal_7231}), .c ({signal_11041, signal_7352}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7336 ( .a ({signal_10382, signal_7022}), .b ({signal_10809, signal_7222}), .c ({signal_11042, signal_7353}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7337 ( .a ({signal_10319, signal_3871}), .b ({signal_10820, signal_7233}), .c ({signal_11043, signal_7354}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7338 ( .a ({signal_10573, signal_7079}), .b ({signal_10811, signal_7224}), .c ({signal_11044, signal_4008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7339 ( .a ({signal_10321, signal_6977}), .b ({signal_10813, signal_7226}), .c ({signal_11045, signal_7355}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7340 ( .a ({signal_10574, signal_7080}), .b ({signal_10814, signal_7227}), .c ({signal_11046, signal_7356}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7341 ( .a ({signal_10576, signal_7082}), .b ({signal_10815, signal_7228}), .c ({signal_11047, signal_4011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7342 ( .a ({signal_10578, signal_7084}), .b ({signal_10816, signal_7229}), .c ({signal_11048, signal_7357}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7343 ( .a ({signal_10580, signal_7086}), .b ({signal_10817, signal_7230}), .c ({signal_11049, signal_7358}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7344 ( .a ({signal_10407, signal_4399}), .b ({signal_10819, signal_7232}), .c ({signal_11050, signal_7359}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7345 ( .a ({signal_10408, signal_3879}), .b ({signal_10821, signal_7234}), .c ({signal_11051, signal_7360}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7346 ( .a ({signal_10582, signal_7088}), .b ({signal_10822, signal_7235}), .c ({signal_11052, signal_4016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7347 ( .a ({signal_10184, signal_6891}), .b ({signal_10823, signal_7236}), .c ({signal_11053, signal_7361}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7348 ( .a ({signal_10837, signal_7251}), .b ({signal_10841, signal_7255}), .c ({signal_11054, signal_7362}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7349 ( .a ({signal_10603, signal_7113}), .b ({signal_10824, signal_7237}), .c ({signal_11055, signal_7363}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7350 ( .a ({signal_10594, signal_7100}), .b ({signal_10825, signal_7238}), .c ({signal_11056, signal_4051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7351 ( .a ({signal_10595, signal_7101}), .b ({signal_10826, signal_7239}), .c ({signal_11057, signal_7364}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7352 ( .a ({signal_10596, signal_7102}), .b ({signal_10827, signal_7240}), .c ({signal_11058, signal_7365}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7353 ( .a ({signal_10351, signal_4439}), .b ({signal_10847, signal_7261}), .c ({signal_11059, signal_7366}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7354 ( .a ({signal_10352, signal_3919}), .b ({signal_10849, signal_7263}), .c ({signal_11060, signal_7367}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7355 ( .a ({signal_10594, signal_7100}), .b ({signal_10828, signal_7241}), .c ({signal_11061, signal_4027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7356 ( .a ({signal_10595, signal_7101}), .b ({signal_10829, signal_7242}), .c ({signal_11062, signal_7368}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7357 ( .a ({signal_10597, signal_7105}), .b ({signal_10830, signal_7243}), .c ({signal_11063, signal_4056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7358 ( .a ({signal_10596, signal_7102}), .b ({signal_10831, signal_7244}), .c ({signal_11064, signal_7369}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7359 ( .a ({signal_10414, signal_4447}), .b ({signal_10836, signal_7250}), .c ({signal_11065, signal_7370}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7360 ( .a ({signal_10415, signal_3927}), .b ({signal_10838, signal_7252}), .c ({signal_11066, signal_7371}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7361 ( .a ({signal_10597, signal_7105}), .b ({signal_10832, signal_7245}), .c ({signal_11067, signal_4032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7362 ( .a ({signal_10417, signal_7037}), .b ({signal_10840, signal_7254}), .c ({signal_11068, signal_7372}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7363 ( .a ({signal_10598, signal_7107}), .b ({signal_10833, signal_7247}), .c ({signal_11069, signal_4035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7364 ( .a ({signal_10599, signal_7108}), .b ({signal_10834, signal_7248}), .c ({signal_11070, signal_7373}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7365 ( .a ({signal_10600, signal_7109}), .b ({signal_10835, signal_7249}), .c ({signal_11071, signal_7374}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7366 ( .a ({signal_10311, signal_4423}), .b ({signal_10846, signal_7260}), .c ({signal_11072, signal_7375}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7367 ( .a ({signal_10354, signal_7010}), .b ({signal_10837, signal_7251}), .c ({signal_11073, signal_7376}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7368 ( .a ({signal_10312, signal_3903}), .b ({signal_10848, signal_7262}), .c ({signal_11074, signal_7377}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7369 ( .a ({signal_10601, signal_7111}), .b ({signal_10839, signal_7253}), .c ({signal_11075, signal_4040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7370 ( .a ({signal_10314, signal_6941}), .b ({signal_10841, signal_7255}), .c ({signal_11076, signal_7378}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7371 ( .a ({signal_10602, signal_7112}), .b ({signal_10842, signal_7256}), .c ({signal_11077, signal_7379}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7372 ( .a ({signal_10604, signal_7114}), .b ({signal_10843, signal_7257}), .c ({signal_11078, signal_4043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7373 ( .a ({signal_10606, signal_7116}), .b ({signal_10844, signal_7258}), .c ({signal_11079, signal_7380}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7374 ( .a ({signal_10608, signal_7118}), .b ({signal_10845, signal_7259}), .c ({signal_11080, signal_7381}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7375 ( .a ({signal_10386, signal_4431}), .b ({signal_10847, signal_7261}), .c ({signal_11081, signal_7382}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7376 ( .a ({signal_10387, signal_3911}), .b ({signal_10849, signal_7263}), .c ({signal_11082, signal_7383}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7377 ( .a ({signal_10610, signal_7120}), .b ({signal_10850, signal_7264}), .c ({signal_11083, signal_4048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7378 ( .a ({signal_10140, signal_6847}), .b ({signal_10851, signal_7265}), .c ({signal_11084, signal_7384}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7379 ( .a ({signal_10865, signal_7280}), .b ({signal_10869, signal_7284}), .c ({signal_11085, signal_7385}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7380 ( .a ({signal_10631, signal_7145}), .b ({signal_10852, signal_7266}), .c ({signal_11086, signal_7386}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7381 ( .a ({signal_10622, signal_7132}), .b ({signal_10853, signal_7267}), .c ({signal_11087, signal_4083}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7382 ( .a ({signal_10623, signal_7133}), .b ({signal_10854, signal_7268}), .c ({signal_11088, signal_7387}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7383 ( .a ({signal_10624, signal_7134}), .b ({signal_10855, signal_7269}), .c ({signal_11089, signal_7388}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7384 ( .a ({signal_10421, signal_4471}), .b ({signal_10875, signal_7290}), .c ({signal_11090, signal_7389}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7385 ( .a ({signal_10422, signal_3951}), .b ({signal_10877, signal_7292}), .c ({signal_11091, signal_7390}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7386 ( .a ({signal_10622, signal_7132}), .b ({signal_10856, signal_7270}), .c ({signal_11092, signal_4059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7387 ( .a ({signal_10623, signal_7133}), .b ({signal_10857, signal_7271}), .c ({signal_11093, signal_7391}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7388 ( .a ({signal_10625, signal_7137}), .b ({signal_10858, signal_7272}), .c ({signal_11094, signal_4088}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7389 ( .a ({signal_10624, signal_7134}), .b ({signal_10859, signal_7273}), .c ({signal_11095, signal_7392}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7390 ( .a ({signal_10393, signal_4479}), .b ({signal_10864, signal_7279}), .c ({signal_11096, signal_7393}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7391 ( .a ({signal_10394, signal_3959}), .b ({signal_10866, signal_7281}), .c ({signal_11097, signal_7394}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7392 ( .a ({signal_10625, signal_7137}), .b ({signal_10860, signal_7274}), .c ({signal_11098, signal_4064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7393 ( .a ({signal_10396, signal_7028}), .b ({signal_10868, signal_7283}), .c ({signal_11099, signal_7395}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7394 ( .a ({signal_10626, signal_7139}), .b ({signal_10861, signal_7276}), .c ({signal_11100, signal_4067}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7395 ( .a ({signal_10627, signal_7140}), .b ({signal_10862, signal_7277}), .c ({signal_11101, signal_7396}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7396 ( .a ({signal_10628, signal_7141}), .b ({signal_10863, signal_7278}), .c ({signal_11102, signal_7397}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7397 ( .a ({signal_10304, signal_4455}), .b ({signal_10874, signal_7289}), .c ({signal_11103, signal_7398}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7398 ( .a ({signal_10424, signal_7040}), .b ({signal_10865, signal_7280}), .c ({signal_11104, signal_7399}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7399 ( .a ({signal_10305, signal_3935}), .b ({signal_10876, signal_7291}), .c ({signal_11105, signal_7400}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7400 ( .a ({signal_10629, signal_7143}), .b ({signal_10867, signal_7282}), .c ({signal_11106, signal_4072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7401 ( .a ({signal_10307, signal_6905}), .b ({signal_10869, signal_7284}), .c ({signal_11107, signal_7401}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7402 ( .a ({signal_10630, signal_7144}), .b ({signal_10870, signal_7285}), .c ({signal_11108, signal_7402}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7403 ( .a ({signal_10632, signal_7146}), .b ({signal_10871, signal_7286}), .c ({signal_11109, signal_4075}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7404 ( .a ({signal_10634, signal_7148}), .b ({signal_10872, signal_7287}), .c ({signal_11110, signal_7403}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7405 ( .a ({signal_10636, signal_7150}), .b ({signal_10873, signal_7288}), .c ({signal_11111, signal_7404}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7406 ( .a ({signal_10358, signal_4463}), .b ({signal_10875, signal_7290}), .c ({signal_11112, signal_7405}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7407 ( .a ({signal_10359, signal_3943}), .b ({signal_10877, signal_7292}), .c ({signal_11113, signal_7406}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7408 ( .a ({signal_10638, signal_7152}), .b ({signal_10878, signal_7293}), .c ({signal_11114, signal_4080}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7409 ( .a ({signal_10250, signal_6963}), .b ({signal_10879, signal_7294}), .c ({signal_11115, signal_7407}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7410 ( .a ({signal_10897, signal_7312}), .b ({signal_10901, signal_7316}), .c ({signal_11116, signal_7408}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7411 ( .a ({signal_10659, signal_7173}), .b ({signal_10880, signal_7295}), .c ({signal_11117, signal_7409}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7412 ( .a ({signal_10650, signal_7164}), .b ({signal_10881, signal_7296}), .c ({signal_11118, signal_4115}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7413 ( .a ({signal_10651, signal_7165}), .b ({signal_10882, signal_7297}), .c ({signal_11119, signal_7410}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7414 ( .a ({signal_10652, signal_7166}), .b ({signal_10883, signal_7298}), .c ({signal_11120, signal_7411}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7415 ( .a ({signal_10400, signal_4503}), .b ({signal_10907, signal_7322}), .c ({signal_11121, signal_7412}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7416 ( .a ({signal_10401, signal_3983}), .b ({signal_10909, signal_7324}), .c ({signal_11122, signal_7413}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7417 ( .a ({signal_10650, signal_7164}), .b ({signal_10884, signal_7299}), .c ({signal_11123, signal_4091}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7418 ( .a ({signal_10651, signal_7165}), .b ({signal_10885, signal_7300}), .c ({signal_11124, signal_7414}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7419 ( .a ({signal_10653, signal_7167}), .b ({signal_10886, signal_7301}), .c ({signal_11125, signal_4120}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7420 ( .a ({signal_10652, signal_7166}), .b ({signal_10887, signal_7302}), .c ({signal_11126, signal_7415}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7421 ( .a ({signal_10372, signal_4511}), .b ({signal_10895, signal_7310}), .c ({signal_11127, signal_7416}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7422 ( .a ({signal_10373, signal_3991}), .b ({signal_10898, signal_7313}), .c ({signal_11128, signal_7417}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7423 ( .a ({signal_10653, signal_7167}), .b ({signal_10890, signal_7305}), .c ({signal_11129, signal_4096}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7424 ( .a ({signal_10375, signal_7019}), .b ({signal_10900, signal_7315}), .c ({signal_11130, signal_7418}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7425 ( .a ({signal_10658, signal_7172}), .b ({signal_10891, signal_7306}), .c ({signal_11131, signal_7419}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7426 ( .a ({signal_10654, signal_7168}), .b ({signal_10892, signal_7307}), .c ({signal_11132, signal_4099}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7427 ( .a ({signal_10655, signal_7169}), .b ({signal_10893, signal_7308}), .c ({signal_11133, signal_7420}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7428 ( .a ({signal_10656, signal_7170}), .b ({signal_10894, signal_7309}), .c ({signal_11134, signal_7421}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7429 ( .a ({signal_10365, signal_4487}), .b ({signal_10906, signal_7321}), .c ({signal_11135, signal_7422}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7430 ( .a ({signal_10403, signal_7031}), .b ({signal_10897, signal_7312}), .c ({signal_11136, signal_7423}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7431 ( .a ({signal_10366, signal_3967}), .b ({signal_10908, signal_7323}), .c ({signal_11137, signal_7424}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7432 ( .a ({signal_10657, signal_7171}), .b ({signal_10899, signal_7314}), .c ({signal_11138, signal_4104}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7433 ( .a ({signal_10368, signal_7016}), .b ({signal_10901, signal_7316}), .c ({signal_11139, signal_7425}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7434 ( .a ({signal_10658, signal_7172}), .b ({signal_10902, signal_7317}), .c ({signal_11140, signal_7426}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7435 ( .a ({signal_10660, signal_7174}), .b ({signal_10903, signal_7318}), .c ({signal_11141, signal_4107}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7436 ( .a ({signal_10662, signal_7176}), .b ({signal_10904, signal_7319}), .c ({signal_11142, signal_7427}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7437 ( .a ({signal_10664, signal_7178}), .b ({signal_10905, signal_7320}), .c ({signal_11143, signal_7428}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7438 ( .a ({signal_10428, signal_4495}), .b ({signal_10907, signal_7322}), .c ({signal_11144, signal_7429}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7439 ( .a ({signal_10429, signal_3975}), .b ({signal_10909, signal_7324}), .c ({signal_11145, signal_7430}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7440 ( .a ({signal_10666, signal_7180}), .b ({signal_10910, signal_7325}), .c ({signal_11146, signal_4112}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7441 ( .a ({signal_10217, signal_6927}), .b ({signal_10911, signal_7326}), .c ({signal_11147, signal_7431}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7442 ( .a ({signal_7838, signal_4369}), .b ({signal_10913, signal_7328}), .c ({signal_11148, signal_7432}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7443 ( .a ({signal_7796, signal_4371}), .b ({signal_10914, signal_4211}), .c ({signal_11149, signal_4243}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7444 ( .a ({signal_7763, signal_4372}), .b ({signal_10915, signal_7329}), .c ({signal_11150, signal_7433}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7445 ( .a ({signal_7742, signal_4373}), .b ({signal_10916, signal_7330}), .c ({signal_11151, signal_7434}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7446 ( .a ({signal_7721, signal_4374}), .b ({signal_10917, signal_4214}), .c ({signal_11152, signal_4246}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7447 ( .a ({signal_7688, signal_4375}), .b ({signal_10918, signal_4215}), .c ({signal_11153, signal_4247}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7448 ( .a ({signal_7655, signal_4376}), .b ({signal_10919, signal_4216}), .c ({signal_11154, signal_4248}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7449 ( .a ({signal_7634, signal_4355}), .b ({signal_10920, signal_4195}), .c ({signal_11155, signal_4227}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7450 ( .a ({signal_7631, signal_4356}), .b ({signal_10921, signal_7331}), .c ({signal_11156, signal_7435}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7451 ( .a ({signal_7628, signal_4357}), .b ({signal_10922, signal_7332}), .c ({signal_11157, signal_7436}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7452 ( .a ({signal_7625, signal_4358}), .b ({signal_10923, signal_4198}), .c ({signal_11158, signal_4230}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7453 ( .a ({signal_7622, signal_4377}), .b ({signal_10924, signal_7333}), .c ({signal_11159, signal_7437}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7454 ( .a ({signal_7619, signal_4359}), .b ({signal_10925, signal_4199}), .c ({signal_11160, signal_4231}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7455 ( .a ({signal_7616, signal_4360}), .b ({signal_10926, signal_4200}), .c ({signal_11161, signal_4232}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7456 ( .a ({signal_7613, signal_4361}), .b ({signal_10927, signal_7334}), .c ({signal_11162, signal_7438}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7457 ( .a ({signal_7607, signal_4363}), .b ({signal_10929, signal_4203}), .c ({signal_11163, signal_4235}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7458 ( .a ({signal_7604, signal_4364}), .b ({signal_10930, signal_7336}), .c ({signal_11164, signal_7439}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7459 ( .a ({signal_7601, signal_4365}), .b ({signal_10931, signal_7337}), .c ({signal_11165, signal_7440}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7460 ( .a ({signal_7598, signal_4366}), .b ({signal_10932, signal_4206}), .c ({signal_11166, signal_4238}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7461 ( .a ({signal_7595, signal_4367}), .b ({signal_10933, signal_4207}), .c ({signal_11167, signal_4239}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7462 ( .a ({signal_7562, signal_4368}), .b ({signal_10934, signal_4208}), .c ({signal_11168, signal_4240}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7463 ( .a ({signal_11024, signal_7340}), .b ({signal_11276, signal_4018}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7464 ( .a ({signal_11026, signal_7341}), .b ({signal_11277, signal_4020}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7465 ( .a ({signal_11027, signal_7342}), .b ({signal_11278, signal_4021}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7466 ( .a ({signal_11031, signal_7345}), .b ({signal_11279, signal_3996}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7467 ( .a ({signal_11033, signal_7346}), .b ({signal_11280, signal_3997}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7468 ( .a ({signal_11039, signal_7350}), .b ({signal_11281, signal_4004}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7469 ( .a ({signal_11040, signal_7351}), .b ({signal_11282, signal_4005}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7470 ( .a ({signal_11046, signal_7356}), .b ({signal_11283, signal_4010}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7471 ( .a ({signal_11048, signal_7357}), .b ({signal_11284, signal_4012}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7472 ( .a ({signal_11049, signal_7358}), .b ({signal_11285, signal_4013}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7473 ( .a ({signal_11053, signal_7361}), .b ({signal_11286, signal_4026}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7474 ( .a ({signal_11055, signal_7363}), .b ({signal_11287, signal_4050}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7475 ( .a ({signal_11057, signal_7364}), .b ({signal_11288, signal_4052}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7476 ( .a ({signal_11058, signal_7365}), .b ({signal_11289, signal_4053}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7477 ( .a ({signal_11062, signal_7368}), .b ({signal_11290, signal_4028}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7478 ( .a ({signal_11064, signal_7369}), .b ({signal_11291, signal_4029}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7479 ( .a ({signal_11070, signal_7373}), .b ({signal_11292, signal_4036}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7480 ( .a ({signal_11071, signal_7374}), .b ({signal_11293, signal_4037}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7481 ( .a ({signal_11077, signal_7379}), .b ({signal_11294, signal_4042}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7482 ( .a ({signal_11079, signal_7380}), .b ({signal_11295, signal_4044}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7483 ( .a ({signal_11080, signal_7381}), .b ({signal_11296, signal_4045}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7484 ( .a ({signal_11084, signal_7384}), .b ({signal_11297, signal_4058}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7485 ( .a ({signal_11086, signal_7386}), .b ({signal_11298, signal_4082}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7486 ( .a ({signal_11088, signal_7387}), .b ({signal_11299, signal_4084}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7487 ( .a ({signal_11089, signal_7388}), .b ({signal_11300, signal_4085}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7488 ( .a ({signal_11093, signal_7391}), .b ({signal_11301, signal_4060}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7489 ( .a ({signal_11095, signal_7392}), .b ({signal_11302, signal_4061}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7490 ( .a ({signal_11101, signal_7396}), .b ({signal_11303, signal_4068}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7491 ( .a ({signal_11102, signal_7397}), .b ({signal_11304, signal_4069}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7492 ( .a ({signal_11108, signal_7402}), .b ({signal_11305, signal_4074}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7493 ( .a ({signal_11110, signal_7403}), .b ({signal_11306, signal_4076}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7494 ( .a ({signal_11111, signal_7404}), .b ({signal_11307, signal_4077}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7495 ( .a ({signal_11115, signal_7407}), .b ({signal_11308, signal_4090}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7496 ( .a ({signal_11117, signal_7409}), .b ({signal_11309, signal_4114}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7497 ( .a ({signal_11119, signal_7410}), .b ({signal_11310, signal_4116}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7498 ( .a ({signal_11120, signal_7411}), .b ({signal_11311, signal_4117}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7499 ( .a ({signal_11124, signal_7414}), .b ({signal_11312, signal_4092}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7500 ( .a ({signal_11126, signal_7415}), .b ({signal_11313, signal_4093}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7501 ( .a ({signal_11131, signal_7419}), .b ({signal_11314, signal_4098}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7502 ( .a ({signal_11133, signal_7420}), .b ({signal_11315, signal_4100}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7503 ( .a ({signal_11134, signal_7421}), .b ({signal_11316, signal_4101}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7504 ( .a ({signal_11140, signal_7426}), .b ({signal_11317, signal_4106}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7505 ( .a ({signal_11142, signal_7427}), .b ({signal_11318, signal_4108}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7506 ( .a ({signal_11143, signal_7428}), .b ({signal_11319, signal_4109}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7507 ( .a ({signal_11147, signal_7431}), .b ({signal_11320, signal_4122}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7508 ( .a ({signal_11148, signal_7432}), .b ({signal_11321, signal_4241}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7509 ( .a ({signal_11150, signal_7433}), .b ({signal_11322, signal_4244}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7510 ( .a ({signal_11151, signal_7434}), .b ({signal_11323, signal_4245}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7511 ( .a ({signal_11156, signal_7435}), .b ({signal_11324, signal_4228}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7512 ( .a ({signal_11157, signal_7436}), .b ({signal_11325, signal_4229}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7513 ( .a ({signal_11159, signal_7437}), .b ({signal_11326, signal_4249}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7514 ( .a ({signal_11162, signal_7438}), .b ({signal_11327, signal_4233}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7515 ( .a ({signal_11164, signal_7439}), .b ({signal_11328, signal_4236}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7516 ( .a ({signal_11165, signal_7440}), .b ({signal_11329, signal_4237}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7517 ( .a ({signal_10410, signal_7034}), .b ({signal_11023, signal_7339}), .c ({signal_11330, signal_7441}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7518 ( .a ({signal_10772, signal_7071}), .b ({signal_11028, signal_7343}), .c ({signal_11331, signal_4022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7519 ( .a ({signal_10773, signal_7072}), .b ({signal_11029, signal_7344}), .c ({signal_11332, signal_4023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7520 ( .a ({signal_10772, signal_7071}), .b ({signal_11034, signal_7347}), .c ({signal_11333, signal_3998}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7521 ( .a ({signal_10773, signal_7072}), .b ({signal_11035, signal_7348}), .c ({signal_11334, signal_3999}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7522 ( .a ({signal_10775, signal_7078}), .b ({signal_11037, signal_7349}), .c ({signal_11335, signal_7442}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7523 ( .a ({signal_10808, signal_7221}), .b ({signal_11041, signal_7352}), .c ({signal_11336, signal_4006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7524 ( .a ({signal_10775, signal_7078}), .b ({signal_11042, signal_7353}), .c ({signal_11337, signal_7443}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7525 ( .a ({signal_10810, signal_7223}), .b ({signal_11043, signal_7354}), .c ({signal_11338, signal_4007}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7526 ( .a ({signal_10812, signal_7225}), .b ({signal_11045, signal_7355}), .c ({signal_11339, signal_7444}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7527 ( .a ({signal_10818, signal_7231}), .b ({signal_11050, signal_7359}), .c ({signal_11340, signal_4014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7528 ( .a ({signal_10820, signal_7233}), .b ({signal_11051, signal_7360}), .c ({signal_11341, signal_4015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7529 ( .a ({signal_10389, signal_7025}), .b ({signal_11054, signal_7362}), .c ({signal_11342, signal_7445}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7530 ( .a ({signal_10776, signal_7103}), .b ({signal_11059, signal_7366}), .c ({signal_11343, signal_4054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7531 ( .a ({signal_10777, signal_7104}), .b ({signal_11060, signal_7367}), .c ({signal_11344, signal_4055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7532 ( .a ({signal_10776, signal_7103}), .b ({signal_11065, signal_7370}), .c ({signal_11345, signal_4030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7533 ( .a ({signal_10777, signal_7104}), .b ({signal_11066, signal_7371}), .c ({signal_11346, signal_4031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7534 ( .a ({signal_10779, signal_7110}), .b ({signal_11068, signal_7372}), .c ({signal_11347, signal_7446}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7535 ( .a ({signal_10836, signal_7250}), .b ({signal_11072, signal_7375}), .c ({signal_11348, signal_4038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7536 ( .a ({signal_10779, signal_7110}), .b ({signal_11073, signal_7376}), .c ({signal_11349, signal_7447}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7537 ( .a ({signal_10838, signal_7252}), .b ({signal_11074, signal_7377}), .c ({signal_11350, signal_4039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7538 ( .a ({signal_10840, signal_7254}), .b ({signal_11076, signal_7378}), .c ({signal_11351, signal_7448}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7539 ( .a ({signal_10846, signal_7260}), .b ({signal_11081, signal_7382}), .c ({signal_11352, signal_4046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7540 ( .a ({signal_10848, signal_7262}), .b ({signal_11082, signal_7383}), .c ({signal_11353, signal_4047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7541 ( .a ({signal_10361, signal_7013}), .b ({signal_11085, signal_7385}), .c ({signal_11354, signal_7449}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7542 ( .a ({signal_10780, signal_7135}), .b ({signal_11090, signal_7389}), .c ({signal_11355, signal_4086}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7543 ( .a ({signal_10781, signal_7136}), .b ({signal_11091, signal_7390}), .c ({signal_11356, signal_4087}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7544 ( .a ({signal_10780, signal_7135}), .b ({signal_11096, signal_7393}), .c ({signal_11357, signal_4062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7545 ( .a ({signal_10781, signal_7136}), .b ({signal_11097, signal_7394}), .c ({signal_11358, signal_4063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7546 ( .a ({signal_10783, signal_7142}), .b ({signal_11099, signal_7395}), .c ({signal_11359, signal_7450}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7547 ( .a ({signal_10864, signal_7279}), .b ({signal_11103, signal_7398}), .c ({signal_11360, signal_4070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7548 ( .a ({signal_10783, signal_7142}), .b ({signal_11104, signal_7399}), .c ({signal_11361, signal_7451}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7549 ( .a ({signal_10866, signal_7281}), .b ({signal_11105, signal_7400}), .c ({signal_11362, signal_4071}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7550 ( .a ({signal_10868, signal_7283}), .b ({signal_11107, signal_7401}), .c ({signal_11363, signal_7452}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7551 ( .a ({signal_10874, signal_7289}), .b ({signal_11112, signal_7405}), .c ({signal_11364, signal_4078}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7552 ( .a ({signal_10876, signal_7291}), .b ({signal_11113, signal_7406}), .c ({signal_11365, signal_4079}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7553 ( .a ({signal_10431, signal_7043}), .b ({signal_11116, signal_7408}), .c ({signal_11366, signal_7453}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7554 ( .a ({signal_10888, signal_7303}), .b ({signal_11121, signal_7412}), .c ({signal_11367, signal_4118}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7555 ( .a ({signal_10889, signal_7304}), .b ({signal_11122, signal_7413}), .c ({signal_11368, signal_4119}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7556 ( .a ({signal_10888, signal_7303}), .b ({signal_11127, signal_7416}), .c ({signal_11369, signal_4094}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7557 ( .a ({signal_10889, signal_7304}), .b ({signal_11128, signal_7417}), .c ({signal_11370, signal_4095}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7558 ( .a ({signal_10896, signal_7311}), .b ({signal_11130, signal_7418}), .c ({signal_11371, signal_7454}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7559 ( .a ({signal_10895, signal_7310}), .b ({signal_11135, signal_7422}), .c ({signal_11372, signal_4102}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7560 ( .a ({signal_10896, signal_7311}), .b ({signal_11136, signal_7423}), .c ({signal_11373, signal_7455}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7561 ( .a ({signal_10898, signal_7313}), .b ({signal_11137, signal_7424}), .c ({signal_11374, signal_4103}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7562 ( .a ({signal_10900, signal_7315}), .b ({signal_11139, signal_7425}), .c ({signal_11375, signal_7456}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7563 ( .a ({signal_10906, signal_7321}), .b ({signal_11144, signal_7429}), .c ({signal_11376, signal_4110}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_7564 ( .a ({signal_10908, signal_7323}), .b ({signal_11145, signal_7430}), .c ({signal_11377, signal_4111}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7565 ( .a ({signal_11330, signal_7441}), .b ({signal_11559, signal_4017}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7566 ( .a ({signal_11335, signal_7442}), .b ({signal_11560, signal_4001}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7567 ( .a ({signal_11337, signal_7443}), .b ({signal_11561, signal_4025}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7568 ( .a ({signal_11339, signal_7444}), .b ({signal_11562, signal_4009}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7569 ( .a ({signal_11342, signal_7445}), .b ({signal_11563, signal_4049}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7570 ( .a ({signal_11347, signal_7446}), .b ({signal_11564, signal_4033}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7571 ( .a ({signal_11349, signal_7447}), .b ({signal_11565, signal_4057}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7572 ( .a ({signal_11351, signal_7448}), .b ({signal_11566, signal_4041}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7573 ( .a ({signal_11354, signal_7449}), .b ({signal_11567, signal_4081}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7574 ( .a ({signal_11359, signal_7450}), .b ({signal_11568, signal_4065}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7575 ( .a ({signal_11361, signal_7451}), .b ({signal_11569, signal_4089}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7576 ( .a ({signal_11363, signal_7452}), .b ({signal_11570, signal_4073}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7577 ( .a ({signal_11366, signal_7453}), .b ({signal_11571, signal_4113}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7578 ( .a ({signal_11371, signal_7454}), .b ({signal_11572, signal_4097}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7579 ( .a ({signal_11373, signal_7455}), .b ({signal_11573, signal_4121}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_7580 ( .a ({signal_11375, signal_7456}), .b ({signal_11574, signal_4105}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_293 ( .clk (signal_12469), .D ({signal_11592, signal_421}), .Q ({signal_7530, signal_3870}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_296 ( .clk (signal_12469), .D ({signal_11758, signal_423}), .Q ({signal_7623, signal_3869}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_299 ( .clk (signal_12469), .D ({signal_11459, signal_425}), .Q ({signal_7656, signal_3868}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_302 ( .clk (signal_12469), .D ({signal_11594, signal_427}), .Q ({signal_7689, signal_3867}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_305 ( .clk (signal_12469), .D ({signal_11596, signal_429}), .Q ({signal_7722, signal_3866}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_308 ( .clk (signal_12469), .D ({signal_11598, signal_431}), .Q ({signal_7743, signal_3865}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_311 ( .clk (signal_12469), .D ({signal_11600, signal_433}), .Q ({signal_7764, signal_3864}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_314 ( .clk (signal_12469), .D ({signal_11461, signal_435}), .Q ({signal_7797, signal_3863}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_317 ( .clk (signal_12469), .D ({signal_11602, signal_437}), .Q ({signal_7824, signal_3862}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_320 ( .clk (signal_12469), .D ({signal_11760, signal_439}), .Q ({signal_7839, signal_3861}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_323 ( .clk (signal_12469), .D ({signal_11463, signal_441}), .Q ({signal_7563, signal_3860}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_326 ( .clk (signal_12469), .D ({signal_11604, signal_443}), .Q ({signal_7596, signal_3859}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_329 ( .clk (signal_12469), .D ({signal_11606, signal_445}), .Q ({signal_7599, signal_3858}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_332 ( .clk (signal_12469), .D ({signal_11608, signal_447}), .Q ({signal_7602, signal_3857}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_335 ( .clk (signal_12469), .D ({signal_11610, signal_449}), .Q ({signal_7605, signal_3856}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_338 ( .clk (signal_12469), .D ({signal_11465, signal_451}), .Q ({signal_7608, signal_3855}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_341 ( .clk (signal_12469), .D ({signal_11612, signal_453}), .Q ({signal_7611, signal_3854}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_344 ( .clk (signal_12469), .D ({signal_11762, signal_455}), .Q ({signal_7614, signal_3853}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_347 ( .clk (signal_12469), .D ({signal_11467, signal_457}), .Q ({signal_7617, signal_3852}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_350 ( .clk (signal_12469), .D ({signal_11614, signal_459}), .Q ({signal_7620, signal_3851}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_353 ( .clk (signal_12469), .D ({signal_11616, signal_461}), .Q ({signal_7626, signal_3850}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_356 ( .clk (signal_12469), .D ({signal_11618, signal_463}), .Q ({signal_7629, signal_3849}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_359 ( .clk (signal_12469), .D ({signal_11620, signal_465}), .Q ({signal_7632, signal_3848}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_362 ( .clk (signal_12469), .D ({signal_11469, signal_467}), .Q ({signal_7635, signal_3847}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_365 ( .clk (signal_12469), .D ({signal_11622, signal_469}), .Q ({signal_7638, signal_3846}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_368 ( .clk (signal_12469), .D ({signal_11764, signal_471}), .Q ({signal_7641, signal_3845}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_371 ( .clk (signal_12469), .D ({signal_11471, signal_473}), .Q ({signal_7644, signal_3844}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_374 ( .clk (signal_12469), .D ({signal_11624, signal_475}), .Q ({signal_7647, signal_3843}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_377 ( .clk (signal_12469), .D ({signal_11626, signal_477}), .Q ({signal_7650, signal_3842}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_380 ( .clk (signal_12469), .D ({signal_11628, signal_479}), .Q ({signal_7653, signal_3841}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_383 ( .clk (signal_12469), .D ({signal_11630, signal_481}), .Q ({signal_7659, signal_3840}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_386 ( .clk (signal_12469), .D ({signal_11473, signal_483}), .Q ({signal_7662, signal_3839}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_389 ( .clk (signal_12469), .D ({signal_11632, signal_485}), .Q ({signal_7665, signal_3838}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_392 ( .clk (signal_12469), .D ({signal_11766, signal_487}), .Q ({signal_7668, signal_3837}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_395 ( .clk (signal_12469), .D ({signal_11475, signal_489}), .Q ({signal_7671, signal_3836}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_398 ( .clk (signal_12469), .D ({signal_11634, signal_491}), .Q ({signal_7674, signal_3835}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_401 ( .clk (signal_12469), .D ({signal_11636, signal_493}), .Q ({signal_7677, signal_3834}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_404 ( .clk (signal_12469), .D ({signal_11638, signal_495}), .Q ({signal_7680, signal_3833}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_407 ( .clk (signal_12469), .D ({signal_11640, signal_497}), .Q ({signal_7683, signal_3832}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_410 ( .clk (signal_12469), .D ({signal_11477, signal_499}), .Q ({signal_7686, signal_3831}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_413 ( .clk (signal_12469), .D ({signal_11642, signal_501}), .Q ({signal_7692, signal_3830}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_416 ( .clk (signal_12469), .D ({signal_11768, signal_503}), .Q ({signal_7695, signal_3829}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_419 ( .clk (signal_12469), .D ({signal_11479, signal_505}), .Q ({signal_7698, signal_3828}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_422 ( .clk (signal_12469), .D ({signal_11644, signal_507}), .Q ({signal_7701, signal_3827}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_425 ( .clk (signal_12469), .D ({signal_11646, signal_509}), .Q ({signal_7704, signal_3826}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_428 ( .clk (signal_12469), .D ({signal_11648, signal_511}), .Q ({signal_7707, signal_3825}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_431 ( .clk (signal_12469), .D ({signal_11650, signal_513}), .Q ({signal_7710, signal_3824}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_434 ( .clk (signal_12469), .D ({signal_11481, signal_515}), .Q ({signal_7713, signal_3823}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_437 ( .clk (signal_12469), .D ({signal_11652, signal_517}), .Q ({signal_7716, signal_3822}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_440 ( .clk (signal_12469), .D ({signal_11770, signal_519}), .Q ({signal_7719, signal_3821}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_443 ( .clk (signal_12469), .D ({signal_11483, signal_521}), .Q ({signal_7725, signal_3820}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_446 ( .clk (signal_12469), .D ({signal_11654, signal_523}), .Q ({signal_7728, signal_3819}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_449 ( .clk (signal_12469), .D ({signal_11656, signal_525}), .Q ({signal_7731, signal_3818}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_452 ( .clk (signal_12469), .D ({signal_11658, signal_527}), .Q ({signal_7734, signal_3817}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_455 ( .clk (signal_12469), .D ({signal_11660, signal_529}), .Q ({signal_7737, signal_3816}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_458 ( .clk (signal_12469), .D ({signal_11485, signal_531}), .Q ({signal_7740, signal_3815}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_461 ( .clk (signal_12469), .D ({signal_11662, signal_533}), .Q ({signal_7481, signal_3814}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_464 ( .clk (signal_12469), .D ({signal_11772, signal_535}), .Q ({signal_7484, signal_3813}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_467 ( .clk (signal_12469), .D ({signal_11487, signal_537}), .Q ({signal_7487, signal_3812}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_470 ( .clk (signal_12469), .D ({signal_11664, signal_539}), .Q ({signal_7490, signal_3811}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_473 ( .clk (signal_12469), .D ({signal_11666, signal_541}), .Q ({signal_7493, signal_3810}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_476 ( .clk (signal_12469), .D ({signal_11668, signal_543}), .Q ({signal_7496, signal_3809}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_479 ( .clk (signal_12469), .D ({signal_11670, signal_545}), .Q ({signal_7499, signal_3808}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_482 ( .clk (signal_12469), .D ({signal_11489, signal_547}), .Q ({signal_7502, signal_3807}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_485 ( .clk (signal_12469), .D ({signal_11672, signal_549}), .Q ({signal_7746, signal_3806}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_488 ( .clk (signal_12469), .D ({signal_11774, signal_551}), .Q ({signal_7749, signal_3805}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_491 ( .clk (signal_12469), .D ({signal_11491, signal_553}), .Q ({signal_7752, signal_3804}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_494 ( .clk (signal_12469), .D ({signal_11674, signal_555}), .Q ({signal_7755, signal_3803}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_497 ( .clk (signal_12469), .D ({signal_11676, signal_557}), .Q ({signal_7758, signal_3802}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_500 ( .clk (signal_12469), .D ({signal_11678, signal_559}), .Q ({signal_7761, signal_3801}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_503 ( .clk (signal_12469), .D ({signal_11680, signal_561}), .Q ({signal_7767, signal_3800}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_506 ( .clk (signal_12469), .D ({signal_11493, signal_563}), .Q ({signal_7770, signal_3799}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_509 ( .clk (signal_12469), .D ({signal_11682, signal_565}), .Q ({signal_7773, signal_3798}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_512 ( .clk (signal_12469), .D ({signal_11776, signal_567}), .Q ({signal_7776, signal_3797}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_515 ( .clk (signal_12469), .D ({signal_11495, signal_569}), .Q ({signal_7779, signal_3796}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_518 ( .clk (signal_12469), .D ({signal_11684, signal_571}), .Q ({signal_7782, signal_3795}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_521 ( .clk (signal_12469), .D ({signal_11686, signal_573}), .Q ({signal_7785, signal_3794}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_524 ( .clk (signal_12469), .D ({signal_11688, signal_575}), .Q ({signal_7788, signal_3793}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_527 ( .clk (signal_12469), .D ({signal_11690, signal_577}), .Q ({signal_7791, signal_3792}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_530 ( .clk (signal_12469), .D ({signal_11497, signal_579}), .Q ({signal_7794, signal_3791}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_533 ( .clk (signal_12469), .D ({signal_11692, signal_581}), .Q ({signal_7800, signal_3790}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_536 ( .clk (signal_12469), .D ({signal_11778, signal_583}), .Q ({signal_7803, signal_3789}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_539 ( .clk (signal_12469), .D ({signal_11499, signal_585}), .Q ({signal_7806, signal_3788}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_542 ( .clk (signal_12469), .D ({signal_11694, signal_587}), .Q ({signal_7809, signal_3787}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_545 ( .clk (signal_12469), .D ({signal_11696, signal_589}), .Q ({signal_7812, signal_3786}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_548 ( .clk (signal_12469), .D ({signal_11698, signal_591}), .Q ({signal_7815, signal_3785}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_551 ( .clk (signal_12469), .D ({signal_11700, signal_593}), .Q ({signal_7818, signal_3784}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_554 ( .clk (signal_12469), .D ({signal_11501, signal_595}), .Q ({signal_7821, signal_3783}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_557 ( .clk (signal_12469), .D ({signal_11702, signal_597}), .Q ({signal_7505, signal_3782}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_560 ( .clk (signal_12469), .D ({signal_11780, signal_599}), .Q ({signal_7508, signal_3781}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_563 ( .clk (signal_12469), .D ({signal_11503, signal_601}), .Q ({signal_7511, signal_3780}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_566 ( .clk (signal_12469), .D ({signal_11704, signal_603}), .Q ({signal_7514, signal_3779}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_569 ( .clk (signal_12469), .D ({signal_11706, signal_605}), .Q ({signal_7517, signal_3778}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_572 ( .clk (signal_12469), .D ({signal_11708, signal_607}), .Q ({signal_7520, signal_3777}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_575 ( .clk (signal_12469), .D ({signal_11710, signal_609}), .Q ({signal_7523, signal_3776}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_578 ( .clk (signal_12469), .D ({signal_11505, signal_611}), .Q ({signal_7526, signal_3775}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_581 ( .clk (signal_12469), .D ({signal_11712, signal_613}), .Q ({signal_7827, signal_3774}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_584 ( .clk (signal_12469), .D ({signal_11782, signal_615}), .Q ({signal_7830, signal_3773}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_587 ( .clk (signal_12469), .D ({signal_11507, signal_617}), .Q ({signal_7833, signal_3772}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_590 ( .clk (signal_12469), .D ({signal_11714, signal_619}), .Q ({signal_7836, signal_3771}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_593 ( .clk (signal_12469), .D ({signal_11716, signal_621}), .Q ({signal_7533, signal_3770}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_596 ( .clk (signal_12469), .D ({signal_11718, signal_623}), .Q ({signal_7536, signal_3769}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_599 ( .clk (signal_12469), .D ({signal_11720, signal_625}), .Q ({signal_7539, signal_3768}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_602 ( .clk (signal_12469), .D ({signal_11509, signal_627}), .Q ({signal_7542, signal_3767}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_605 ( .clk (signal_12469), .D ({signal_11722, signal_629}), .Q ({signal_7545, signal_3766}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_608 ( .clk (signal_12469), .D ({signal_11784, signal_631}), .Q ({signal_7548, signal_3765}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_611 ( .clk (signal_12469), .D ({signal_11511, signal_633}), .Q ({signal_7551, signal_3764}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_614 ( .clk (signal_12469), .D ({signal_11724, signal_635}), .Q ({signal_7554, signal_3763}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_617 ( .clk (signal_12469), .D ({signal_11726, signal_637}), .Q ({signal_7557, signal_3762}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_620 ( .clk (signal_12469), .D ({signal_11728, signal_639}), .Q ({signal_7560, signal_3761}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_623 ( .clk (signal_12469), .D ({signal_11730, signal_641}), .Q ({signal_7566, signal_3760}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_626 ( .clk (signal_12469), .D ({signal_11513, signal_643}), .Q ({signal_7569, signal_3759}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_629 ( .clk (signal_12469), .D ({signal_11732, signal_645}), .Q ({signal_7572, signal_3758}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_632 ( .clk (signal_12469), .D ({signal_11786, signal_647}), .Q ({signal_7575, signal_3757}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_635 ( .clk (signal_12469), .D ({signal_11515, signal_649}), .Q ({signal_7578, signal_3756}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_638 ( .clk (signal_12469), .D ({signal_11734, signal_651}), .Q ({signal_7581, signal_3755}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_641 ( .clk (signal_12469), .D ({signal_11736, signal_653}), .Q ({signal_7584, signal_3754}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_644 ( .clk (signal_12469), .D ({signal_11738, signal_655}), .Q ({signal_7587, signal_3753}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_647 ( .clk (signal_12469), .D ({signal_11740, signal_657}), .Q ({signal_7590, signal_3752}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_650 ( .clk (signal_12469), .D ({signal_11517, signal_659}), .Q ({signal_7593, signal_3751}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_653 ( .clk (signal_12469), .D ({signal_11742, signal_661}), .Q ({signal_7457, signal_3750}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_656 ( .clk (signal_12469), .D ({signal_11788, signal_663}), .Q ({signal_7460, signal_3749}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_659 ( .clk (signal_12469), .D ({signal_11519, signal_665}), .Q ({signal_7463, signal_3748}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_662 ( .clk (signal_12469), .D ({signal_11744, signal_667}), .Q ({signal_7466, signal_3747}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_665 ( .clk (signal_12469), .D ({signal_11746, signal_669}), .Q ({signal_7469, signal_3746}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_668 ( .clk (signal_12469), .D ({signal_11748, signal_671}), .Q ({signal_7472, signal_3745}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_671 ( .clk (signal_12469), .D ({signal_11750, signal_673}), .Q ({signal_7475, signal_3744}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_674 ( .clk (signal_12469), .D ({signal_11521, signal_675}), .Q ({signal_7478, signal_3743}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3157 ( .clk (signal_12469), .D ({signal_11202, signal_2853}), .Q ({signal_7529, signal_4378}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3160 ( .clk (signal_12469), .D ({signal_11523, signal_2855}), .Q ({signal_7622, signal_4377}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3163 ( .clk (signal_12469), .D ({signal_11204, signal_2857}), .Q ({signal_7655, signal_4376}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3166 ( .clk (signal_12469), .D ({signal_11206, signal_2859}), .Q ({signal_7688, signal_4375}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3169 ( .clk (signal_12469), .D ({signal_11208, signal_2861}), .Q ({signal_7721, signal_4374}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3172 ( .clk (signal_12469), .D ({signal_11525, signal_2863}), .Q ({signal_7742, signal_4373}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3175 ( .clk (signal_12469), .D ({signal_11527, signal_2865}), .Q ({signal_7763, signal_4372}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3178 ( .clk (signal_12469), .D ({signal_11210, signal_2867}), .Q ({signal_7796, signal_4371}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3181 ( .clk (signal_12469), .D ({signal_11212, signal_2869}), .Q ({signal_7823, signal_4370}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3184 ( .clk (signal_12469), .D ({signal_11529, signal_2871}), .Q ({signal_7838, signal_4369}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3187 ( .clk (signal_12469), .D ({signal_11214, signal_2873}), .Q ({signal_7562, signal_4368}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3190 ( .clk (signal_12469), .D ({signal_11216, signal_2875}), .Q ({signal_7595, signal_4367}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3193 ( .clk (signal_12469), .D ({signal_11218, signal_2877}), .Q ({signal_7598, signal_4366}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3196 ( .clk (signal_12469), .D ({signal_11531, signal_2879}), .Q ({signal_7601, signal_4365}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3199 ( .clk (signal_12469), .D ({signal_11533, signal_2881}), .Q ({signal_7604, signal_4364}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3202 ( .clk (signal_12469), .D ({signal_11220, signal_2883}), .Q ({signal_7607, signal_4363}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3205 ( .clk (signal_12469), .D ({signal_11222, signal_2885}), .Q ({signal_7610, signal_4362}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3208 ( .clk (signal_12469), .D ({signal_11535, signal_2887}), .Q ({signal_7613, signal_4361}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3211 ( .clk (signal_12469), .D ({signal_11224, signal_2889}), .Q ({signal_7616, signal_4360}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3214 ( .clk (signal_12469), .D ({signal_11226, signal_2891}), .Q ({signal_7619, signal_4359}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3217 ( .clk (signal_12469), .D ({signal_11228, signal_2893}), .Q ({signal_7625, signal_4358}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3220 ( .clk (signal_12469), .D ({signal_11537, signal_2895}), .Q ({signal_7628, signal_4357}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3223 ( .clk (signal_12469), .D ({signal_11539, signal_2897}), .Q ({signal_7631, signal_4356}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3226 ( .clk (signal_12469), .D ({signal_11230, signal_2899}), .Q ({signal_7634, signal_4355}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3229 ( .clk (signal_12469), .D ({signal_11541, signal_2901}), .Q ({signal_7637, signal_4354}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3232 ( .clk (signal_12469), .D ({signal_11752, signal_2903}), .Q ({signal_7640, signal_4353}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3235 ( .clk (signal_12469), .D ({signal_11543, signal_2905}), .Q ({signal_7643, signal_4352}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3238 ( .clk (signal_12469), .D ({signal_11545, signal_2907}), .Q ({signal_7646, signal_4351}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3241 ( .clk (signal_12469), .D ({signal_11547, signal_2909}), .Q ({signal_7649, signal_4350}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3244 ( .clk (signal_12469), .D ({signal_11754, signal_2911}), .Q ({signal_7652, signal_4349}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3247 ( .clk (signal_12469), .D ({signal_11756, signal_2913}), .Q ({signal_7658, signal_4348}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3250 ( .clk (signal_12469), .D ({signal_11549, signal_2915}), .Q ({signal_7661, signal_4347}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3253 ( .clk (signal_12469), .D ({signal_10937, signal_2917}), .Q ({signal_7664, signal_4346}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3256 ( .clk (signal_12469), .D ({signal_11232, signal_2919}), .Q ({signal_7667, signal_4345}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3259 ( .clk (signal_12469), .D ({signal_10939, signal_2921}), .Q ({signal_7670, signal_4344}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3262 ( .clk (signal_12469), .D ({signal_10941, signal_2923}), .Q ({signal_7673, signal_4343}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3265 ( .clk (signal_12469), .D ({signal_10943, signal_2925}), .Q ({signal_7676, signal_4342}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3268 ( .clk (signal_12469), .D ({signal_11234, signal_2927}), .Q ({signal_7679, signal_4341}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3271 ( .clk (signal_12469), .D ({signal_11236, signal_2929}), .Q ({signal_7682, signal_4340}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3274 ( .clk (signal_12469), .D ({signal_10945, signal_2931}), .Q ({signal_7685, signal_4339}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3277 ( .clk (signal_12469), .D ({signal_10947, signal_2933}), .Q ({signal_7691, signal_4338}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3280 ( .clk (signal_12469), .D ({signal_11238, signal_2935}), .Q ({signal_7694, signal_4337}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3283 ( .clk (signal_12469), .D ({signal_10949, signal_2937}), .Q ({signal_7697, signal_4336}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3286 ( .clk (signal_12469), .D ({signal_10951, signal_2939}), .Q ({signal_7700, signal_4335}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3289 ( .clk (signal_12469), .D ({signal_10953, signal_2941}), .Q ({signal_7703, signal_4334}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3292 ( .clk (signal_12469), .D ({signal_11240, signal_2943}), .Q ({signal_7706, signal_4333}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3295 ( .clk (signal_12469), .D ({signal_11242, signal_2945}), .Q ({signal_7709, signal_4332}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3298 ( .clk (signal_12469), .D ({signal_10955, signal_2947}), .Q ({signal_7712, signal_4331}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3301 ( .clk (signal_12469), .D ({signal_10957, signal_2949}), .Q ({signal_7715, signal_4330}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3304 ( .clk (signal_12469), .D ({signal_11244, signal_2951}), .Q ({signal_7718, signal_4329}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3307 ( .clk (signal_12469), .D ({signal_10959, signal_2953}), .Q ({signal_7724, signal_4328}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3310 ( .clk (signal_12469), .D ({signal_10961, signal_2955}), .Q ({signal_7727, signal_4327}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3313 ( .clk (signal_12469), .D ({signal_10963, signal_2957}), .Q ({signal_7730, signal_4326}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3316 ( .clk (signal_12469), .D ({signal_11246, signal_2959}), .Q ({signal_7733, signal_4325}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3319 ( .clk (signal_12469), .D ({signal_11248, signal_2961}), .Q ({signal_7736, signal_4324}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3322 ( .clk (signal_12469), .D ({signal_10965, signal_2963}), .Q ({signal_7739, signal_4323}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3325 ( .clk (signal_12469), .D ({signal_11250, signal_2965}), .Q ({signal_7482, signal_4322}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3328 ( .clk (signal_12469), .D ({signal_11551, signal_2967}), .Q ({signal_7485, signal_4321}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3331 ( .clk (signal_12469), .D ({signal_11252, signal_2969}), .Q ({signal_7488, signal_4320}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3334 ( .clk (signal_12469), .D ({signal_11254, signal_2971}), .Q ({signal_7491, signal_4319}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3337 ( .clk (signal_12469), .D ({signal_11256, signal_2973}), .Q ({signal_7494, signal_4318}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3340 ( .clk (signal_12469), .D ({signal_11553, signal_2975}), .Q ({signal_7497, signal_4317}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3343 ( .clk (signal_12469), .D ({signal_11555, signal_2977}), .Q ({signal_7500, signal_4316}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3346 ( .clk (signal_12469), .D ({signal_11258, signal_2979}), .Q ({signal_7503, signal_4315}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3349 ( .clk (signal_12469), .D ({signal_10707, signal_2981}), .Q ({signal_7745, signal_4314}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3352 ( .clk (signal_12469), .D ({signal_10967, signal_2983}), .Q ({signal_7748, signal_4313}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3355 ( .clk (signal_12469), .D ({signal_10709, signal_2985}), .Q ({signal_7751, signal_4312}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3358 ( .clk (signal_12469), .D ({signal_10711, signal_2987}), .Q ({signal_7754, signal_4311}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3361 ( .clk (signal_12469), .D ({signal_10713, signal_2989}), .Q ({signal_7757, signal_4310}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3364 ( .clk (signal_12469), .D ({signal_10969, signal_2991}), .Q ({signal_7760, signal_4309}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3367 ( .clk (signal_12469), .D ({signal_10971, signal_2993}), .Q ({signal_7766, signal_4308}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3370 ( .clk (signal_12469), .D ({signal_10715, signal_2995}), .Q ({signal_7769, signal_4307}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3373 ( .clk (signal_12469), .D ({signal_10717, signal_2997}), .Q ({signal_7772, signal_4306}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3376 ( .clk (signal_12469), .D ({signal_10973, signal_2999}), .Q ({signal_7775, signal_4305}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3379 ( .clk (signal_12469), .D ({signal_10719, signal_3001}), .Q ({signal_7778, signal_4304}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3382 ( .clk (signal_12469), .D ({signal_10721, signal_3003}), .Q ({signal_7781, signal_4303}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3385 ( .clk (signal_12469), .D ({signal_10723, signal_3005}), .Q ({signal_7784, signal_4302}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3388 ( .clk (signal_12469), .D ({signal_10975, signal_3007}), .Q ({signal_7787, signal_4301}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3391 ( .clk (signal_12469), .D ({signal_10977, signal_3009}), .Q ({signal_7790, signal_4300}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3394 ( .clk (signal_12469), .D ({signal_10725, signal_3011}), .Q ({signal_7793, signal_4299}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3397 ( .clk (signal_12469), .D ({signal_10727, signal_3013}), .Q ({signal_7799, signal_4298}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3400 ( .clk (signal_12469), .D ({signal_10979, signal_3015}), .Q ({signal_7802, signal_4297}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3403 ( .clk (signal_12469), .D ({signal_10729, signal_3017}), .Q ({signal_7805, signal_4296}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3406 ( .clk (signal_12469), .D ({signal_10731, signal_3019}), .Q ({signal_7808, signal_4295}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3409 ( .clk (signal_12469), .D ({signal_10733, signal_3021}), .Q ({signal_7811, signal_4294}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3412 ( .clk (signal_12469), .D ({signal_10981, signal_3023}), .Q ({signal_7814, signal_4293}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3415 ( .clk (signal_12469), .D ({signal_10983, signal_3025}), .Q ({signal_7817, signal_4292}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3418 ( .clk (signal_12469), .D ({signal_10735, signal_3027}), .Q ({signal_7820, signal_4291}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3421 ( .clk (signal_12469), .D ({signal_10985, signal_3029}), .Q ({signal_7506, signal_4290}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3424 ( .clk (signal_12469), .D ({signal_11260, signal_3031}), .Q ({signal_7509, signal_4289}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3427 ( .clk (signal_12469), .D ({signal_10987, signal_3033}), .Q ({signal_7512, signal_4288}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3430 ( .clk (signal_12469), .D ({signal_10989, signal_3035}), .Q ({signal_7515, signal_4287}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3433 ( .clk (signal_12469), .D ({signal_10991, signal_3037}), .Q ({signal_7518, signal_4286}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3436 ( .clk (signal_12469), .D ({signal_11262, signal_3039}), .Q ({signal_7521, signal_4285}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3439 ( .clk (signal_12469), .D ({signal_11264, signal_3041}), .Q ({signal_7524, signal_4284}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3442 ( .clk (signal_12469), .D ({signal_10993, signal_3043}), .Q ({signal_7527, signal_4283}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3445 ( .clk (signal_12469), .D ({signal_10457, signal_3045}), .Q ({signal_7826, signal_4282}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3448 ( .clk (signal_12469), .D ({signal_10737, signal_3047}), .Q ({signal_7829, signal_4281}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3451 ( .clk (signal_12469), .D ({signal_10459, signal_3049}), .Q ({signal_7832, signal_4280}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3454 ( .clk (signal_12469), .D ({signal_10461, signal_3051}), .Q ({signal_7835, signal_4279}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3457 ( .clk (signal_12469), .D ({signal_10463, signal_3053}), .Q ({signal_7532, signal_4278}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3460 ( .clk (signal_12469), .D ({signal_10739, signal_3055}), .Q ({signal_7535, signal_4277}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3463 ( .clk (signal_12469), .D ({signal_10741, signal_3057}), .Q ({signal_7538, signal_4276}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3466 ( .clk (signal_12469), .D ({signal_10465, signal_3059}), .Q ({signal_7541, signal_4275}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3469 ( .clk (signal_12469), .D ({signal_10467, signal_3061}), .Q ({signal_7544, signal_4274}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3472 ( .clk (signal_12469), .D ({signal_10743, signal_3063}), .Q ({signal_7547, signal_4273}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3475 ( .clk (signal_12469), .D ({signal_10469, signal_3065}), .Q ({signal_7550, signal_4272}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3478 ( .clk (signal_12469), .D ({signal_10471, signal_3067}), .Q ({signal_7553, signal_4271}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3481 ( .clk (signal_12469), .D ({signal_10473, signal_3069}), .Q ({signal_7556, signal_4270}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3484 ( .clk (signal_12469), .D ({signal_10745, signal_3071}), .Q ({signal_7559, signal_4269}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3487 ( .clk (signal_12469), .D ({signal_10747, signal_3073}), .Q ({signal_7565, signal_4268}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3490 ( .clk (signal_12469), .D ({signal_10475, signal_3075}), .Q ({signal_7568, signal_4267}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3493 ( .clk (signal_12469), .D ({signal_10477, signal_3077}), .Q ({signal_7571, signal_4266}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3496 ( .clk (signal_12469), .D ({signal_10749, signal_3079}), .Q ({signal_7574, signal_4265}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3499 ( .clk (signal_12469), .D ({signal_10479, signal_3081}), .Q ({signal_7577, signal_4264}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3502 ( .clk (signal_12469), .D ({signal_10481, signal_3083}), .Q ({signal_7580, signal_4263}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3505 ( .clk (signal_12469), .D ({signal_10483, signal_3085}), .Q ({signal_7583, signal_4262}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3508 ( .clk (signal_12469), .D ({signal_10751, signal_3087}), .Q ({signal_7586, signal_4261}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3511 ( .clk (signal_12469), .D ({signal_10753, signal_3089}), .Q ({signal_7589, signal_4260}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3514 ( .clk (signal_12469), .D ({signal_10485, signal_3091}), .Q ({signal_7592, signal_4259}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3517 ( .clk (signal_12469), .D ({signal_10755, signal_3093}), .Q ({signal_7458, signal_4258}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3520 ( .clk (signal_12469), .D ({signal_10995, signal_3095}), .Q ({signal_7461, signal_4257}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3523 ( .clk (signal_12469), .D ({signal_10757, signal_3097}), .Q ({signal_7464, signal_4256}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3526 ( .clk (signal_12469), .D ({signal_10759, signal_3099}), .Q ({signal_7467, signal_4255}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3529 ( .clk (signal_12469), .D ({signal_10761, signal_3101}), .Q ({signal_7470, signal_4254}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3532 ( .clk (signal_12469), .D ({signal_10997, signal_3103}), .Q ({signal_7473, signal_4253}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3535 ( .clk (signal_12469), .D ({signal_10999, signal_3105}), .Q ({signal_7476, signal_4252}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3538 ( .clk (signal_12469), .D ({signal_10763, signal_3107}), .Q ({signal_7479, signal_4251}) ) ;
    DFF_X1 cell_4202 ( .CK (signal_12469), .D (signal_3612), .Q (signal_4388), .QN () ) ;
    DFF_X1 cell_4204 ( .CK (signal_12469), .D (signal_3610), .Q (signal_4387), .QN () ) ;
    DFF_X1 cell_4206 ( .CK (signal_12469), .D (signal_3607), .Q (signal_4386), .QN () ) ;
    DFF_X1 cell_4208 ( .CK (signal_12469), .D (signal_3608), .Q (signal_4385), .QN () ) ;
endmodule
