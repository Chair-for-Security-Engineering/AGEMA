/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 10 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 11 register stage(s) in total */

module sbox_HPC2_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [3:0] SI_s3 ;
    input [77:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    output [3:0] SO_s3 ;
    wire N9 ;
    wire N12 ;
    wire N19 ;
    wire N27 ;
    wire n40 ;
    wire n41 ;
    wire n42 ;
    wire n43 ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire new_AGEMA_signal_37 ;
    wire new_AGEMA_signal_38 ;
    wire new_AGEMA_signal_39 ;
    wire new_AGEMA_signal_46 ;
    wire new_AGEMA_signal_47 ;
    wire new_AGEMA_signal_48 ;
    wire new_AGEMA_signal_52 ;
    wire new_AGEMA_signal_53 ;
    wire new_AGEMA_signal_54 ;
    wire new_AGEMA_signal_55 ;
    wire new_AGEMA_signal_56 ;
    wire new_AGEMA_signal_57 ;
    wire new_AGEMA_signal_58 ;
    wire new_AGEMA_signal_59 ;
    wire new_AGEMA_signal_60 ;
    wire new_AGEMA_signal_61 ;
    wire new_AGEMA_signal_62 ;
    wire new_AGEMA_signal_63 ;
    wire new_AGEMA_signal_64 ;
    wire new_AGEMA_signal_65 ;
    wire new_AGEMA_signal_66 ;
    wire new_AGEMA_signal_67 ;
    wire new_AGEMA_signal_68 ;
    wire new_AGEMA_signal_69 ;
    wire new_AGEMA_signal_70 ;
    wire new_AGEMA_signal_71 ;
    wire new_AGEMA_signal_72 ;
    wire new_AGEMA_signal_73 ;
    wire new_AGEMA_signal_74 ;
    wire new_AGEMA_signal_75 ;
    wire new_AGEMA_signal_76 ;
    wire new_AGEMA_signal_77 ;
    wire new_AGEMA_signal_78 ;
    wire new_AGEMA_signal_79 ;
    wire new_AGEMA_signal_80 ;
    wire new_AGEMA_signal_81 ;
    wire new_AGEMA_signal_82 ;
    wire new_AGEMA_signal_83 ;
    wire new_AGEMA_signal_84 ;
    wire new_AGEMA_signal_85 ;
    wire new_AGEMA_signal_86 ;
    wire new_AGEMA_signal_87 ;
    wire new_AGEMA_signal_88 ;
    wire new_AGEMA_signal_89 ;
    wire new_AGEMA_signal_90 ;
    wire new_AGEMA_signal_91 ;
    wire new_AGEMA_signal_92 ;
    wire new_AGEMA_signal_93 ;
    wire new_AGEMA_signal_94 ;
    wire new_AGEMA_signal_95 ;
    wire new_AGEMA_signal_96 ;
    wire new_AGEMA_signal_97 ;
    wire new_AGEMA_signal_98 ;
    wire new_AGEMA_signal_99 ;
    wire new_AGEMA_signal_100 ;
    wire new_AGEMA_signal_101 ;
    wire new_AGEMA_signal_102 ;
    wire new_AGEMA_signal_193 ;
    wire new_AGEMA_signal_194 ;
    wire new_AGEMA_signal_195 ;
    wire new_AGEMA_signal_196 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_201 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_206 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_213 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_224 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) U50 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_39, new_AGEMA_signal_38, new_AGEMA_signal_37, n53}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U53 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, n52}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U59 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n51}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_23 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_25 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_27 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_29 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( new_AGEMA_signal_199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_31 ( .C ( clk ), .D ( n53 ), .Q ( new_AGEMA_signal_201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_33 ( .C ( clk ), .D ( new_AGEMA_signal_37 ), .Q ( new_AGEMA_signal_203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_35 ( .C ( clk ), .D ( new_AGEMA_signal_38 ), .Q ( new_AGEMA_signal_205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_37 ( .C ( clk ), .D ( new_AGEMA_signal_39 ), .Q ( new_AGEMA_signal_207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_39 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_41 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_43 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_45 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( new_AGEMA_signal_215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_47 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_49 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_51 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_53 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( new_AGEMA_signal_223 ) ) ;

    /* cells in depth 2 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U51 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_48, new_AGEMA_signal_47, new_AGEMA_signal_46, n40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) U52 ( .a ({new_AGEMA_signal_48, new_AGEMA_signal_47, new_AGEMA_signal_46, n40}), .b ({new_AGEMA_signal_200, new_AGEMA_signal_198, new_AGEMA_signal_196, new_AGEMA_signal_194}), .c ({new_AGEMA_signal_66, new_AGEMA_signal_65, new_AGEMA_signal_64, N12}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U54 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, n52}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, n41}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(1)) U55 ( .a ({new_AGEMA_signal_208, new_AGEMA_signal_206, new_AGEMA_signal_204, new_AGEMA_signal_202}), .b ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, n41}), .c ({new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, n42}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U57 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_57, new_AGEMA_signal_56, new_AGEMA_signal_55, n43}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U60 ( .a ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n51}), .b ({new_AGEMA_signal_39, new_AGEMA_signal_38, new_AGEMA_signal_37, n53}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_75, new_AGEMA_signal_74, new_AGEMA_signal_73, n45}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U61 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, n48}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U67 ( .a ({new_AGEMA_signal_54, new_AGEMA_signal_53, new_AGEMA_signal_52, n52}), .b ({new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n51}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, n54}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) U68 ( .a ({new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, n54}), .b ({new_AGEMA_signal_208, new_AGEMA_signal_206, new_AGEMA_signal_204, new_AGEMA_signal_202}), .c ({new_AGEMA_signal_93, new_AGEMA_signal_92, new_AGEMA_signal_91, N9}) ) ;
    buf_clk new_AGEMA_reg_buffer_24 ( .C ( clk ), .D ( new_AGEMA_signal_193 ), .Q ( new_AGEMA_signal_194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_26 ( .C ( clk ), .D ( new_AGEMA_signal_195 ), .Q ( new_AGEMA_signal_196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_28 ( .C ( clk ), .D ( new_AGEMA_signal_197 ), .Q ( new_AGEMA_signal_198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_30 ( .C ( clk ), .D ( new_AGEMA_signal_199 ), .Q ( new_AGEMA_signal_200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_32 ( .C ( clk ), .D ( new_AGEMA_signal_201 ), .Q ( new_AGEMA_signal_202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_34 ( .C ( clk ), .D ( new_AGEMA_signal_203 ), .Q ( new_AGEMA_signal_204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_36 ( .C ( clk ), .D ( new_AGEMA_signal_205 ), .Q ( new_AGEMA_signal_206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_38 ( .C ( clk ), .D ( new_AGEMA_signal_207 ), .Q ( new_AGEMA_signal_208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_40 ( .C ( clk ), .D ( new_AGEMA_signal_209 ), .Q ( new_AGEMA_signal_210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_42 ( .C ( clk ), .D ( new_AGEMA_signal_211 ), .Q ( new_AGEMA_signal_212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_44 ( .C ( clk ), .D ( new_AGEMA_signal_213 ), .Q ( new_AGEMA_signal_214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_46 ( .C ( clk ), .D ( new_AGEMA_signal_215 ), .Q ( new_AGEMA_signal_216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_48 ( .C ( clk ), .D ( new_AGEMA_signal_217 ), .Q ( new_AGEMA_signal_218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_50 ( .C ( clk ), .D ( new_AGEMA_signal_219 ), .Q ( new_AGEMA_signal_220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_52 ( .C ( clk ), .D ( new_AGEMA_signal_221 ), .Q ( new_AGEMA_signal_222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_54 ( .C ( clk ), .D ( new_AGEMA_signal_223 ), .Q ( new_AGEMA_signal_224 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_55 ( .C ( clk ), .D ( n45 ), .Q ( new_AGEMA_signal_225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_57 ( .C ( clk ), .D ( new_AGEMA_signal_73 ), .Q ( new_AGEMA_signal_227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_59 ( .C ( clk ), .D ( new_AGEMA_signal_74 ), .Q ( new_AGEMA_signal_229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_61 ( .C ( clk ), .D ( new_AGEMA_signal_75 ), .Q ( new_AGEMA_signal_231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_63 ( .C ( clk ), .D ( new_AGEMA_signal_210 ), .Q ( new_AGEMA_signal_233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_67 ( .C ( clk ), .D ( new_AGEMA_signal_212 ), .Q ( new_AGEMA_signal_237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_71 ( .C ( clk ), .D ( new_AGEMA_signal_214 ), .Q ( new_AGEMA_signal_241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_75 ( .C ( clk ), .D ( new_AGEMA_signal_216 ), .Q ( new_AGEMA_signal_245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_103 ( .C ( clk ), .D ( N9 ), .Q ( new_AGEMA_signal_273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_111 ( .C ( clk ), .D ( new_AGEMA_signal_91 ), .Q ( new_AGEMA_signal_281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_119 ( .C ( clk ), .D ( new_AGEMA_signal_92 ), .Q ( new_AGEMA_signal_289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_127 ( .C ( clk ), .D ( new_AGEMA_signal_93 ), .Q ( new_AGEMA_signal_297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_135 ( .C ( clk ), .D ( N12 ), .Q ( new_AGEMA_signal_305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C ( clk ), .D ( new_AGEMA_signal_64 ), .Q ( new_AGEMA_signal_313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C ( clk ), .D ( new_AGEMA_signal_65 ), .Q ( new_AGEMA_signal_321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C ( clk ), .D ( new_AGEMA_signal_66 ), .Q ( new_AGEMA_signal_329 ) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U56 ( .s ({new_AGEMA_signal_216, new_AGEMA_signal_214, new_AGEMA_signal_212, new_AGEMA_signal_210}), .b ({new_AGEMA_signal_87, new_AGEMA_signal_86, new_AGEMA_signal_85, n42}), .a ({new_AGEMA_signal_224, new_AGEMA_signal_222, new_AGEMA_signal_220, new_AGEMA_signal_218}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, N19}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U58 ( .a ({new_AGEMA_signal_57, new_AGEMA_signal_56, new_AGEMA_signal_55, n43}), .b ({new_AGEMA_signal_224, new_AGEMA_signal_222, new_AGEMA_signal_220, new_AGEMA_signal_218}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, n47}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(1)) U62 ( .a ({new_AGEMA_signal_200, new_AGEMA_signal_198, new_AGEMA_signal_196, new_AGEMA_signal_194}), .b ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, n48}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, n44}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U65 ( .a ({new_AGEMA_signal_200, new_AGEMA_signal_198, new_AGEMA_signal_196, new_AGEMA_signal_194}), .b ({new_AGEMA_signal_63, new_AGEMA_signal_62, new_AGEMA_signal_61, n48}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_81, new_AGEMA_signal_80, new_AGEMA_signal_79, n49}) ) ;
    buf_clk new_AGEMA_reg_buffer_56 ( .C ( clk ), .D ( new_AGEMA_signal_225 ), .Q ( new_AGEMA_signal_226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_58 ( .C ( clk ), .D ( new_AGEMA_signal_227 ), .Q ( new_AGEMA_signal_228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_60 ( .C ( clk ), .D ( new_AGEMA_signal_229 ), .Q ( new_AGEMA_signal_230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_62 ( .C ( clk ), .D ( new_AGEMA_signal_231 ), .Q ( new_AGEMA_signal_232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_64 ( .C ( clk ), .D ( new_AGEMA_signal_233 ), .Q ( new_AGEMA_signal_234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_68 ( .C ( clk ), .D ( new_AGEMA_signal_237 ), .Q ( new_AGEMA_signal_238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_72 ( .C ( clk ), .D ( new_AGEMA_signal_241 ), .Q ( new_AGEMA_signal_242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_76 ( .C ( clk ), .D ( new_AGEMA_signal_245 ), .Q ( new_AGEMA_signal_246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_104 ( .C ( clk ), .D ( new_AGEMA_signal_273 ), .Q ( new_AGEMA_signal_274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_112 ( .C ( clk ), .D ( new_AGEMA_signal_281 ), .Q ( new_AGEMA_signal_282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_120 ( .C ( clk ), .D ( new_AGEMA_signal_289 ), .Q ( new_AGEMA_signal_290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_128 ( .C ( clk ), .D ( new_AGEMA_signal_297 ), .Q ( new_AGEMA_signal_298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_136 ( .C ( clk ), .D ( new_AGEMA_signal_305 ), .Q ( new_AGEMA_signal_306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C ( clk ), .D ( new_AGEMA_signal_313 ), .Q ( new_AGEMA_signal_314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_152 ( .C ( clk ), .D ( new_AGEMA_signal_321 ), .Q ( new_AGEMA_signal_322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_160 ( .C ( clk ), .D ( new_AGEMA_signal_329 ), .Q ( new_AGEMA_signal_330 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_65 ( .C ( clk ), .D ( new_AGEMA_signal_234 ), .Q ( new_AGEMA_signal_235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_69 ( .C ( clk ), .D ( new_AGEMA_signal_238 ), .Q ( new_AGEMA_signal_239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_73 ( .C ( clk ), .D ( new_AGEMA_signal_242 ), .Q ( new_AGEMA_signal_243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_77 ( .C ( clk ), .D ( new_AGEMA_signal_246 ), .Q ( new_AGEMA_signal_247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_79 ( .C ( clk ), .D ( n47 ), .Q ( new_AGEMA_signal_249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_81 ( .C ( clk ), .D ( new_AGEMA_signal_70 ), .Q ( new_AGEMA_signal_251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_83 ( .C ( clk ), .D ( new_AGEMA_signal_71 ), .Q ( new_AGEMA_signal_253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_85 ( .C ( clk ), .D ( new_AGEMA_signal_72 ), .Q ( new_AGEMA_signal_255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_87 ( .C ( clk ), .D ( n49 ), .Q ( new_AGEMA_signal_257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_91 ( .C ( clk ), .D ( new_AGEMA_signal_79 ), .Q ( new_AGEMA_signal_261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_95 ( .C ( clk ), .D ( new_AGEMA_signal_80 ), .Q ( new_AGEMA_signal_265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_99 ( .C ( clk ), .D ( new_AGEMA_signal_81 ), .Q ( new_AGEMA_signal_269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_105 ( .C ( clk ), .D ( new_AGEMA_signal_274 ), .Q ( new_AGEMA_signal_275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_113 ( .C ( clk ), .D ( new_AGEMA_signal_282 ), .Q ( new_AGEMA_signal_283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_121 ( .C ( clk ), .D ( new_AGEMA_signal_290 ), .Q ( new_AGEMA_signal_291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_129 ( .C ( clk ), .D ( new_AGEMA_signal_298 ), .Q ( new_AGEMA_signal_299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C ( clk ), .D ( new_AGEMA_signal_306 ), .Q ( new_AGEMA_signal_307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C ( clk ), .D ( new_AGEMA_signal_314 ), .Q ( new_AGEMA_signal_315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C ( clk ), .D ( new_AGEMA_signal_322 ), .Q ( new_AGEMA_signal_323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C ( clk ), .D ( new_AGEMA_signal_330 ), .Q ( new_AGEMA_signal_331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C ( clk ), .D ( N19 ), .Q ( new_AGEMA_signal_337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C ( clk ), .D ( new_AGEMA_signal_94 ), .Q ( new_AGEMA_signal_343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C ( clk ), .D ( new_AGEMA_signal_95 ), .Q ( new_AGEMA_signal_349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C ( clk ), .D ( new_AGEMA_signal_96 ), .Q ( new_AGEMA_signal_355 ) ) ;

    /* cells in depth 6 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U63 ( .a ({new_AGEMA_signal_232, new_AGEMA_signal_230, new_AGEMA_signal_228, new_AGEMA_signal_226}), .b ({new_AGEMA_signal_78, new_AGEMA_signal_77, new_AGEMA_signal_76, n44}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_90, new_AGEMA_signal_89, new_AGEMA_signal_88, n46}) ) ;
    buf_clk new_AGEMA_reg_buffer_66 ( .C ( clk ), .D ( new_AGEMA_signal_235 ), .Q ( new_AGEMA_signal_236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_70 ( .C ( clk ), .D ( new_AGEMA_signal_239 ), .Q ( new_AGEMA_signal_240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_74 ( .C ( clk ), .D ( new_AGEMA_signal_243 ), .Q ( new_AGEMA_signal_244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_78 ( .C ( clk ), .D ( new_AGEMA_signal_247 ), .Q ( new_AGEMA_signal_248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_80 ( .C ( clk ), .D ( new_AGEMA_signal_249 ), .Q ( new_AGEMA_signal_250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_82 ( .C ( clk ), .D ( new_AGEMA_signal_251 ), .Q ( new_AGEMA_signal_252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_84 ( .C ( clk ), .D ( new_AGEMA_signal_253 ), .Q ( new_AGEMA_signal_254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_86 ( .C ( clk ), .D ( new_AGEMA_signal_255 ), .Q ( new_AGEMA_signal_256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_88 ( .C ( clk ), .D ( new_AGEMA_signal_257 ), .Q ( new_AGEMA_signal_258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_92 ( .C ( clk ), .D ( new_AGEMA_signal_261 ), .Q ( new_AGEMA_signal_262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_96 ( .C ( clk ), .D ( new_AGEMA_signal_265 ), .Q ( new_AGEMA_signal_266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_100 ( .C ( clk ), .D ( new_AGEMA_signal_269 ), .Q ( new_AGEMA_signal_270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_106 ( .C ( clk ), .D ( new_AGEMA_signal_275 ), .Q ( new_AGEMA_signal_276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_114 ( .C ( clk ), .D ( new_AGEMA_signal_283 ), .Q ( new_AGEMA_signal_284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_122 ( .C ( clk ), .D ( new_AGEMA_signal_291 ), .Q ( new_AGEMA_signal_292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_130 ( .C ( clk ), .D ( new_AGEMA_signal_299 ), .Q ( new_AGEMA_signal_300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C ( clk ), .D ( new_AGEMA_signal_307 ), .Q ( new_AGEMA_signal_308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C ( clk ), .D ( new_AGEMA_signal_315 ), .Q ( new_AGEMA_signal_316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C ( clk ), .D ( new_AGEMA_signal_323 ), .Q ( new_AGEMA_signal_324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C ( clk ), .D ( new_AGEMA_signal_331 ), .Q ( new_AGEMA_signal_332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_168 ( .C ( clk ), .D ( new_AGEMA_signal_337 ), .Q ( new_AGEMA_signal_338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C ( clk ), .D ( new_AGEMA_signal_343 ), .Q ( new_AGEMA_signal_344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C ( clk ), .D ( new_AGEMA_signal_349 ), .Q ( new_AGEMA_signal_350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C ( clk ), .D ( new_AGEMA_signal_355 ), .Q ( new_AGEMA_signal_356 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_89 ( .C ( clk ), .D ( new_AGEMA_signal_258 ), .Q ( new_AGEMA_signal_259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_93 ( .C ( clk ), .D ( new_AGEMA_signal_262 ), .Q ( new_AGEMA_signal_263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_97 ( .C ( clk ), .D ( new_AGEMA_signal_266 ), .Q ( new_AGEMA_signal_267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_101 ( .C ( clk ), .D ( new_AGEMA_signal_270 ), .Q ( new_AGEMA_signal_271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_107 ( .C ( clk ), .D ( new_AGEMA_signal_276 ), .Q ( new_AGEMA_signal_277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_115 ( .C ( clk ), .D ( new_AGEMA_signal_284 ), .Q ( new_AGEMA_signal_285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_123 ( .C ( clk ), .D ( new_AGEMA_signal_292 ), .Q ( new_AGEMA_signal_293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_131 ( .C ( clk ), .D ( new_AGEMA_signal_300 ), .Q ( new_AGEMA_signal_301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C ( clk ), .D ( new_AGEMA_signal_308 ), .Q ( new_AGEMA_signal_309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C ( clk ), .D ( new_AGEMA_signal_316 ), .Q ( new_AGEMA_signal_317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C ( clk ), .D ( new_AGEMA_signal_324 ), .Q ( new_AGEMA_signal_325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C ( clk ), .D ( new_AGEMA_signal_332 ), .Q ( new_AGEMA_signal_333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C ( clk ), .D ( new_AGEMA_signal_338 ), .Q ( new_AGEMA_signal_339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C ( clk ), .D ( new_AGEMA_signal_344 ), .Q ( new_AGEMA_signal_345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C ( clk ), .D ( new_AGEMA_signal_350 ), .Q ( new_AGEMA_signal_351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C ( clk ), .D ( new_AGEMA_signal_356 ), .Q ( new_AGEMA_signal_357 ) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U64 ( .s ({new_AGEMA_signal_248, new_AGEMA_signal_244, new_AGEMA_signal_240, new_AGEMA_signal_236}), .b ({new_AGEMA_signal_256, new_AGEMA_signal_254, new_AGEMA_signal_252, new_AGEMA_signal_250}), .a ({new_AGEMA_signal_90, new_AGEMA_signal_89, new_AGEMA_signal_88, n46}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, n50}) ) ;
    buf_clk new_AGEMA_reg_buffer_90 ( .C ( clk ), .D ( new_AGEMA_signal_259 ), .Q ( new_AGEMA_signal_260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_94 ( .C ( clk ), .D ( new_AGEMA_signal_263 ), .Q ( new_AGEMA_signal_264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_98 ( .C ( clk ), .D ( new_AGEMA_signal_267 ), .Q ( new_AGEMA_signal_268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_102 ( .C ( clk ), .D ( new_AGEMA_signal_271 ), .Q ( new_AGEMA_signal_272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_108 ( .C ( clk ), .D ( new_AGEMA_signal_277 ), .Q ( new_AGEMA_signal_278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_116 ( .C ( clk ), .D ( new_AGEMA_signal_285 ), .Q ( new_AGEMA_signal_286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_124 ( .C ( clk ), .D ( new_AGEMA_signal_293 ), .Q ( new_AGEMA_signal_294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_132 ( .C ( clk ), .D ( new_AGEMA_signal_301 ), .Q ( new_AGEMA_signal_302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C ( clk ), .D ( new_AGEMA_signal_309 ), .Q ( new_AGEMA_signal_310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C ( clk ), .D ( new_AGEMA_signal_317 ), .Q ( new_AGEMA_signal_318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C ( clk ), .D ( new_AGEMA_signal_325 ), .Q ( new_AGEMA_signal_326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C ( clk ), .D ( new_AGEMA_signal_333 ), .Q ( new_AGEMA_signal_334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C ( clk ), .D ( new_AGEMA_signal_339 ), .Q ( new_AGEMA_signal_340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C ( clk ), .D ( new_AGEMA_signal_345 ), .Q ( new_AGEMA_signal_346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C ( clk ), .D ( new_AGEMA_signal_351 ), .Q ( new_AGEMA_signal_352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C ( clk ), .D ( new_AGEMA_signal_357 ), .Q ( new_AGEMA_signal_358 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_109 ( .C ( clk ), .D ( new_AGEMA_signal_278 ), .Q ( new_AGEMA_signal_279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_117 ( .C ( clk ), .D ( new_AGEMA_signal_286 ), .Q ( new_AGEMA_signal_287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_125 ( .C ( clk ), .D ( new_AGEMA_signal_294 ), .Q ( new_AGEMA_signal_295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_133 ( .C ( clk ), .D ( new_AGEMA_signal_302 ), .Q ( new_AGEMA_signal_303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C ( clk ), .D ( new_AGEMA_signal_310 ), .Q ( new_AGEMA_signal_311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C ( clk ), .D ( new_AGEMA_signal_318 ), .Q ( new_AGEMA_signal_319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C ( clk ), .D ( new_AGEMA_signal_326 ), .Q ( new_AGEMA_signal_327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C ( clk ), .D ( new_AGEMA_signal_334 ), .Q ( new_AGEMA_signal_335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C ( clk ), .D ( new_AGEMA_signal_340 ), .Q ( new_AGEMA_signal_341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C ( clk ), .D ( new_AGEMA_signal_346 ), .Q ( new_AGEMA_signal_347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C ( clk ), .D ( new_AGEMA_signal_352 ), .Q ( new_AGEMA_signal_353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C ( clk ), .D ( new_AGEMA_signal_358 ), .Q ( new_AGEMA_signal_359 ) ) ;

    /* cells in depth 10 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U66 ( .a ({new_AGEMA_signal_99, new_AGEMA_signal_98, new_AGEMA_signal_97, n50}), .b ({new_AGEMA_signal_272, new_AGEMA_signal_268, new_AGEMA_signal_264, new_AGEMA_signal_260}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_102, new_AGEMA_signal_101, new_AGEMA_signal_100, N27}) ) ;
    buf_clk new_AGEMA_reg_buffer_110 ( .C ( clk ), .D ( new_AGEMA_signal_279 ), .Q ( new_AGEMA_signal_280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_118 ( .C ( clk ), .D ( new_AGEMA_signal_287 ), .Q ( new_AGEMA_signal_288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_126 ( .C ( clk ), .D ( new_AGEMA_signal_295 ), .Q ( new_AGEMA_signal_296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_134 ( .C ( clk ), .D ( new_AGEMA_signal_303 ), .Q ( new_AGEMA_signal_304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C ( clk ), .D ( new_AGEMA_signal_311 ), .Q ( new_AGEMA_signal_312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C ( clk ), .D ( new_AGEMA_signal_319 ), .Q ( new_AGEMA_signal_320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C ( clk ), .D ( new_AGEMA_signal_327 ), .Q ( new_AGEMA_signal_328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C ( clk ), .D ( new_AGEMA_signal_335 ), .Q ( new_AGEMA_signal_336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C ( clk ), .D ( new_AGEMA_signal_341 ), .Q ( new_AGEMA_signal_342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C ( clk ), .D ( new_AGEMA_signal_347 ), .Q ( new_AGEMA_signal_348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C ( clk ), .D ( new_AGEMA_signal_353 ), .Q ( new_AGEMA_signal_354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C ( clk ), .D ( new_AGEMA_signal_359 ), .Q ( new_AGEMA_signal_360 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_304, new_AGEMA_signal_296, new_AGEMA_signal_288, new_AGEMA_signal_280}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_336, new_AGEMA_signal_328, new_AGEMA_signal_320, new_AGEMA_signal_312}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_360, new_AGEMA_signal_354, new_AGEMA_signal_348, new_AGEMA_signal_342}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_102, new_AGEMA_signal_101, new_AGEMA_signal_100, N27}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
