module Reg1(x, y);
 input [158:0] x;
 output [157:0] y;

  register_stage #(.WIDTH(158)) inst_0(.clk(x[0]), .D({x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[95],x[96],x[97],x[98],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[15],x[16],x[17],x[18],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157]}));
endmodule

module Reg2(x, y);
 input [250:0] x;
 output [249:0] y;

  register_stage #(.WIDTH(250)) inst_0(.clk(x[0]), .D({x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[171],x[172],x[173],x[174],x[175],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[71],x[72],x[73],x[74],x[75],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[205],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [365:0] x;
 output [207:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx29 Fx29_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx30 Fx30_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx34 Fx34_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx35 Fx35_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx39 Fx39_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx40 Fx40_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx44 Fx44_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx45 Fx45_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx49 Fx49_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx50 Fx50_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx54 Fx54_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx55 Fx55_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx59 Fx59_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx60 Fx60_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx64 Fx64_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx65 Fx65_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx69 Fx69_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx70 Fx70_inst(.x({x[46], x[45], x[44], x[43], x[42]}), .y(y[28]));
  Fx71 Fx71_inst(.x({x[47], x[45]}), .y(y[29]));
  Fx72 Fx72_inst(.x({x[48], x[44]}), .y(y[30]));
  Fx73 Fx73_inst(.x({x[49], x[43]}), .y(y[31]));
  Fx74 Fx74_inst(.x({x[50], x[42]}), .y(y[32]));
  Fx75 Fx75_inst(.x({x[55], x[54], x[53], x[52], x[51]}), .y(y[33]));
  Fx76 Fx76_inst(.x({x[56], x[54]}), .y(y[34]));
  Fx77 Fx77_inst(.x({x[57], x[53]}), .y(y[35]));
  Fx78 Fx78_inst(.x({x[58], x[52]}), .y(y[36]));
  Fx79 Fx79_inst(.x({x[59], x[51]}), .y(y[37]));
  Fx80 Fx80_inst(.x({x[64], x[63], x[62], x[61], x[60]}), .y(y[38]));
  Fx81 Fx81_inst(.x({x[65], x[63]}), .y(y[39]));
  Fx82 Fx82_inst(.x({x[66], x[62]}), .y(y[40]));
  Fx83 Fx83_inst(.x({x[67], x[61]}), .y(y[41]));
  Fx84 Fx84_inst(.x({x[68], x[60]}), .y(y[42]));
  Fx85 Fx85_inst(.x({x[73], x[72], x[71], x[70], x[69]}), .y(y[43]));
  Fx86 Fx86_inst(.x({x[74], x[72]}), .y(y[44]));
  Fx87 Fx87_inst(.x({x[75], x[71]}), .y(y[45]));
  Fx88 Fx88_inst(.x({x[76], x[70]}), .y(y[46]));
  Fx89 Fx89_inst(.x({x[77], x[69]}), .y(y[47]));
  Fx90 Fx90_inst(.x({x[82], x[81], x[80], x[79], x[78]}), .y(y[48]));
  Fx91 Fx91_inst(.x({x[83], x[81]}), .y(y[49]));
  Fx92 Fx92_inst(.x({x[84], x[80]}), .y(y[50]));
  Fx93 Fx93_inst(.x({x[85], x[79]}), .y(y[51]));
  Fx94 Fx94_inst(.x({x[86], x[78]}), .y(y[52]));
  Fx95 Fx95_inst(.x({x[91], x[90], x[89], x[88], x[87]}), .y(y[53]));
  Fx96 Fx96_inst(.x({x[92], x[90]}), .y(y[54]));
  Fx97 Fx97_inst(.x({x[93], x[89]}), .y(y[55]));
  Fx98 Fx98_inst(.x({x[94], x[88]}), .y(y[56]));
  Fx99 Fx99_inst(.x({x[95], x[87]}), .y(y[57]));
  Fx100 Fx100_inst(.x({x[100], x[99], x[98], x[97], x[96]}), .y(y[58]));
  Fx101 Fx101_inst(.x({x[101], x[99]}), .y(y[59]));
  Fx102 Fx102_inst(.x({x[102], x[98]}), .y(y[60]));
  Fx103 Fx103_inst(.x({x[103], x[97]}), .y(y[61]));
  Fx104 Fx104_inst(.x({x[104], x[96]}), .y(y[62]));
  Fx105 Fx105_inst(.x({x[109], x[108], x[107], x[106], x[105]}), .y(y[63]));
  Fx106 Fx106_inst(.x({x[110], x[108]}), .y(y[64]));
  Fx107 Fx107_inst(.x({x[111], x[107]}), .y(y[65]));
  Fx108 Fx108_inst(.x({x[112], x[106]}), .y(y[66]));
  Fx109 Fx109_inst(.x({x[113], x[105]}), .y(y[67]));
  Fx110 Fx110_inst(.x({x[118], x[117], x[116], x[115], x[114]}), .y(y[68]));
  Fx111 Fx111_inst(.x({x[119], x[117]}), .y(y[69]));
  Fx112 Fx112_inst(.x({x[120], x[116]}), .y(y[70]));
  Fx113 Fx113_inst(.x({x[121], x[115]}), .y(y[71]));
  Fx114 Fx114_inst(.x({x[122], x[114]}), .y(y[72]));
  Fx115 Fx115_inst(.x({x[127], x[126], x[125], x[124], x[123]}), .y(y[73]));
  Fx116 Fx116_inst(.x({x[128], x[126]}), .y(y[74]));
  Fx117 Fx117_inst(.x({x[129], x[125]}), .y(y[75]));
  Fx118 Fx118_inst(.x({x[130], x[124]}), .y(y[76]));
  Fx119 Fx119_inst(.x({x[131], x[123]}), .y(y[77]));
  Fx120 Fx120_inst(.x({x[136], x[135], x[134], x[133], x[132]}), .y(y[78]));
  Fx121 Fx121_inst(.x({x[137], x[135]}), .y(y[79]));
  Fx122 Fx122_inst(.x({x[138], x[134]}), .y(y[80]));
  Fx123 Fx123_inst(.x({x[139], x[133]}), .y(y[81]));
  Fx124 Fx124_inst(.x({x[140], x[132]}), .y(y[82]));
  Fx125 Fx125_inst(.x({x[145], x[144], x[143], x[142], x[141]}), .y(y[83]));
  Fx126 Fx126_inst(.x({x[146], x[144]}), .y(y[84]));
  Fx127 Fx127_inst(.x({x[147], x[143]}), .y(y[85]));
  Fx128 Fx128_inst(.x({x[148], x[142]}), .y(y[86]));
  Fx129 Fx129_inst(.x({x[149], x[141]}), .y(y[87]));
  Fx130 Fx130_inst(.x({x[154], x[153], x[152], x[151], x[150]}), .y(y[88]));
  Fx131 Fx131_inst(.x({x[155], x[153]}), .y(y[89]));
  Fx132 Fx132_inst(.x({x[156], x[152]}), .y(y[90]));
  Fx133 Fx133_inst(.x({x[157], x[151]}), .y(y[91]));
  Fx134 Fx134_inst(.x({x[158], x[150]}), .y(y[92]));
  Fx135 Fx135_inst(.x({x[163], x[162], x[161], x[160], x[159]}), .y(y[93]));
  Fx136 Fx136_inst(.x({x[164], x[162]}), .y(y[94]));
  Fx137 Fx137_inst(.x({x[165], x[161]}), .y(y[95]));
  Fx138 Fx138_inst(.x({x[166], x[160]}), .y(y[96]));
  Fx139 Fx139_inst(.x({x[167], x[159]}), .y(y[97]));
  Fx140 Fx140_inst(.x({x[172], x[171], x[170], x[169], x[168]}), .y(y[98]));
  Fx141 Fx141_inst(.x({x[173], x[171]}), .y(y[99]));
  Fx142 Fx142_inst(.x({x[174], x[170]}), .y(y[100]));
  Fx143 Fx143_inst(.x({x[175], x[169]}), .y(y[101]));
  Fx144 Fx144_inst(.x({x[176], x[168]}), .y(y[102]));
  Fx145 Fx145_inst(.x({x[181], x[180], x[179], x[178], x[177]}), .y(y[103]));
  Fx146 Fx146_inst(.x({x[182], x[180]}), .y(y[104]));
  Fx147 Fx147_inst(.x({x[183], x[179]}), .y(y[105]));
  Fx148 Fx148_inst(.x({x[184], x[178]}), .y(y[106]));
  Fx149 Fx149_inst(.x({x[185], x[177]}), .y(y[107]));
  Fx150 Fx150_inst(.x({x[190], x[189], x[188], x[187], x[186]}), .y(y[108]));
  Fx151 Fx151_inst(.x({x[191], x[189]}), .y(y[109]));
  Fx152 Fx152_inst(.x({x[192], x[188]}), .y(y[110]));
  Fx153 Fx153_inst(.x({x[193], x[187]}), .y(y[111]));
  Fx154 Fx154_inst(.x({x[194], x[186]}), .y(y[112]));
  Fx155 Fx155_inst(.x({x[199], x[198], x[197], x[196], x[195]}), .y(y[113]));
  Fx156 Fx156_inst(.x({x[200], x[198]}), .y(y[114]));
  Fx157 Fx157_inst(.x({x[201], x[197]}), .y(y[115]));
  Fx158 Fx158_inst(.x({x[202], x[196]}), .y(y[116]));
  Fx159 Fx159_inst(.x({x[203], x[195]}), .y(y[117]));
  Fx160 Fx160_inst(.x({x[208], x[207], x[206], x[205], x[204]}), .y(y[118]));
  Fx161 Fx161_inst(.x({x[209], x[207]}), .y(y[119]));
  Fx162 Fx162_inst(.x({x[210], x[206]}), .y(y[120]));
  Fx163 Fx163_inst(.x({x[211], x[205]}), .y(y[121]));
  Fx164 Fx164_inst(.x({x[212], x[204]}), .y(y[122]));
  Fx165 Fx165_inst(.x({x[217], x[216], x[215], x[214], x[213]}), .y(y[123]));
  Fx166 Fx166_inst(.x({x[218], x[216]}), .y(y[124]));
  Fx167 Fx167_inst(.x({x[219], x[215]}), .y(y[125]));
  Fx168 Fx168_inst(.x({x[220], x[214]}), .y(y[126]));
  Fx169 Fx169_inst(.x({x[221], x[213]}), .y(y[127]));
  Fx170 Fx170_inst(.x({x[226], x[225], x[224], x[223], x[222]}), .y(y[128]));
  Fx171 Fx171_inst(.x({x[227], x[225]}), .y(y[129]));
  Fx172 Fx172_inst(.x({x[228], x[224]}), .y(y[130]));
  Fx173 Fx173_inst(.x({x[229], x[223]}), .y(y[131]));
  Fx174 Fx174_inst(.x({x[230], x[222]}), .y(y[132]));
  Fx175 Fx175_inst(.x({x[235], x[234], x[233], x[232], x[231]}), .y(y[133]));
  Fx176 Fx176_inst(.x({x[236], x[234]}), .y(y[134]));
  Fx177 Fx177_inst(.x({x[237], x[233]}), .y(y[135]));
  Fx178 Fx178_inst(.x({x[238], x[232]}), .y(y[136]));
  Fx179 Fx179_inst(.x({x[239], x[231]}), .y(y[137]));
  Fx180 Fx180_inst(.x({x[244], x[243], x[242], x[241], x[240]}), .y(y[138]));
  Fx181 Fx181_inst(.x({x[245], x[243]}), .y(y[139]));
  Fx182 Fx182_inst(.x({x[246], x[242]}), .y(y[140]));
  Fx183 Fx183_inst(.x({x[247], x[241]}), .y(y[141]));
  Fx184 Fx184_inst(.x({x[248], x[240]}), .y(y[142]));
  Fx185 Fx185_inst(.x({x[253], x[252], x[251], x[250], x[249]}), .y(y[143]));
  Fx186 Fx186_inst(.x({x[254], x[252]}), .y(y[144]));
  Fx187 Fx187_inst(.x({x[255], x[251]}), .y(y[145]));
  Fx188 Fx188_inst(.x({x[256], x[250]}), .y(y[146]));
  Fx189 Fx189_inst(.x({x[257], x[249]}), .y(y[147]));
  Fx190 Fx190_inst(.x({x[262], x[261], x[260], x[259], x[258]}), .y(y[148]));
  Fx191 Fx191_inst(.x({x[263], x[261]}), .y(y[149]));
  Fx192 Fx192_inst(.x({x[264], x[260]}), .y(y[150]));
  Fx193 Fx193_inst(.x({x[265], x[259]}), .y(y[151]));
  Fx194 Fx194_inst(.x({x[266], x[258]}), .y(y[152]));
  Fx195 Fx195_inst(.x({x[271], x[270], x[269], x[268], x[267]}), .y(y[153]));
  Fx196 Fx196_inst(.x({x[272], x[270]}), .y(y[154]));
  Fx197 Fx197_inst(.x({x[273], x[269]}), .y(y[155]));
  Fx198 Fx198_inst(.x({x[274], x[268]}), .y(y[156]));
  Fx199 Fx199_inst(.x({x[275], x[267]}), .y(y[157]));
  Fx200 Fx200_inst(.x({x[280], x[279], x[278], x[277], x[276]}), .y(y[158]));
  Fx201 Fx201_inst(.x({x[281], x[279]}), .y(y[159]));
  Fx202 Fx202_inst(.x({x[282], x[278]}), .y(y[160]));
  Fx203 Fx203_inst(.x({x[283], x[277]}), .y(y[161]));
  Fx204 Fx204_inst(.x({x[284], x[276]}), .y(y[162]));
  Fx205 Fx205_inst(.x({x[289], x[288], x[287], x[286], x[285]}), .y(y[163]));
  Fx206 Fx206_inst(.x({x[290], x[288]}), .y(y[164]));
  Fx207 Fx207_inst(.x({x[291], x[287]}), .y(y[165]));
  Fx208 Fx208_inst(.x({x[292], x[286]}), .y(y[166]));
  Fx209 Fx209_inst(.x({x[293], x[285]}), .y(y[167]));
  Fx210 Fx210_inst(.x({x[298], x[297], x[296], x[295], x[294]}), .y(y[168]));
  Fx211 Fx211_inst(.x({x[299], x[297]}), .y(y[169]));
  Fx212 Fx212_inst(.x({x[300], x[296]}), .y(y[170]));
  Fx213 Fx213_inst(.x({x[301], x[295]}), .y(y[171]));
  Fx214 Fx214_inst(.x({x[302], x[294]}), .y(y[172]));
  Fx215 Fx215_inst(.x({x[307], x[306], x[305], x[304], x[303]}), .y(y[173]));
  Fx216 Fx216_inst(.x({x[308], x[306]}), .y(y[174]));
  Fx217 Fx217_inst(.x({x[309], x[305]}), .y(y[175]));
  Fx218 Fx218_inst(.x({x[310], x[304]}), .y(y[176]));
  Fx219 Fx219_inst(.x({x[311], x[303]}), .y(y[177]));
  Fx220 Fx220_inst(.x({x[316], x[315], x[314], x[313], x[312]}), .y(y[178]));
  Fx221 Fx221_inst(.x({x[317], x[315]}), .y(y[179]));
  Fx222 Fx222_inst(.x({x[318], x[314]}), .y(y[180]));
  Fx223 Fx223_inst(.x({x[319], x[313]}), .y(y[181]));
  Fx224 Fx224_inst(.x({x[320], x[312]}), .y(y[182]));
  Fx225 Fx225_inst(.x({x[325], x[324], x[323], x[322], x[321]}), .y(y[183]));
  Fx226 Fx226_inst(.x({x[326], x[324]}), .y(y[184]));
  Fx227 Fx227_inst(.x({x[327], x[323]}), .y(y[185]));
  Fx228 Fx228_inst(.x({x[328], x[322]}), .y(y[186]));
  Fx229 Fx229_inst(.x({x[329], x[321]}), .y(y[187]));
  Fx230 Fx230_inst(.x({x[334], x[333], x[332], x[331], x[330]}), .y(y[188]));
  Fx231 Fx231_inst(.x({x[335], x[333]}), .y(y[189]));
  Fx232 Fx232_inst(.x({x[336], x[332]}), .y(y[190]));
  Fx233 Fx233_inst(.x({x[337], x[331]}), .y(y[191]));
  Fx234 Fx234_inst(.x({x[338], x[330]}), .y(y[192]));
  Fx235 Fx235_inst(.x({x[343], x[342], x[341], x[340], x[339]}), .y(y[193]));
  Fx236 Fx236_inst(.x({x[344], x[342]}), .y(y[194]));
  Fx237 Fx237_inst(.x({x[345], x[341]}), .y(y[195]));
  Fx238 Fx238_inst(.x({x[346], x[340]}), .y(y[196]));
  Fx239 Fx239_inst(.x({x[347], x[339]}), .y(y[197]));
  Fx240 Fx240_inst(.x({x[352], x[351], x[350], x[349], x[348]}), .y(y[198]));
  Fx241 Fx241_inst(.x({x[353], x[351]}), .y(y[199]));
  Fx242 Fx242_inst(.x({x[354], x[350]}), .y(y[200]));
  Fx243 Fx243_inst(.x({x[355], x[349]}), .y(y[201]));
  Fx244 Fx244_inst(.x({x[356], x[348]}), .y(y[202]));
  Fx245 Fx245_inst(.x({x[361], x[360], x[359], x[358], x[357]}), .y(y[203]));
  Fx246 Fx246_inst(.x({x[362], x[360]}), .y(y[204]));
  Fx247 Fx247_inst(.x({x[363], x[359]}), .y(y[205]));
  Fx248 Fx248_inst(.x({x[364], x[358]}), .y(y[206]));
  Fx249 Fx249_inst(.x({x[365], x[357]}), .y(y[207]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [23:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[16] | t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = ~(t[15]);
  assign t[13] = t[21] ^ x[2];
  assign t[14] = t[22] ^ x[5];
  assign t[15] = t[23] ^ x[8];
  assign t[16] = t[24] ^ x[11];
  assign t[17] = t[25] ^ x[14];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[20];
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = t[28] ^ x[23];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[3] & x[4]);
  assign t[23] = (x[6] & x[7]);
  assign t[24] = (x[9] & x[10]);
  assign t[25] = (x[12] & x[13]);
  assign t[26] = (x[15] & x[16]);
  assign t[27] = (x[18] & x[19]);
  assign t[28] = (x[21] & x[22]);
  assign t[2] = ~(t[13] | t[14]);
  assign t[3] = ~(t[6] | t[15]);
  assign t[4] = ~(t[13] | t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[16]);
  assign t[7] = ~(t[14] & t[10]);
  assign t[8] = ~(t[17] & t[18]);
  assign t[9] = ~(t[19] & t[20]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind66(x, y);
 input [41:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] ^ t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[26]);
  assign t[1] = ~(t[5] & t[44]);
  assign t[20] = t[25] ? t[46] : t[27];
  assign t[21] = t[25] ? t[47] : t[28];
  assign t[22] = t[25] ? t[48] : t[29];
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[13]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = t[25] ? t[49] : t[34];
  assign t[27] = t[50] ^ t[51];
  assign t[28] = t[48] ^ t[52];
  assign t[29] = t[45] ^ t[53];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[54] | t[35]);
  assign t[31] = ~(t[36]);
  assign t[32] = ~(t[37] & t[38]);
  assign t[33] = ~(t[54] & t[39]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = ~(t[57] & t[40]);
  assign t[36] = ~(t[37] & t[41]);
  assign t[37] = ~(t[58]);
  assign t[38] = ~(t[57]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[45]);
  assign t[40] = ~(t[58] | t[42]);
  assign t[41] = t[43] & t[59];
  assign t[42] = ~(t[39]);
  assign t[43] = ~(t[54] | t[57]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[10];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[14];
  assign t[49] = t[65] ^ x[16];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[66] ^ x[18];
  assign t[51] = t[67] ^ x[21];
  assign t[52] = t[68] ^ x[23];
  assign t[53] = t[69] ^ x[25];
  assign t[54] = t[70] ^ x[28];
  assign t[55] = t[71] ^ x[30];
  assign t[56] = t[72] ^ x[32];
  assign t[57] = t[73] ^ x[35];
  assign t[58] = t[74] ^ x[38];
  assign t[59] = t[75] ^ x[41];
  assign t[5] = ~(t[7] | t[6]);
  assign t[60] = (x[0] & x[1]);
  assign t[61] = (x[3] & x[4]);
  assign t[62] = (x[8] & x[9]);
  assign t[63] = (x[8] & x[11]);
  assign t[64] = (x[3] & x[13]);
  assign t[65] = (x[8] & x[15]);
  assign t[66] = (x[3] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[19] & x[22]);
  assign t[69] = (x[19] & x[24]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[26] & x[27]);
  assign t[71] = (x[3] & x[29]);
  assign t[72] = (x[19] & x[31]);
  assign t[73] = (x[33] & x[34]);
  assign t[74] = (x[36] & x[37]);
  assign t[75] = (x[39] & x[40]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[7] : t[11];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind67(x, y);
 input [41:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[26] | t[21]);
  assign t[1] = ~(t[5] & t[51]);
  assign t[20] = t[27] ? t[29] : t[28];
  assign t[21] = ~(t[30]);
  assign t[22] = ~(t[27] ^ t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[13]);
  assign t[25] = ~(t[34] | t[35]);
  assign t[26] = ~(t[27] | t[31]);
  assign t[27] = t[25] ? t[53] : t[36];
  assign t[28] = t[25] ? t[54] : t[37];
  assign t[29] = ~(t[28] & t[38]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[25] ? t[55] : t[39];
  assign t[31] = t[25] ? t[56] : t[40];
  assign t[32] = ~(t[57] | t[41]);
  assign t[33] = ~(t[42]);
  assign t[34] = ~(t[43] & t[44]);
  assign t[35] = ~(t[57] & t[45]);
  assign t[36] = t[56] ^ t[58];
  assign t[37] = t[52] ^ t[59];
  assign t[38] = ~(t[46] & t[21]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[52]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] & t[47]);
  assign t[42] = ~(t[43] & t[48]);
  assign t[43] = ~(t[65]);
  assign t[44] = ~(t[64]);
  assign t[45] = ~(t[66]);
  assign t[46] = ~(t[31]);
  assign t[47] = ~(t[65] | t[49]);
  assign t[48] = t[50] & t[66];
  assign t[49] = ~(t[45]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = ~(t[57] | t[64]);
  assign t[51] = t[67] ^ x[2];
  assign t[52] = t[68] ^ x[5];
  assign t[53] = t[69] ^ x[10];
  assign t[54] = t[70] ^ x[12];
  assign t[55] = t[71] ^ x[14];
  assign t[56] = t[72] ^ x[16];
  assign t[57] = t[73] ^ x[19];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[24];
  assign t[5] = ~(t[7] | t[6]);
  assign t[60] = t[76] ^ x[26];
  assign t[61] = t[77] ^ x[28];
  assign t[62] = t[78] ^ x[30];
  assign t[63] = t[79] ^ x[32];
  assign t[64] = t[80] ^ x[35];
  assign t[65] = t[81] ^ x[38];
  assign t[66] = t[82] ^ x[41];
  assign t[67] = (x[0] & x[1]);
  assign t[68] = (x[3] & x[4]);
  assign t[69] = (x[8] & x[9]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[8] & x[11]);
  assign t[71] = (x[8] & x[13]);
  assign t[72] = (x[3] & x[15]);
  assign t[73] = (x[17] & x[18]);
  assign t[74] = (x[20] & x[21]);
  assign t[75] = (x[20] & x[23]);
  assign t[76] = (x[3] & x[25]);
  assign t[77] = (x[20] & x[27]);
  assign t[78] = (x[3] & x[29]);
  assign t[79] = (x[20] & x[31]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[33] & x[34]);
  assign t[81] = (x[36] & x[37]);
  assign t[82] = (x[39] & x[40]);
  assign t[8] = x[6] ? x[7] : t[11];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind68(x, y);
 input [41:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[5] & t[55]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = t[32] ? t[20] : t[28];
  assign t[23] = ~(t[33] | t[34]);
  assign t[24] = ~(t[13]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[26] = t[25] ? t[57] : t[37];
  assign t[27] = ~(t[38] | t[39]);
  assign t[28] = t[25] ? t[58] : t[40];
  assign t[29] = ~(t[41] & t[31]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[32] | t[42]);
  assign t[31] = ~(t[26]);
  assign t[32] = t[25] ? t[59] : t[43];
  assign t[33] = ~(t[60] | t[44]);
  assign t[34] = ~(t[45]);
  assign t[35] = ~(t[46] & t[47]);
  assign t[36] = ~(t[60] & t[48]);
  assign t[37] = t[56] ^ t[61];
  assign t[38] = ~(t[32]);
  assign t[39] = ~(t[41] & t[49]);
  assign t[3] = ~(t[56]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[42]);
  assign t[42] = t[25] ? t[64] : t[50];
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[51]);
  assign t[45] = ~(t[46] & t[52]);
  assign t[46] = ~(t[67]);
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[68]);
  assign t[49] = ~(t[28]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[69] ^ t[70];
  assign t[51] = ~(t[67] | t[53]);
  assign t[52] = t[54] & t[68];
  assign t[53] = ~(t[48]);
  assign t[54] = ~(t[60] | t[66]);
  assign t[55] = t[71] ^ x[2];
  assign t[56] = t[72] ^ x[5];
  assign t[57] = t[73] ^ x[10];
  assign t[58] = t[74] ^ x[12];
  assign t[59] = t[75] ^ x[14];
  assign t[5] = ~(t[7] | t[6]);
  assign t[60] = t[76] ^ x[17];
  assign t[61] = t[77] ^ x[20];
  assign t[62] = t[78] ^ x[22];
  assign t[63] = t[79] ^ x[24];
  assign t[64] = t[80] ^ x[26];
  assign t[65] = t[81] ^ x[28];
  assign t[66] = t[82] ^ x[31];
  assign t[67] = t[83] ^ x[34];
  assign t[68] = t[84] ^ x[37];
  assign t[69] = t[85] ^ x[39];
  assign t[6] = ~(t[9]);
  assign t[70] = t[86] ^ x[41];
  assign t[71] = (x[0] & x[1]);
  assign t[72] = (x[3] & x[4]);
  assign t[73] = (x[8] & x[9]);
  assign t[74] = (x[8] & x[11]);
  assign t[75] = (x[8] & x[13]);
  assign t[76] = (x[15] & x[16]);
  assign t[77] = (x[18] & x[19]);
  assign t[78] = (x[3] & x[21]);
  assign t[79] = (x[18] & x[23]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[3] & x[25]);
  assign t[81] = (x[18] & x[27]);
  assign t[82] = (x[29] & x[30]);
  assign t[83] = (x[32] & x[33]);
  assign t[84] = (x[35] & x[36]);
  assign t[85] = (x[3] & x[38]);
  assign t[86] = (x[18] & x[40]);
  assign t[8] = x[6] ? x[7] : t[11];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind69(x, y);
 input [41:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26]);
  assign t[18] = ~(x[6]);
  assign t[19] = t[26] ? t[53] : t[27];
  assign t[1] = ~(t[5] & t[51]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[22] = ~(t[19] | t[32]);
  assign t[23] = ~(t[28]);
  assign t[24] = ~(t[33] | t[34]);
  assign t[25] = ~(t[13]);
  assign t[26] = ~(t[35] | t[36]);
  assign t[27] = t[52] ^ t[54];
  assign t[28] = t[26] ? t[55] : t[37];
  assign t[29] = ~(t[38] & t[30]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[39]);
  assign t[31] = ~(t[38] & t[23]);
  assign t[32] = t[26] ? t[52] : t[40];
  assign t[33] = ~(t[56] | t[41]);
  assign t[34] = ~(t[42]);
  assign t[35] = ~(t[43] & t[44]);
  assign t[36] = ~(t[56] & t[45]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = ~(t[32]);
  assign t[39] = t[26] ? t[59] : t[46];
  assign t[3] = ~(t[52]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[62] & t[47]);
  assign t[42] = ~(t[43] & t[48]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[62]);
  assign t[45] = ~(t[64]);
  assign t[46] = t[65] ^ t[66];
  assign t[47] = ~(t[63] | t[49]);
  assign t[48] = t[50] & t[64];
  assign t[49] = ~(t[45]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = ~(t[56] | t[62]);
  assign t[51] = t[67] ^ x[2];
  assign t[52] = t[68] ^ x[5];
  assign t[53] = t[69] ^ x[10];
  assign t[54] = t[70] ^ x[13];
  assign t[55] = t[71] ^ x[15];
  assign t[56] = t[72] ^ x[18];
  assign t[57] = t[73] ^ x[20];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[24];
  assign t[5] = ~(t[7] | t[6]);
  assign t[60] = t[76] ^ x[26];
  assign t[61] = t[77] ^ x[28];
  assign t[62] = t[78] ^ x[31];
  assign t[63] = t[79] ^ x[34];
  assign t[64] = t[80] ^ x[37];
  assign t[65] = t[81] ^ x[39];
  assign t[66] = t[82] ^ x[41];
  assign t[67] = (x[0] & x[1]);
  assign t[68] = (x[3] & x[4]);
  assign t[69] = (x[8] & x[9]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[11] & x[12]);
  assign t[71] = (x[8] & x[14]);
  assign t[72] = (x[16] & x[17]);
  assign t[73] = (x[3] & x[19]);
  assign t[74] = (x[11] & x[21]);
  assign t[75] = (x[8] & x[23]);
  assign t[76] = (x[3] & x[25]);
  assign t[77] = (x[11] & x[27]);
  assign t[78] = (x[29] & x[30]);
  assign t[79] = (x[32] & x[33]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[35] & x[36]);
  assign t[81] = (x[3] & x[38]);
  assign t[82] = (x[11] & x[40]);
  assign t[8] = x[6] ? x[7] : t[11];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind70(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind71(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind72(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind73(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind74(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind75(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind76(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind77(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind78(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind79(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind80(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind81(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind82(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind83(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind84(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind85(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind86(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[9] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind87(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind88(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind89(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind90(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[9] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind91(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind92(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind93(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind94(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[9] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind95(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind96(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind97(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind98(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind99(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind100(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind101(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind102(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind103(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind104(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind105(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind106(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind107(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind108(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind109(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind110(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind111(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind112(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind113(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind114(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind115(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind116(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind117(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind118(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind119(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind120(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind121(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind122(x, y);
 input [21:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[33] & t[21]);
  assign t[17] = ~(t[22] | t[23]);
  assign t[18] = ~(t[7]);
  assign t[19] = ~(t[34]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[33] | t[24]);
  assign t[23] = ~(t[25]);
  assign t[24] = ~(t[35] & t[26]);
  assign t[25] = ~(t[19] & t[27]);
  assign t[26] = ~(t[34] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[33] | t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[8];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = t[42] ^ x[18];
  assign t[36] = t[43] ^ x[21];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[3] & x[7]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[10] & x[11]);
  assign t[41] = (x[13] & x[14]);
  assign t[42] = (x[16] & x[17]);
  assign t[43] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[9] : t[32];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind123(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[33] & t[21]);
  assign t[17] = ~(t[22] | t[23]);
  assign t[18] = ~(t[7]);
  assign t[19] = ~(t[34]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[33] | t[24]);
  assign t[23] = ~(t[25]);
  assign t[24] = ~(t[35] & t[26]);
  assign t[25] = ~(t[19] & t[27]);
  assign t[26] = ~(t[34] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[33] | t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind124(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[33] & t[21]);
  assign t[17] = ~(t[22] | t[23]);
  assign t[18] = ~(t[7]);
  assign t[19] = ~(t[34]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[33] | t[24]);
  assign t[23] = ~(t[25]);
  assign t[24] = ~(t[35] & t[26]);
  assign t[25] = ~(t[19] & t[27]);
  assign t[26] = ~(t[34] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[33] | t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind125(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[33] & t[21]);
  assign t[17] = ~(t[22] | t[23]);
  assign t[18] = ~(t[7]);
  assign t[19] = ~(t[34]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[33] | t[24]);
  assign t[23] = ~(t[25]);
  assign t[24] = ~(t[35] & t[26]);
  assign t[25] = ~(t[19] & t[27]);
  assign t[26] = ~(t[34] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[33] | t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind126(x, y);
 input [24:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[33] ^ t[34];
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[35] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[7]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[35] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[37] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[38];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[35] | t[37]);
  assign t[31] = t[39] ^ x[2];
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[12];
  assign t[35] = t[43] ^ x[15];
  assign t[36] = t[44] ^ x[18];
  assign t[37] = t[45] ^ x[21];
  assign t[38] = t[46] ^ x[24];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[3] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[7] : t[12];
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind127(x, y);
 input [25:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[33] ^ t[34];
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[35] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[7]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[35] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[37] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[38];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[35] | t[37]);
  assign t[31] = t[39] ^ x[2];
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[46] = (x[23] & x[24]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[7] : t[12];
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind128(x, y);
 input [25:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[33] ^ t[34];
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[35] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[7]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[35] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[37] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[38];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[35] | t[37]);
  assign t[31] = t[39] ^ x[2];
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[46] = (x[23] & x[24]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[7] : t[12];
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind129(x, y);
 input [25:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[33] ^ t[34];
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[35] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[7]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[35] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[37] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[38];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[35] | t[37]);
  assign t[31] = t[39] ^ x[2];
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[46] = (x[23] & x[24]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = x[6] ? x[7] : t[12];
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind130(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind131(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind132(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind133(x, y);
 input [25:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = t[35] ^ t[36];
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[6]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~(t[5] & t[33]);
  assign t[20] = ~(t[37] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[37] & t[28]);
  assign t[24] = ~(t[38] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[39]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[40]);
  assign t[29] = ~(t[39] | t[31]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[32] & t[40];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[37] | t[38]);
  assign t[33] = t[41] ^ x[2];
  assign t[34] = t[42] ^ x[5];
  assign t[35] = t[43] ^ x[10];
  assign t[36] = t[44] ^ x[13];
  assign t[37] = t[45] ^ x[16];
  assign t[38] = t[46] ^ x[19];
  assign t[39] = t[47] ^ x[22];
  assign t[3] = ~(t[34]);
  assign t[40] = t[48] ^ x[25];
  assign t[41] = (x[0] & x[1]);
  assign t[42] = (x[3] & x[4]);
  assign t[43] = (x[8] & x[9]);
  assign t[44] = (x[11] & x[12]);
  assign t[45] = (x[14] & x[15]);
  assign t[46] = (x[17] & x[18]);
  assign t[47] = (x[20] & x[21]);
  assign t[48] = (x[23] & x[24]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[7] : t[11];
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind134(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[3] & x[7]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind135(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind136(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind137(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(x[6]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[35] | t[23]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[25] & t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[36]);
  assign t[27] = ~(t[38]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[38];
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[27]);
  assign t[31] = ~(t[35] | t[36]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[9];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[34];
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind138(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[9] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind139(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind140(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind141(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind142(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[3] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[9] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind143(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind144(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind145(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[37]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[9];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[16];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = x[6] ? x[10] : t[33];
  assign t[9] = ~(t[2]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind146(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind147(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind148(x, y);
 input [21:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[8];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[15];
  assign t[35] = t[42] ^ x[18];
  assign t[36] = t[43] ^ x[21];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[0] & x[7]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[10] & x[11]);
  assign t[41] = (x[13] & x[14]);
  assign t[42] = (x[16] & x[17]);
  assign t[43] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[9] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind149(x, y);
 input [19:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[7]);
  assign t[16] = ~(t[34] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[7]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[35] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[36] | t[28]);
  assign t[24] = ~(t[36]);
  assign t[25] = t[29] & t[37];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[34] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[35]);
  assign t[31] = ~(t[37]);
  assign t[32] = t[38] ^ x[2];
  assign t[33] = t[39] ^ x[5];
  assign t[34] = t[40] ^ x[10];
  assign t[35] = t[41] ^ x[13];
  assign t[36] = t[42] ^ x[16];
  assign t[37] = t[43] ^ x[19];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[8] & x[9]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[6] : t[33];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind150(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind151(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind152(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind153(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind154(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind155(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind156(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind157(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind158(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind159(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind160(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind161(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[6]);
  assign t[18] = ~(t[34] & t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[35] | t[26]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[27] & t[36];
  assign t[24] = ~(t[22] & t[28]);
  assign t[25] = ~(t[33] & t[29]);
  assign t[26] = ~(t[29]);
  assign t[27] = ~(t[33] | t[34]);
  assign t[28] = ~(t[34]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[9];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[6] ? x[10] : t[32];
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind162(x, y);
 input [22:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[32] | t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[33] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[22]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[34] | t[23]);
  assign t[1] = ~(t[5] & t[29]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[24] & t[35];
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20] & t[28]);
  assign t[26] = ~(t[32] & t[27]);
  assign t[27] = ~(t[35]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[36] ^ x[2];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[37] ^ x[5];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[16];
  assign t[34] = t[41] ^ x[19];
  assign t[35] = t[42] ^ x[22];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = ~(t[30]);
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = x[6] ? x[10] : t[31];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind163(x, y);
 input [22:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[32] | t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[33] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[22]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[34] | t[23]);
  assign t[1] = ~(t[5] & t[29]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[24] & t[35];
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20] & t[28]);
  assign t[26] = ~(t[32] & t[27]);
  assign t[27] = ~(t[35]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[36] ^ x[2];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[37] ^ x[5];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[16];
  assign t[34] = t[41] ^ x[19];
  assign t[35] = t[42] ^ x[22];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = ~(t[30]);
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = x[6] ? x[10] : t[31];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind164(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind165(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind166(x, y);
 input [22:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[32] | t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[33] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[22]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[34] | t[23]);
  assign t[1] = ~(t[5] & t[29]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[24] & t[35];
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20] & t[28]);
  assign t[26] = ~(t[32] & t[27]);
  assign t[27] = ~(t[35]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[36] ^ x[2];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[37] ^ x[5];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[16];
  assign t[34] = t[41] ^ x[19];
  assign t[35] = t[42] ^ x[22];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = ~(t[30]);
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = x[6] ? x[10] : t[31];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind167(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[15]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[15]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[7];
  assign t[34] = t[41] ^ x[11];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[0] & x[6]);
  assign t[41] = (x[9] & x[10]);
  assign t[42] = (x[12] & x[13]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[8] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind168(x, y);
 input [19:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[33] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[34] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[13]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[13]);
  assign t[21] = ~(t[35] | t[25]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[26] & t[36];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[33] & t[29]);
  assign t[29] = ~(t[36]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[34]);
  assign t[31] = t[37] ^ x[2];
  assign t[32] = t[38] ^ x[5];
  assign t[33] = t[39] ^ x[9];
  assign t[34] = t[40] ^ x[12];
  assign t[35] = t[41] ^ x[16];
  assign t[36] = t[42] ^ x[19];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[7] & x[8]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[10] & x[11]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[6] : t[32];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind169(x, y);
 input [22:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[32] | t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[33] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[22]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[34] | t[23]);
  assign t[1] = ~(t[5] & t[29]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[24] & t[35];
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20] & t[28]);
  assign t[26] = ~(t[32] & t[27]);
  assign t[27] = ~(t[35]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[36] ^ x[2];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[37] ^ x[5];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[16];
  assign t[34] = t[41] ^ x[19];
  assign t[35] = t[42] ^ x[22];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = ~(t[30]);
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = x[6] ? x[10] : t[31];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind170(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind171(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind172(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind173(x, y);
 input [22:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[32] | t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[33] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[22]);
  assign t[18] = ~(x[6]);
  assign t[19] = ~(t[34] | t[23]);
  assign t[1] = ~(t[5] & t[29]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[24] & t[35];
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20] & t[28]);
  assign t[26] = ~(t[32] & t[27]);
  assign t[27] = ~(t[35]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[36] ^ x[2];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[37] ^ x[5];
  assign t[31] = t[38] ^ x[9];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[16];
  assign t[34] = t[41] ^ x[19];
  assign t[35] = t[42] ^ x[22];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = ~(t[30]);
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = x[6] ? x[10] : t[31];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind174(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind175(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind176(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind177(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind178(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind179(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind180(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind181(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind182(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind183(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind184(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind185(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind186(x, y);
 input [21:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[9]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[9]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[7];
  assign t[35] = t[42] ^ x[12];
  assign t[36] = t[43] ^ x[15];
  assign t[37] = t[44] ^ x[18];
  assign t[38] = t[45] ^ x[21];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[0] & x[6]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[8] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind187(x, y);
 input [19:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[7]);
  assign t[16] = ~(t[34] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[7]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[35] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[36] | t[28]);
  assign t[24] = ~(t[36]);
  assign t[25] = t[29] & t[37];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[34] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[35]);
  assign t[31] = ~(t[37]);
  assign t[32] = t[38] ^ x[2];
  assign t[33] = t[39] ^ x[5];
  assign t[34] = t[40] ^ x[10];
  assign t[35] = t[41] ^ x[13];
  assign t[36] = t[42] ^ x[16];
  assign t[37] = t[43] ^ x[19];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[8] & x[9]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[14] & x[15]);
  assign t[43] = (x[17] & x[18]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[6] : t[33];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind188(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind189(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind190(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind191(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind192(x, y);
 input [22:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[16]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[16]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[8];
  assign t[34] = t[41] ^ x[12];
  assign t[35] = t[42] ^ x[15];
  assign t[36] = t[43] ^ x[19];
  assign t[37] = t[44] ^ x[22];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[17] & x[18]);
  assign t[44] = (x[20] & x[21]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[9] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind193(x, y);
 input [21:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[2]);
  assign t[11] = ~(t[34] | t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[13]);
  assign t[15] = ~(t[20]);
  assign t[16] = ~(t[35] & t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(x[15]);
  assign t[1] = ~(t[5] & t[31]);
  assign t[20] = ~(x[15]);
  assign t[21] = ~(t[36] | t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = t[26] & t[37];
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[22] & t[30]);
  assign t[28] = ~(t[34] & t[29]);
  assign t[29] = ~(t[37]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[35]);
  assign t[31] = t[38] ^ x[2];
  assign t[32] = t[39] ^ x[5];
  assign t[33] = t[40] ^ x[7];
  assign t[34] = t[41] ^ x[11];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = t[43] ^ x[18];
  assign t[37] = t[44] ^ x[21];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[32]);
  assign t[40] = (x[0] & x[6]);
  assign t[41] = (x[9] & x[10]);
  assign t[42] = (x[12] & x[13]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[4] = ~(t[8] & t[9]);
  assign t[5] = ~(t[8] | t[10]);
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[15] ? x[8] : t[33];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind194(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind195(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind196(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind197(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind198(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind199(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind200(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind201(x, y);
 input [22:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(x[10]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[10]);
  assign t[1] = ~(t[5] & t[32]);
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = t[39] ^ x[2];
  assign t[33] = t[40] ^ x[5];
  assign t[34] = t[41] ^ x[8];
  assign t[35] = t[42] ^ x[13];
  assign t[36] = t[43] ^ x[16];
  assign t[37] = t[44] ^ x[19];
  assign t[38] = t[45] ^ x[22];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[33]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[6] & x[7]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[44] = (x[17] & x[18]);
  assign t[45] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[11] ? x[9] : t[34];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind202(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[15]);
  assign t[11] = ~(x[10]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[7]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(x[10]);
  assign t[17] = ~(t[33] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[33] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[23] & t[27]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[25]);
  assign t[29] = ~(t[33] | t[34]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[8];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] ? x[9] : t[32];
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind203(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[15]);
  assign t[11] = ~(x[10]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[7]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(x[10]);
  assign t[17] = ~(t[33] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[33] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[23] & t[27]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[25]);
  assign t[29] = ~(t[33] | t[34]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[8];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] ? x[9] : t[32];
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind204(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[15]);
  assign t[11] = ~(x[10]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[7]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(x[10]);
  assign t[17] = ~(t[33] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[33] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[23] & t[27]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[25]);
  assign t[29] = ~(t[33] | t[34]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[8];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] ? x[9] : t[32];
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind205(x, y);
 input [22:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[15]);
  assign t[11] = ~(x[10]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[7]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(x[10]);
  assign t[17] = ~(t[33] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[5] & t[30]);
  assign t[20] = ~(t[33] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[23] & t[27]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] | t[28]);
  assign t[27] = t[29] & t[36];
  assign t[28] = ~(t[25]);
  assign t[29] = ~(t[33] | t[34]);
  assign t[2] = ~(t[6]);
  assign t[30] = t[37] ^ x[2];
  assign t[31] = t[38] ^ x[5];
  assign t[32] = t[39] ^ x[8];
  assign t[33] = t[40] ^ x[13];
  assign t[34] = t[41] ^ x[16];
  assign t[35] = t[42] ^ x[19];
  assign t[36] = t[43] ^ x[22];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[31]);
  assign t[40] = (x[11] & x[12]);
  assign t[41] = (x[14] & x[15]);
  assign t[42] = (x[17] & x[18]);
  assign t[43] = (x[20] & x[21]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[7] | t[6]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] ? x[9] : t[32];
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind206(x, y);
 input [41:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[18] ? x[3] : t[42];
  assign t[11] = ~(t[2]);
  assign t[12] = ~(t[43] | t[19]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = t[44] ^ t[45];
  assign t[15] = ~(t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(x[13]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[46] & t[25]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[28] ^ t[29]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(x[13]);
  assign t[25] = ~(t[47] | t[34]);
  assign t[26] = ~(t[35]);
  assign t[27] = t[23] ? t[48] : t[36];
  assign t[28] = t[23] ? t[49] : t[37];
  assign t[29] = t[23] ? t[50] : t[14];
  assign t[2] = ~(t[7] & t[8]);
  assign t[30] = ~(t[47]);
  assign t[31] = t[38] & t[51];
  assign t[32] = ~(t[30] & t[39]);
  assign t[33] = ~(t[43] & t[40]);
  assign t[34] = ~(t[40]);
  assign t[35] = t[23] ? t[52] : t[41];
  assign t[36] = t[53] ^ t[54];
  assign t[37] = t[50] ^ t[55];
  assign t[38] = ~(t[43] | t[46]);
  assign t[39] = ~(t[46]);
  assign t[3] = ~(t[42]);
  assign t[40] = ~(t[51]);
  assign t[41] = t[56] ^ t[57];
  assign t[42] = t[58] ^ x[2];
  assign t[43] = t[59] ^ x[6];
  assign t[44] = t[60] ^ x[9];
  assign t[45] = t[61] ^ x[12];
  assign t[46] = t[62] ^ x[16];
  assign t[47] = t[63] ^ x[19];
  assign t[48] = t[64] ^ x[22];
  assign t[49] = t[65] ^ x[24];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[66] ^ x[26];
  assign t[51] = t[67] ^ x[29];
  assign t[52] = t[68] ^ x[31];
  assign t[53] = t[69] ^ x[33];
  assign t[54] = t[70] ^ x[35];
  assign t[55] = t[71] ^ x[37];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[41];
  assign t[58] = (x[0] & x[1]);
  assign t[59] = (x[4] & x[5]);
  assign t[5] = ~(t[9] | t[11]);
  assign t[60] = (x[7] & x[8]);
  assign t[61] = (x[10] & x[11]);
  assign t[62] = (x[14] & x[15]);
  assign t[63] = (x[17] & x[18]);
  assign t[64] = (x[20] & x[21]);
  assign t[65] = (x[20] & x[23]);
  assign t[66] = (x[7] & x[25]);
  assign t[67] = (x[27] & x[28]);
  assign t[68] = (x[20] & x[30]);
  assign t[69] = (x[7] & x[32]);
  assign t[6] = t[12] ? t[14] : t[13];
  assign t[70] = (x[10] & x[34]);
  assign t[71] = (x[10] & x[36]);
  assign t[72] = (x[7] & x[38]);
  assign t[73] = (x[10] & x[40]);
  assign t[7] = ~(t[12] | t[15]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind207(x, y);
 input [44:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[18] ? x[6] : t[50];
  assign t[11] = ~(t[2]);
  assign t[12] = ~(t[51] | t[19]);
  assign t[13] = ~(t[20] | t[21]);
  assign t[14] = t[52] ^ t[53];
  assign t[15] = ~(t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(x[16]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[54] & t[25]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(x[16]);
  assign t[25] = ~(t[55] | t[34]);
  assign t[26] = ~(t[35] | t[28]);
  assign t[27] = t[36] ? t[38] : t[37];
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[36] ^ t[40]);
  assign t[2] = ~(t[7] & t[8]);
  assign t[30] = ~(t[55]);
  assign t[31] = t[41] & t[56];
  assign t[32] = ~(t[30] & t[42]);
  assign t[33] = ~(t[51] & t[43]);
  assign t[34] = ~(t[43]);
  assign t[35] = ~(t[36] | t[40]);
  assign t[36] = t[23] ? t[57] : t[44];
  assign t[37] = t[23] ? t[58] : t[14];
  assign t[38] = ~(t[37] & t[45]);
  assign t[39] = t[23] ? t[59] : t[46];
  assign t[3] = ~(t[49]);
  assign t[40] = t[23] ? t[60] : t[47];
  assign t[41] = ~(t[51] | t[54]);
  assign t[42] = ~(t[54]);
  assign t[43] = ~(t[56]);
  assign t[44] = t[60] ^ t[61];
  assign t[45] = ~(t[48] & t[28]);
  assign t[46] = t[62] ^ t[63];
  assign t[47] = t[64] ^ t[65];
  assign t[48] = ~(t[40]);
  assign t[49] = t[66] ^ x[2];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[67] ^ x[5];
  assign t[51] = t[68] ^ x[9];
  assign t[52] = t[69] ^ x[12];
  assign t[53] = t[70] ^ x[15];
  assign t[54] = t[71] ^ x[19];
  assign t[55] = t[72] ^ x[22];
  assign t[56] = t[73] ^ x[25];
  assign t[57] = t[74] ^ x[28];
  assign t[58] = t[75] ^ x[30];
  assign t[59] = t[76] ^ x[32];
  assign t[5] = ~(t[9] | t[11]);
  assign t[60] = t[77] ^ x[34];
  assign t[61] = t[78] ^ x[36];
  assign t[62] = t[79] ^ x[38];
  assign t[63] = t[80] ^ x[40];
  assign t[64] = t[81] ^ x[42];
  assign t[65] = t[82] ^ x[44];
  assign t[66] = (x[0] & x[1]);
  assign t[67] = (x[3] & x[4]);
  assign t[68] = (x[7] & x[8]);
  assign t[69] = (x[10] & x[11]);
  assign t[6] = t[12] ? t[14] : t[13];
  assign t[70] = (x[13] & x[14]);
  assign t[71] = (x[17] & x[18]);
  assign t[72] = (x[20] & x[21]);
  assign t[73] = (x[23] & x[24]);
  assign t[74] = (x[26] & x[27]);
  assign t[75] = (x[26] & x[29]);
  assign t[76] = (x[26] & x[31]);
  assign t[77] = (x[10] & x[33]);
  assign t[78] = (x[13] & x[35]);
  assign t[79] = (x[10] & x[37]);
  assign t[7] = ~(t[12] | t[15]);
  assign t[80] = (x[13] & x[39]);
  assign t[81] = (x[10] & x[41]);
  assign t[82] = (x[13] & x[43]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind208(x, y);
 input [44:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[18] ? x[6] : t[54];
  assign t[11] = ~(t[2]);
  assign t[12] = ~(t[55] | t[19]);
  assign t[13] = ~(t[20] & t[21]);
  assign t[14] = t[56] ^ t[57];
  assign t[15] = ~(t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(x[16]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[58] & t[25]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[20] = ~(t[26] & t[27]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(x[16]);
  assign t[25] = ~(t[59] | t[34]);
  assign t[26] = ~(t[35] | t[36]);
  assign t[27] = ~(t[37] & t[38]);
  assign t[28] = ~(t[39] | t[40]);
  assign t[29] = t[41] ? t[27] : t[37];
  assign t[2] = ~(t[7] & t[8]);
  assign t[30] = ~(t[59]);
  assign t[31] = t[42] & t[60];
  assign t[32] = ~(t[30] & t[43]);
  assign t[33] = ~(t[55] & t[44]);
  assign t[34] = ~(t[44]);
  assign t[35] = t[23] ? t[61] : t[14];
  assign t[36] = ~(t[45] | t[46]);
  assign t[37] = t[23] ? t[62] : t[47];
  assign t[38] = ~(t[48] & t[40]);
  assign t[39] = ~(t[41] | t[49]);
  assign t[3] = ~(t[53]);
  assign t[40] = ~(t[35]);
  assign t[41] = t[23] ? t[63] : t[50];
  assign t[42] = ~(t[55] | t[58]);
  assign t[43] = ~(t[58]);
  assign t[44] = ~(t[60]);
  assign t[45] = ~(t[41]);
  assign t[46] = ~(t[48] & t[51]);
  assign t[47] = t[64] ^ t[65];
  assign t[48] = ~(t[49]);
  assign t[49] = t[23] ? t[66] : t[52];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[66] ^ t[67];
  assign t[51] = ~(t[37]);
  assign t[52] = t[68] ^ t[69];
  assign t[53] = t[70] ^ x[2];
  assign t[54] = t[71] ^ x[5];
  assign t[55] = t[72] ^ x[9];
  assign t[56] = t[73] ^ x[12];
  assign t[57] = t[74] ^ x[15];
  assign t[58] = t[75] ^ x[19];
  assign t[59] = t[76] ^ x[22];
  assign t[5] = ~(t[9] | t[11]);
  assign t[60] = t[77] ^ x[25];
  assign t[61] = t[78] ^ x[28];
  assign t[62] = t[79] ^ x[30];
  assign t[63] = t[80] ^ x[32];
  assign t[64] = t[81] ^ x[34];
  assign t[65] = t[82] ^ x[36];
  assign t[66] = t[83] ^ x[38];
  assign t[67] = t[84] ^ x[40];
  assign t[68] = t[85] ^ x[42];
  assign t[69] = t[86] ^ x[44];
  assign t[6] = t[12] ? t[14] : t[13];
  assign t[70] = (x[0] & x[1]);
  assign t[71] = (x[3] & x[4]);
  assign t[72] = (x[7] & x[8]);
  assign t[73] = (x[10] & x[11]);
  assign t[74] = (x[13] & x[14]);
  assign t[75] = (x[17] & x[18]);
  assign t[76] = (x[20] & x[21]);
  assign t[77] = (x[23] & x[24]);
  assign t[78] = (x[26] & x[27]);
  assign t[79] = (x[26] & x[29]);
  assign t[7] = ~(t[12] | t[15]);
  assign t[80] = (x[26] & x[31]);
  assign t[81] = (x[10] & x[33]);
  assign t[82] = (x[13] & x[35]);
  assign t[83] = (x[10] & x[37]);
  assign t[84] = (x[13] & x[39]);
  assign t[85] = (x[10] & x[41]);
  assign t[86] = (x[13] & x[43]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind209(x, y);
 input [44:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[18] ? x[6] : t[50];
  assign t[11] = ~(t[2]);
  assign t[12] = ~(t[51] | t[19]);
  assign t[13] = ~(t[20] & t[21]);
  assign t[14] = t[52] ^ t[53];
  assign t[15] = ~(t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(x[16]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[54] & t[25]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[20] = t[26] ? t[28] : t[27];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = ~(t[33] | t[34]);
  assign t[24] = ~(x[16]);
  assign t[25] = ~(t[55] | t[35]);
  assign t[26] = t[23] ? t[56] : t[14];
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = ~(t[26] | t[40]);
  assign t[2] = ~(t[7] & t[8]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[55]);
  assign t[32] = t[41] & t[57];
  assign t[33] = ~(t[31] & t[42]);
  assign t[34] = ~(t[51] & t[43]);
  assign t[35] = ~(t[43]);
  assign t[36] = t[23] ? t[58] : t[44];
  assign t[37] = ~(t[45] & t[38]);
  assign t[38] = ~(t[46]);
  assign t[39] = ~(t[45] & t[30]);
  assign t[3] = ~(t[49]);
  assign t[40] = t[23] ? t[52] : t[47];
  assign t[41] = ~(t[51] | t[54]);
  assign t[42] = ~(t[54]);
  assign t[43] = ~(t[57]);
  assign t[44] = t[59] ^ t[60];
  assign t[45] = ~(t[40]);
  assign t[46] = t[23] ? t[61] : t[48];
  assign t[47] = t[62] ^ t[63];
  assign t[48] = t[64] ^ t[65];
  assign t[49] = t[66] ^ x[2];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[67] ^ x[5];
  assign t[51] = t[68] ^ x[9];
  assign t[52] = t[69] ^ x[12];
  assign t[53] = t[70] ^ x[15];
  assign t[54] = t[71] ^ x[19];
  assign t[55] = t[72] ^ x[22];
  assign t[56] = t[73] ^ x[25];
  assign t[57] = t[74] ^ x[28];
  assign t[58] = t[75] ^ x[30];
  assign t[59] = t[76] ^ x[32];
  assign t[5] = ~(t[9] | t[11]);
  assign t[60] = t[77] ^ x[34];
  assign t[61] = t[78] ^ x[36];
  assign t[62] = t[79] ^ x[38];
  assign t[63] = t[80] ^ x[40];
  assign t[64] = t[81] ^ x[42];
  assign t[65] = t[82] ^ x[44];
  assign t[66] = (x[0] & x[1]);
  assign t[67] = (x[3] & x[4]);
  assign t[68] = (x[7] & x[8]);
  assign t[69] = (x[10] & x[11]);
  assign t[6] = t[12] ? t[14] : t[13];
  assign t[70] = (x[13] & x[14]);
  assign t[71] = (x[17] & x[18]);
  assign t[72] = (x[20] & x[21]);
  assign t[73] = (x[23] & x[24]);
  assign t[74] = (x[26] & x[27]);
  assign t[75] = (x[23] & x[29]);
  assign t[76] = (x[10] & x[31]);
  assign t[77] = (x[13] & x[33]);
  assign t[78] = (x[23] & x[35]);
  assign t[79] = (x[10] & x[37]);
  assign t[7] = ~(t[12] | t[15]);
  assign t[80] = (x[13] & x[39]);
  assign t[81] = (x[10] & x[41]);
  assign t[82] = (x[13] & x[43]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind210(x, y);
 input [24:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[18] ^ x[3];
  assign t[11] = t[19] ^ x[6];
  assign t[12] = t[20] ^ x[9];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[15];
  assign t[15] = t[23] ^ x[18];
  assign t[16] = t[24] ^ x[21];
  assign t[17] = t[25] ^ x[24];
  assign t[18] = (x[1] & x[2]);
  assign t[19] = (x[4] & x[5]);
  assign t[1] = ~(x[0]);
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[24] = (x[19] & x[20]);
  assign t[25] = (x[22] & x[23]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[7] & t[11];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14] & t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = t[0] & t[1];
endmodule

module R1ind211(x, y);
 input [24:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[28] ^ t[2]);
  assign t[10] = ~(t[31]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14] | t[15]);
  assign t[13] = ~(t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[32] & t[19]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[33]);
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[32] | t[22]);
  assign t[21] = ~(t[23]);
  assign t[22] = ~(t[34] & t[24]);
  assign t[23] = ~(t[17] & t[25]);
  assign t[24] = ~(t[33] | t[26]);
  assign t[25] = t[27] & t[35];
  assign t[26] = ~(t[19]);
  assign t[27] = ~(t[32] | t[34]);
  assign t[28] = t[36] ^ x[2];
  assign t[29] = t[37] ^ x[5];
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = t[38] ^ x[8];
  assign t[31] = t[39] ^ x[12];
  assign t[32] = t[40] ^ x[15];
  assign t[33] = t[41] ^ x[18];
  assign t[34] = t[42] ^ x[21];
  assign t[35] = t[43] ^ x[24];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[6] & x[7]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[4] = ~(t[29]);
  assign t[5] = ~(t[7] & t[30]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(x[9]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind212(x, y);
 input [21:0] x;
 output y;

 wire [39:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[29] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[32]);
  assign t[18] = ~(t[29] | t[20]);
  assign t[19] = ~(t[21]);
  assign t[1] = t[26] ^ t[3];
  assign t[20] = ~(t[31] & t[22]);
  assign t[21] = ~(t[15] & t[23]);
  assign t[22] = ~(t[30] | t[24]);
  assign t[23] = t[25] & t[32];
  assign t[24] = ~(t[17]);
  assign t[25] = ~(t[29] | t[31]);
  assign t[26] = t[33] ^ x[2];
  assign t[27] = t[34] ^ x[5];
  assign t[28] = t[35] ^ x[9];
  assign t[29] = t[36] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[37] ^ x[15];
  assign t[31] = t[38] ^ x[18];
  assign t[32] = t[39] ^ x[21];
  assign t[33] = (x[0] & x[1]);
  assign t[34] = (x[3] & x[4]);
  assign t[35] = (x[7] & x[8]);
  assign t[36] = (x[10] & x[11]);
  assign t[37] = (x[13] & x[14]);
  assign t[38] = (x[16] & x[17]);
  assign t[39] = (x[19] & x[20]);
  assign t[3] = ~(t[5] & t[27]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(x[6]);
  assign t[8] = ~(t[28]);
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind213(x, y);
 input [18:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[2] ^ t[25]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[27] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[27] & t[20]);
  assign t[16] = ~(t[28] & t[21]);
  assign t[17] = ~(t[18] & t[22]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[29] | t[23]);
  assign t[22] = t[24] & t[30];
  assign t[23] = ~(t[20]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = t[31] ^ x[2];
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[9];
  assign t[28] = t[34] ^ x[12];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = t[36] ^ x[18];
  assign t[31] = (x[0] & x[1]);
  assign t[32] = (x[3] & x[4]);
  assign t[33] = (x[7] & x[8]);
  assign t[34] = (x[10] & x[11]);
  assign t[35] = (x[13] & x[14]);
  assign t[36] = (x[16] & x[17]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~(t[26]);
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = ~(x[6]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind214(x, y);
 input [15:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[25] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[17] & t[19]);
  assign t[15] = ~(t[24] & t[20]);
  assign t[16] = ~(t[26] | t[21]);
  assign t[17] = ~(t[26]);
  assign t[18] = t[22] & t[27];
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[20]);
  assign t[22] = ~(t[24] | t[25]);
  assign t[23] = t[28] ^ x[2];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[12];
  assign t[27] = t[32] ^ x[15];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[4] & x[5]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[7] & x[8]);
  assign t[31] = (x[10] & x[11]);
  assign t[32] = (x[13] & x[14]);
  assign t[3] = ~(t[23]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(x[3]);
  assign t[9] = ~(t[24] | t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind215(x, y);
 input [39:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[11] & t[24]);
  assign t[11] = t[25] & t[12];
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17]);
  assign t[15] = ~(t[26]);
  assign t[16] = t[18] & t[27];
  assign t[17] = ~(t[19] | t[20]);
  assign t[18] = ~(t[28] | t[29]);
  assign t[19] = ~(t[30] & t[31]);
  assign t[1] = t[21] ? t[4] : t[3];
  assign t[20] = ~(t[32] & t[33]);
  assign t[21] = t[34] ^ x[2];
  assign t[22] = t[35] ^ x[6];
  assign t[23] = t[36] ^ x[9];
  assign t[24] = t[37] ^ x[12];
  assign t[25] = t[38] ^ x[15];
  assign t[26] = t[39] ^ x[18];
  assign t[27] = t[40] ^ x[21];
  assign t[28] = t[41] ^ x[24];
  assign t[29] = t[42] ^ x[27];
  assign t[2] = ~(x[3]);
  assign t[30] = t[43] ^ x[30];
  assign t[31] = t[44] ^ x[33];
  assign t[32] = t[45] ^ x[36];
  assign t[33] = t[46] ^ x[39];
  assign t[34] = (x[0] & x[1]);
  assign t[35] = (x[4] & x[5]);
  assign t[36] = (x[7] & x[8]);
  assign t[37] = (x[10] & x[11]);
  assign t[38] = (x[13] & x[14]);
  assign t[39] = (x[16] & x[17]);
  assign t[3] = t[5] | t[6];
  assign t[40] = (x[19] & x[20]);
  assign t[41] = (x[22] & x[23]);
  assign t[42] = (x[25] & x[26]);
  assign t[43] = (x[28] & x[29]);
  assign t[44] = (x[31] & x[32]);
  assign t[45] = (x[34] & x[35]);
  assign t[46] = (x[37] & x[38]);
  assign t[4] = ~(t[5] | t[7]);
  assign t[5] = ~(t[22]);
  assign t[6] = ~(t[8] & t[23]);
  assign t[7] = t[9] | t[10];
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[23]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind216(x, y);
 input [36:0] x;
 output y;

 wire [39:0] t;
  assign t[0] = t[2] ^ t[16];
  assign t[10] = ~(t[20]);
  assign t[11] = t[13] & t[21];
  assign t[12] = ~(t[14] | t[15]);
  assign t[13] = ~(t[22] | t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = t[28] ^ x[2];
  assign t[17] = t[29] ^ x[6];
  assign t[18] = t[30] ^ x[9];
  assign t[19] = t[31] ^ x[12];
  assign t[1] = ~(t[3]);
  assign t[20] = t[32] ^ x[15];
  assign t[21] = t[33] ^ x[18];
  assign t[22] = t[34] ^ x[21];
  assign t[23] = t[35] ^ x[24];
  assign t[24] = t[36] ^ x[27];
  assign t[25] = t[37] ^ x[30];
  assign t[26] = t[38] ^ x[33];
  assign t[27] = t[39] ^ x[36];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[4] & x[5]);
  assign t[2] = t[4] | t[5];
  assign t[30] = (x[7] & x[8]);
  assign t[31] = (x[10] & x[11]);
  assign t[32] = (x[13] & x[14]);
  assign t[33] = (x[16] & x[17]);
  assign t[34] = (x[19] & x[20]);
  assign t[35] = (x[22] & x[23]);
  assign t[36] = (x[25] & x[26]);
  assign t[37] = (x[28] & x[29]);
  assign t[38] = (x[31] & x[32]);
  assign t[39] = (x[34] & x[35]);
  assign t[3] = ~(x[3]);
  assign t[4] = ~(t[17]);
  assign t[5] = ~(t[6] & t[18]);
  assign t[6] = t[19] & t[7];
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind217(x, y);
 input [33:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[14];
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[19] | t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = ~(t[23] & t[24]);
  assign t[14] = t[25] ^ x[2];
  assign t[15] = t[26] ^ x[5];
  assign t[16] = t[27] ^ x[9];
  assign t[17] = t[28] ^ x[12];
  assign t[18] = t[29] ^ x[15];
  assign t[19] = t[30] ^ x[18];
  assign t[1] = ~(t[3]);
  assign t[20] = t[31] ^ x[21];
  assign t[21] = t[32] ^ x[24];
  assign t[22] = t[33] ^ x[27];
  assign t[23] = t[34] ^ x[30];
  assign t[24] = t[35] ^ x[33];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[7] & x[8]);
  assign t[28] = (x[10] & x[11]);
  assign t[29] = (x[13] & x[14]);
  assign t[2] = ~(t[4] & t[15]);
  assign t[30] = (x[16] & x[17]);
  assign t[31] = (x[19] & x[20]);
  assign t[32] = (x[22] & x[23]);
  assign t[33] = (x[25] & x[26]);
  assign t[34] = (x[28] & x[29]);
  assign t[35] = (x[31] & x[32]);
  assign t[3] = ~(x[6]);
  assign t[4] = t[16] & t[5];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[17]);
  assign t[9] = t[11] & t[18];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind218(x, y);
 input [30:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2] ^ t[13]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = t[23] ^ x[2];
  assign t[14] = t[24] ^ x[5];
  assign t[15] = t[25] ^ x[9];
  assign t[16] = t[26] ^ x[12];
  assign t[17] = t[27] ^ x[15];
  assign t[18] = t[28] ^ x[18];
  assign t[19] = t[29] ^ x[21];
  assign t[1] = ~(t[3]);
  assign t[20] = t[30] ^ x[24];
  assign t[21] = t[31] ^ x[27];
  assign t[22] = t[32] ^ x[30];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[7] & x[8]);
  assign t[26] = (x[10] & x[11]);
  assign t[27] = (x[13] & x[14]);
  assign t[28] = (x[16] & x[17]);
  assign t[29] = (x[19] & x[20]);
  assign t[2] = t[14] & t[4];
  assign t[30] = (x[22] & x[23]);
  assign t[31] = (x[25] & x[26]);
  assign t[32] = (x[28] & x[29]);
  assign t[3] = ~(x[6]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[15]);
  assign t[8] = t[10] & t[16];
  assign t[9] = ~(t[11] | t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind219(x, y);
 input [27:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[12] ^ t[2]);
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = t[21] ^ x[2];
  assign t[13] = t[22] ^ x[6];
  assign t[14] = t[23] ^ x[9];
  assign t[15] = t[24] ^ x[12];
  assign t[16] = t[25] ^ x[15];
  assign t[17] = t[26] ^ x[18];
  assign t[18] = t[27] ^ x[21];
  assign t[19] = t[28] ^ x[24];
  assign t[1] = ~(t[3]);
  assign t[20] = t[29] ^ x[27];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[4] & x[5]);
  assign t[23] = (x[7] & x[8]);
  assign t[24] = (x[10] & x[11]);
  assign t[25] = (x[13] & x[14]);
  assign t[26] = (x[16] & x[17]);
  assign t[27] = (x[19] & x[20]);
  assign t[28] = (x[22] & x[23]);
  assign t[29] = (x[25] & x[26]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(x[3]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[9] & t[14];
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind220(x, y);
 input [24:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(x[0]);
  assign t[10] = ~(t[19] & t[20]);
  assign t[11] = ~(t[21] & t[22]);
  assign t[12] = ~(t[18] | t[13]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17]);
  assign t[15] = t[23] ^ x[3];
  assign t[16] = t[24] ^ x[6];
  assign t[17] = t[25] ^ x[9];
  assign t[18] = t[26] ^ x[12];
  assign t[19] = t[27] ^ x[15];
  assign t[1] = ~(t[2] & t[3]);
  assign t[20] = t[28] ^ x[18];
  assign t[21] = t[29] ^ x[21];
  assign t[22] = t[30] ^ x[24];
  assign t[23] = (x[1] & x[2]);
  assign t[24] = (x[4] & x[5]);
  assign t[25] = (x[7] & x[8]);
  assign t[26] = (x[10] & x[11]);
  assign t[27] = (x[13] & x[14]);
  assign t[28] = (x[16] & x[17]);
  assign t[29] = (x[19] & x[20]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = (x[22] & x[23]);
  assign t[3] = ~(t[6] & t[7]);
  assign t[4] = ~(t[15] | t[16]);
  assign t[5] = ~(t[8] | t[17]);
  assign t[6] = ~(t[15] | t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[18]);
  assign t[9] = ~(t[16] & t[12]);
  assign y = t[0] & t[1];
endmodule

module R1ind221(x, y);
 input [39:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[36]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19] & t[10]);
  assign t[16] = ~(t[37] & t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[37] | t[25]);
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[40] & t[41]);
  assign t[24] = ~(t[42] & t[43]);
  assign t[25] = ~(t[36] & t[27]);
  assign t[26] = ~(t[19] & t[28]);
  assign t[27] = ~(t[38] | t[29]);
  assign t[28] = t[30] & t[39];
  assign t[29] = ~(t[20]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[37] | t[36]);
  assign t[31] = t[44] ^ x[3];
  assign t[32] = t[45] ^ x[6];
  assign t[33] = t[46] ^ x[9];
  assign t[34] = t[47] ^ x[12];
  assign t[35] = t[48] ^ x[15];
  assign t[36] = t[49] ^ x[18];
  assign t[37] = t[50] ^ x[21];
  assign t[38] = t[51] ^ x[24];
  assign t[39] = t[52] ^ x[27];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[53] ^ x[30];
  assign t[41] = t[54] ^ x[33];
  assign t[42] = t[55] ^ x[36];
  assign t[43] = t[56] ^ x[39];
  assign t[44] = (x[1] & x[2]);
  assign t[45] = (x[4] & x[5]);
  assign t[46] = (x[7] & x[8]);
  assign t[47] = (x[10] & x[11]);
  assign t[48] = (x[13] & x[14]);
  assign t[49] = (x[16] & x[17]);
  assign t[4] = ~(t[10] | t[11]);
  assign t[50] = (x[19] & x[20]);
  assign t[51] = (x[22] & x[23]);
  assign t[52] = (x[25] & x[26]);
  assign t[53] = (x[28] & x[29]);
  assign t[54] = (x[31] & x[32]);
  assign t[55] = (x[34] & x[35]);
  assign t[56] = (x[37] & x[38]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[31] & t[32]);
  assign t[7] = ~(t[33] & t[34]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[35] & t[5]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind222(x, y);
 input [39:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[33]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[34] & t[35]);
  assign t[15] = ~(t[36] & t[37]);
  assign t[16] = ~(t[24]);
  assign t[17] = ~(t[38] & t[7]);
  assign t[18] = ~(t[39] & t[40]);
  assign t[19] = ~(t[41] & t[42]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[43] | t[25]);
  assign t[21] = ~(t[26]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[27] | t[33]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[25] = ~(t[44] & t[30]);
  assign t[26] = ~(t[27] & t[31]);
  assign t[27] = ~(t[45]);
  assign t[28] = ~(t[27] & t[32]);
  assign t[29] = ~(t[43] & t[10]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[45] | t[4]);
  assign t[31] = t[22] & t[33];
  assign t[32] = ~(t[44]);
  assign t[33] = t[46] ^ x[3];
  assign t[34] = t[47] ^ x[6];
  assign t[35] = t[48] ^ x[9];
  assign t[36] = t[49] ^ x[12];
  assign t[37] = t[50] ^ x[15];
  assign t[38] = t[51] ^ x[18];
  assign t[39] = t[52] ^ x[21];
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = t[53] ^ x[24];
  assign t[41] = t[54] ^ x[27];
  assign t[42] = t[55] ^ x[30];
  assign t[43] = t[56] ^ x[33];
  assign t[44] = t[57] ^ x[36];
  assign t[45] = t[58] ^ x[39];
  assign t[46] = (x[1] & x[2]);
  assign t[47] = (x[4] & x[5]);
  assign t[48] = (x[7] & x[8]);
  assign t[49] = (x[10] & x[11]);
  assign t[4] = ~(t[10]);
  assign t[50] = (x[13] & x[14]);
  assign t[51] = (x[16] & x[17]);
  assign t[52] = (x[19] & x[20]);
  assign t[53] = (x[22] & x[23]);
  assign t[54] = (x[25] & x[26]);
  assign t[55] = (x[28] & x[29]);
  assign t[56] = (x[31] & x[32]);
  assign t[57] = (x[34] & x[35]);
  assign t[58] = (x[37] & x[38]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12] & t[13]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[14] | t[15]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1_ind(x, y);
 input [510:0] x;
 output [222:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[142], x[141], x[191], x[190], x[149], x[148], x[147], x[146], x[145], x[140], x[139], x[144], x[143], x[138], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[146], x[145], x[176], x[175], x[142], x[141], x[191], x[190], x[144], x[143], x[140], x[139], x[138], x[149], x[148], x[147], x[185], x[184], x[187], x[186], x[181], x[180], x[183], x[182], x[179], x[194], x[177], x[189], x[188], x[174], x[193], x[192], x[171]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[146], x[145], x[176], x[175], x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[140], x[139], x[185], x[184], x[144], x[143], x[189], x[188], x[142], x[141], x[138], x[149], x[148], x[147], x[183], x[182], x[181], x[180], x[187], x[186], x[179], x[197], x[177], x[191], x[190], x[174], x[196], x[195], x[171]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[142], x[141], x[191], x[190], x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[146], x[145], x[176], x[175], x[187], x[186], x[144], x[143], x[189], x[188], x[149], x[148], x[147], x[181], x[180], x[140], x[139], x[138], x[183], x[182], x[179], x[200], x[177], x[185], x[184], x[174], x[199], x[198], x[171]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[204], x[199], x[198], x[177], x[173], x[172], x[171], x[203], x[202], x[201]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[207], x[176], x[175], x[174], x[177], x[193], x[192], x[171], x[206], x[205], x[201]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[210], x[189], x[188], x[174], x[177], x[196], x[195], x[171], x[209], x[208], x[201]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[213], x[191], x[190], x[174], x[177], x[199], x[198], x[171], x[212], x[211], x[201]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[217], x[212], x[211], x[177], x[203], x[202], x[201], x[216], x[215], x[214]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[220], x[173], x[172], x[171], x[177], x[206], x[205], x[201], x[219], x[218], x[214]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[223], x[193], x[192], x[171], x[177], x[209], x[208], x[201], x[222], x[221], x[214]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[226], x[196], x[195], x[171], x[177], x[212], x[211], x[201], x[225], x[224], x[214]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[230], x[225], x[224], x[177], x[216], x[215], x[214], x[229], x[228], x[227]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[233], x[203], x[202], x[201], x[177], x[219], x[218], x[214], x[232], x[231], x[227]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[236], x[206], x[205], x[201], x[177], x[222], x[221], x[214], x[235], x[234], x[227]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[239], x[209], x[208], x[201], x[177], x[225], x[224], x[214], x[238], x[237], x[227]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[243], x[238], x[237], x[177], x[229], x[228], x[227], x[242], x[241], x[240]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[246], x[216], x[215], x[214], x[177], x[232], x[231], x[227], x[245], x[244], x[240]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[249], x[219], x[218], x[214], x[177], x[235], x[234], x[227], x[248], x[247], x[240]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[252], x[222], x[221], x[214], x[177], x[238], x[237], x[227], x[251], x[250], x[240]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[256], x[251], x[250], x[177], x[242], x[241], x[240], x[255], x[254], x[253]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[259], x[229], x[228], x[227], x[177], x[245], x[244], x[240], x[258], x[257], x[253]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[262], x[232], x[231], x[227], x[177], x[248], x[247], x[240], x[261], x[260], x[253]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[265], x[235], x[234], x[227], x[177], x[251], x[250], x[240], x[264], x[263], x[253]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[269], x[264], x[263], x[177], x[255], x[254], x[253], x[268], x[267], x[266]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[272], x[242], x[241], x[240], x[177], x[258], x[257], x[253], x[271], x[270], x[266]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[275], x[245], x[244], x[240], x[177], x[261], x[260], x[253], x[274], x[273], x[266]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[278], x[248], x[247], x[240], x[177], x[264], x[263], x[253], x[277], x[276], x[266]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[282], x[277], x[276], x[177], x[268], x[267], x[266], x[281], x[280], x[279]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[285], x[255], x[254], x[253], x[177], x[271], x[270], x[266], x[284], x[283], x[279]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[288], x[258], x[257], x[253], x[177], x[274], x[273], x[266], x[287], x[286], x[279]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[291], x[261], x[260], x[253], x[177], x[277], x[276], x[266], x[290], x[289], x[279]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[295], x[290], x[289], x[177], x[281], x[280], x[279], x[294], x[293], x[292]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[298], x[268], x[267], x[266], x[177], x[284], x[283], x[279], x[297], x[296], x[292]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[301], x[271], x[270], x[266], x[177], x[287], x[286], x[279], x[300], x[299], x[292]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[304], x[274], x[273], x[266], x[177], x[290], x[289], x[279], x[303], x[302], x[292]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[308], x[303], x[302], x[177], x[294], x[293], x[292], x[307], x[306], x[305]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[311], x[281], x[280], x[279], x[177], x[297], x[296], x[292], x[310], x[309], x[305]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[314], x[284], x[283], x[279], x[177], x[300], x[299], x[292], x[313], x[312], x[305]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[317], x[287], x[286], x[279], x[177], x[303], x[302], x[292], x[316], x[315], x[305]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[321], x[316], x[315], x[177], x[307], x[306], x[305], x[320], x[319], x[318]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[324], x[294], x[293], x[292], x[177], x[310], x[309], x[305], x[323], x[322], x[318]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[327], x[297], x[296], x[292], x[177], x[313], x[312], x[305], x[326], x[325], x[318]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[330], x[300], x[299], x[292], x[177], x[316], x[315], x[305], x[329], x[328], x[318]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[334], x[329], x[328], x[177], x[320], x[319], x[318], x[333], x[332], x[331]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[337], x[307], x[306], x[305], x[177], x[323], x[322], x[318], x[336], x[335], x[331]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[340], x[310], x[309], x[305], x[177], x[326], x[325], x[318], x[339], x[338], x[331]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[343], x[313], x[312], x[305], x[177], x[329], x[328], x[318], x[342], x[341], x[331]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[347], x[342], x[341], x[177], x[333], x[332], x[331], x[346], x[345], x[344]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[350], x[320], x[319], x[318], x[177], x[336], x[335], x[331], x[349], x[348], x[344]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[353], x[323], x[322], x[318], x[177], x[339], x[338], x[331], x[352], x[351], x[344]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[356], x[326], x[325], x[318], x[177], x[342], x[341], x[331], x[355], x[354], x[344]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[360], x[355], x[354], x[177], x[346], x[345], x[344], x[359], x[358], x[357]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[363], x[333], x[332], x[331], x[177], x[349], x[348], x[344], x[362], x[361], x[357]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[366], x[336], x[335], x[331], x[177], x[352], x[351], x[344], x[365], x[364], x[357]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[369], x[339], x[338], x[331], x[177], x[355], x[354], x[344], x[368], x[367], x[357]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[373], x[368], x[367], x[177], x[359], x[358], x[357], x[372], x[371], x[370]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[376], x[346], x[345], x[344], x[177], x[362], x[361], x[357], x[375], x[374], x[370]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[379], x[349], x[348], x[344], x[177], x[365], x[364], x[357], x[378], x[377], x[370]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[382], x[352], x[351], x[344], x[177], x[368], x[367], x[357], x[381], x[380], x[370]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[381], x[380], x[389], x[388], x[387], x[386], x[177], x[372], x[371], x[370], x[385], x[384], x[383]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[359], x[358], x[357], x[395], x[394], x[393], x[392], x[177], x[375], x[374], x[370], x[391], x[390], x[383]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[362], x[361], x[357], x[401], x[400], x[399], x[398], x[177], x[378], x[377], x[370], x[397], x[396], x[383]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[365], x[364], x[357], x[407], x[406], x[405], x[404], x[177], x[381], x[380], x[370], x[403], x[402], x[383]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[411], x[403], x[402], x[177], x[385], x[384], x[383], x[410], x[409], x[408]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[414], x[372], x[371], x[370], x[177], x[391], x[390], x[383], x[413], x[412], x[408]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[417], x[375], x[374], x[370], x[177], x[397], x[396], x[383], x[416], x[415], x[408]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[378], x[377], x[370], x[423], x[422], x[421], x[420], x[177], x[403], x[402], x[383], x[419], x[418], x[408]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[427], x[419], x[418], x[177], x[410], x[409], x[408], x[426], x[425], x[424]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[430], x[385], x[384], x[383], x[177], x[413], x[412], x[408], x[429], x[428], x[424]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[433], x[391], x[390], x[383], x[177], x[416], x[415], x[408], x[432], x[431], x[424]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[436], x[397], x[396], x[383], x[177], x[419], x[418], x[408], x[435], x[434], x[424]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[437], x[435], x[434], x[177], x[426], x[425], x[424], x[181], x[180], x[179]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[438], x[410], x[409], x[408], x[177], x[429], x[428], x[424], x[187], x[186], x[179]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[439], x[413], x[412], x[408], x[177], x[432], x[431], x[424], x[183], x[182], x[179]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[442], x[416], x[415], x[408], x[177], x[435], x[434], x[424], x[441], x[440], x[179]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[443], x[441], x[440], x[177], x[181], x[180], x[179], x[176], x[175], x[174]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[444], x[426], x[425], x[424], x[177], x[187], x[186], x[179], x[189], x[188], x[174]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[445], x[429], x[428], x[424], x[177], x[183], x[182], x[179], x[191], x[190], x[174]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[446], x[432], x[431], x[424], x[177], x[441], x[440], x[179], x[185], x[184], x[174]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[447], x[113], x[112], x[111], x[146], x[145], x[138], x[137], x[136], x[129]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[448], x[122], x[121], x[120], x[144], x[143], x[138], x[135], x[134], x[129]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[449], x[131], x[130], x[177], x[142], x[141], x[138], x[133], x[132], x[129]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[450], x[140], x[139], x[138], x[131], x[130], x[129]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[451], x[77], x[76], x[75], x[177], x[137], x[136], x[129], x[128], x[127], x[120]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[452], x[86], x[85], x[84], x[177], x[135], x[134], x[129], x[126], x[125], x[120]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[453], x[95], x[94], x[93], x[177], x[133], x[132], x[129], x[124], x[123], x[120]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[454], x[104], x[103], x[102], x[177], x[131], x[130], x[129], x[122], x[121], x[120]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[455], x[41], x[40], x[39], x[177], x[128], x[127], x[120], x[119], x[118], x[111]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[456], x[50], x[49], x[48], x[177], x[126], x[125], x[120], x[117], x[116], x[111]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[457], x[59], x[58], x[57], x[177], x[124], x[123], x[120], x[115], x[114], x[111]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[458], x[68], x[67], x[66], x[177], x[122], x[121], x[120], x[113], x[112], x[111]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[459], x[11], x[10], x[3], x[119], x[118], x[111], x[110], x[109], x[102]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[460], x[14], x[13], x[12], x[117], x[116], x[111], x[108], x[107], x[102]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[461], x[23], x[22], x[21], x[115], x[114], x[111], x[106], x[105], x[102]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[462], x[32], x[31], x[30], x[177], x[113], x[112], x[111], x[104], x[103], x[102]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[463], x[115], x[114], x[111], x[177], x[110], x[109], x[102], x[101], x[100], x[93]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[464], x[124], x[123], x[120], x[177], x[108], x[107], x[102], x[99], x[98], x[93]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[465], x[133], x[132], x[129], x[106], x[105], x[102], x[97], x[96], x[93]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[466], x[142], x[141], x[138], x[104], x[103], x[102], x[95], x[94], x[93]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[467], x[79], x[78], x[75], x[177], x[101], x[100], x[93], x[92], x[91], x[84]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[468], x[88], x[87], x[99], x[98], x[93], x[90], x[89], x[84]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[469], x[97], x[96], x[93], x[88], x[87], x[84]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[470], x[106], x[105], x[102], x[177], x[95], x[94], x[93], x[86], x[85], x[84]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[471], x[43], x[42], x[39], x[92], x[91], x[84], x[83], x[82], x[75]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[472], x[52], x[51], x[48], x[90], x[89], x[84], x[81], x[80], x[75]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[473], x[61], x[60], x[57], x[88], x[87], x[84], x[79], x[78], x[75]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[474], x[70], x[69], x[66], x[177], x[86], x[85], x[84], x[77], x[76], x[75]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[475], x[9], x[8], x[3], x[83], x[82], x[75], x[74], x[73], x[66]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[476], x[16], x[15], x[12], x[81], x[80], x[75], x[72], x[71], x[66]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[477], x[25], x[24], x[21], x[79], x[78], x[75], x[70], x[69], x[66]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[478], x[34], x[33], x[30], x[77], x[76], x[75], x[68], x[67], x[66]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[479], x[117], x[116], x[111], x[74], x[73], x[66], x[65], x[64], x[57]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[480], x[126], x[125], x[120], x[72], x[71], x[66], x[63], x[62], x[57]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[481], x[135], x[134], x[129], x[70], x[69], x[66], x[61], x[60], x[57]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[482], x[144], x[143], x[138], x[68], x[67], x[66], x[59], x[58], x[57]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[483], x[81], x[80], x[75], x[65], x[64], x[57], x[56], x[55], x[48]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[484], x[90], x[89], x[84], x[63], x[62], x[57], x[54], x[53], x[48]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[485], x[99], x[98], x[93], x[61], x[60], x[57], x[52], x[51], x[48]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[486], x[108], x[107], x[102], x[59], x[58], x[57], x[50], x[49], x[48]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[487], x[45], x[44], x[56], x[55], x[48], x[47], x[46], x[39]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[488], x[54], x[53], x[48], x[45], x[44], x[39]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[489], x[63], x[62], x[57], x[52], x[51], x[48], x[43], x[42], x[39]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[490], x[72], x[71], x[66], x[50], x[49], x[48], x[41], x[40], x[39]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[491], x[7], x[6], x[3], x[47], x[46], x[39], x[38], x[37], x[30]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[492], x[18], x[17], x[12], x[45], x[44], x[39], x[36], x[35], x[30]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[493], x[27], x[26], x[21], x[43], x[42], x[39], x[34], x[33], x[30]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[152], x[151], x[150], x[149], x[148], x[147], x[494], x[36], x[35], x[41], x[40], x[39], x[32], x[31], x[30]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[495], x[119], x[118], x[111], x[38], x[37], x[30], x[29], x[28], x[21]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[496], x[128], x[127], x[120], x[36], x[35], x[30], x[27], x[26], x[21]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[497], x[137], x[136], x[129], x[34], x[33], x[30], x[25], x[24], x[21]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[498], x[146], x[145], x[138], x[32], x[31], x[30], x[23], x[22], x[21]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[499], x[83], x[82], x[75], x[29], x[28], x[21], x[20], x[19], x[12]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[500], x[92], x[91], x[84], x[27], x[26], x[21], x[18], x[17], x[12]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[501], x[101], x[100], x[93], x[25], x[24], x[21], x[16], x[15], x[12]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[502], x[110], x[109], x[102], x[23], x[22], x[21], x[14], x[13], x[12]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[503], x[47], x[46], x[39], x[20], x[19], x[12], x[5], x[4], x[3]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[504], x[56], x[55], x[48], x[18], x[17], x[12], x[7], x[6], x[3]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[505], x[65], x[64], x[57], x[16], x[15], x[12], x[9], x[8], x[3]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[506], x[74], x[73], x[66], x[14], x[13], x[12], x[11], x[10], x[3]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[142], x[141], x[191], x[190], x[140], x[139], x[144], x[143], x[189], x[188], x[187], x[186], x[155], x[154], x[153], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[158], x[157], x[156], x[152], x[151], x[150], x[177], x[146], x[145], x[138], x[176], x[175], x[174], x[149], x[148], x[147], x[507], x[5], x[4], x[3]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[146], x[145], x[176], x[175], x[142], x[141], x[191], x[190], x[140], x[139], x[185], x[184], x[187], x[186], x[181], x[180], x[183], x[182], x[179], x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[177], x[144], x[143], x[138], x[189], x[188], x[174], x[149], x[148], x[147], x[508], x[20], x[19], x[12], x[7], x[6], x[3]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[146], x[145], x[176], x[175], x[140], x[139], x[185], x[184], x[144], x[143], x[189], x[188], x[183], x[182], x[181], x[180], x[187], x[186], x[179], x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[177], x[142], x[141], x[138], x[191], x[190], x[174], x[149], x[148], x[147], x[509], x[29], x[28], x[21], x[9], x[8], x[3]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[142], x[141], x[191], x[190], x[146], x[145], x[176], x[175], x[187], x[186], x[144], x[143], x[189], x[188], x[181], x[180], x[155], x[154], x[153], x[183], x[182], x[179], x[158], x[157], x[156], x[152], x[151], x[150], x[177], x[140], x[139], x[138], x[185], x[184], x[174], x[149], x[148], x[147], x[510], x[38], x[37], x[30], x[11], x[10], x[3]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[152], x[151], x[150], x[149], x[148], x[147], x[155], x[154], x[153], x[158], x[157], x[156], x[177]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[167], x[166], x[165], x[177], x[170], x[169], x[168], x[161], x[160], x[159], x[164], x[163], x[162]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[155], x[154], x[153], x[152], x[151], x[150], x[158], x[157], x[156], x[149], x[148], x[147], x[167], x[166], x[165], x[177], x[170], x[169], x[168], x[161], x[160], x[159]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[167], x[166], x[165], x[170], x[169], x[168]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[155], x[154], x[153], x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[177], x[167], x[166], x[165]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[152], x[151], x[150], x[149], x[148], x[147], x[155], x[154], x[153], x[158], x[157], x[156], x[423], x[422], x[421], x[389], x[388], x[387], x[395], x[394], x[393], x[401], x[400], x[399], x[177], x[407], x[406], x[405]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[152], x[151], x[150], x[149], x[148], x[147], x[155], x[154], x[153], x[158], x[157], x[156], x[423], x[422], x[421], x[389], x[388], x[387], x[395], x[394], x[393], x[177], x[401], x[400], x[399]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[152], x[151], x[150], x[149], x[148], x[147], x[155], x[154], x[153], x[158], x[157], x[156], x[423], x[422], x[421], x[177], x[389], x[388], x[387], x[395], x[394], x[393]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[152], x[151], x[150], x[149], x[148], x[147], x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[423], x[422], x[421], x[389], x[388], x[387]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[152], x[151], x[150], x[149], x[148], x[147], x[155], x[154], x[153], x[158], x[157], x[156], x[177], x[423], x[422], x[421]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[177]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[155], x[154], x[153], x[158], x[157], x[156], x[149], x[148], x[147], x[152], x[151], x[150], x[423], x[422], x[421], x[407], x[406], x[405], x[395], x[394], x[393], x[401], x[400], x[399], x[389], x[388], x[387], x[177]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[158], x[157], x[156], x[152], x[151], x[150], x[149], x[148], x[147], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[423], x[422], x[421], x[407], x[406], x[405], x[395], x[394], x[393], x[401], x[400], x[399], x[389], x[388], x[387], x[155], x[154], x[153], x[177]}), .y(y[222]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [23:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[20] & t[21]);
  assign t[11] = ~(t[17] | t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[14];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[23];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[1];
  assign t[39] = t[55] ^ x[2];
  assign t[3] = ~(t[14] | t[15]);
  assign t[40] = t[56] ^ x[4];
  assign t[41] = t[57] ^ x[5];
  assign t[42] = t[58] ^ x[7];
  assign t[43] = t[59] ^ x[8];
  assign t[44] = t[60] ^ x[10];
  assign t[45] = t[61] ^ x[11];
  assign t[46] = t[62] ^ x[13];
  assign t[47] = t[63] ^ x[14];
  assign t[48] = t[64] ^ x[16];
  assign t[49] = t[65] ^ x[17];
  assign t[4] = ~(t[7] | t[16]);
  assign t[50] = t[66] ^ x[19];
  assign t[51] = t[67] ^ x[20];
  assign t[52] = t[68] ^ x[22];
  assign t[53] = t[69] ^ x[23];
  assign t[54] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[0]);
  assign t[56] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[3]);
  assign t[58] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[14] | t[8]);
  assign t[60] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[9]);
  assign t[62] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[12]);
  assign t[64] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[15]);
  assign t[66] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[18]);
  assign t[68] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[17]);
  assign t[8] = ~(t[15] & t[11]);
  assign t[9] = ~(t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [23:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[20] & t[21]);
  assign t[11] = ~(t[17] | t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[16]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[14];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[23];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[1];
  assign t[39] = t[55] ^ x[2];
  assign t[3] = ~(t[14] | t[15]);
  assign t[40] = t[56] ^ x[4];
  assign t[41] = t[57] ^ x[5];
  assign t[42] = t[58] ^ x[7];
  assign t[43] = t[59] ^ x[8];
  assign t[44] = t[60] ^ x[10];
  assign t[45] = t[61] ^ x[11];
  assign t[46] = t[62] ^ x[13];
  assign t[47] = t[63] ^ x[14];
  assign t[48] = t[64] ^ x[16];
  assign t[49] = t[65] ^ x[17];
  assign t[4] = ~(t[7] | t[16]);
  assign t[50] = t[66] ^ x[19];
  assign t[51] = t[67] ^ x[20];
  assign t[52] = t[68] ^ x[22];
  assign t[53] = t[69] ^ x[23];
  assign t[54] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[55] = (x[0]);
  assign t[56] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[3]);
  assign t[58] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[14] | t[8]);
  assign t[60] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[9]);
  assign t[62] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[12]);
  assign t[64] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[15]);
  assign t[66] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[18]);
  assign t[68] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[17]);
  assign t[8] = ~(t[15] & t[11]);
  assign t[9] = ~(t[18] & t[19]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = (t[19]);
  assign t[12] = (t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[28] ^ x[6];
  assign t[21] = t[29] ^ x[9];
  assign t[22] = t[30] ^ x[12];
  assign t[23] = t[31] ^ x[15];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[24];
  assign t[27] = (~t[35] & t[36]);
  assign t[28] = (~t[37] & t[38]);
  assign t[29] = (~t[39] & t[40]);
  assign t[2] = ~(x[0]);
  assign t[30] = (~t[41] & t[42]);
  assign t[31] = (~t[43] & t[44]);
  assign t[32] = (~t[45] & t[46]);
  assign t[33] = (~t[47] & t[48]);
  assign t[34] = (~t[49] & t[50]);
  assign t[35] = t[51] ^ x[2];
  assign t[36] = t[52] ^ x[3];
  assign t[37] = t[53] ^ x[5];
  assign t[38] = t[54] ^ x[6];
  assign t[39] = t[55] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[9];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[12];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[15];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[18];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[21];
  assign t[49] = t[65] ^ x[23];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[24];
  assign t[51] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[1]);
  assign t[53] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[4]);
  assign t[55] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[7]);
  assign t[57] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[10]);
  assign t[59] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[13]);
  assign t[61] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[16]);
  assign t[63] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[19]);
  assign t[65] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[22]);
  assign t[6] = t[8] & t[12];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[15] & t[16]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = (t[19]);
  assign t[12] = (t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[28] ^ x[6];
  assign t[21] = t[29] ^ x[9];
  assign t[22] = t[30] ^ x[12];
  assign t[23] = t[31] ^ x[15];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[24];
  assign t[27] = (~t[35] & t[36]);
  assign t[28] = (~t[37] & t[38]);
  assign t[29] = (~t[39] & t[40]);
  assign t[2] = ~(x[0]);
  assign t[30] = (~t[41] & t[42]);
  assign t[31] = (~t[43] & t[44]);
  assign t[32] = (~t[45] & t[46]);
  assign t[33] = (~t[47] & t[48]);
  assign t[34] = (~t[49] & t[50]);
  assign t[35] = t[51] ^ x[2];
  assign t[36] = t[52] ^ x[3];
  assign t[37] = t[53] ^ x[5];
  assign t[38] = t[54] ^ x[6];
  assign t[39] = t[55] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[9];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[12];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[15];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[18];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[21];
  assign t[49] = t[65] ^ x[23];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[24];
  assign t[51] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[1]);
  assign t[53] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[4]);
  assign t[55] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[7]);
  assign t[57] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[10]);
  assign t[59] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[13]);
  assign t[61] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[16]);
  assign t[63] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[19]);
  assign t[65] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[22]);
  assign t[6] = t[8] & t[12];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[15] & t[16]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [39:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[4]);
  assign t[101] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[7]);
  assign t[103] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[10]);
  assign t[105] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[13]);
  assign t[107] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[16]);
  assign t[109] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[36] & t[6]);
  assign t[110] = (x[19]);
  assign t[111] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[22]);
  assign t[113] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[25]);
  assign t[115] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[28]);
  assign t[117] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[31]);
  assign t[119] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[37]);
  assign t[120] = (x[34]);
  assign t[121] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[37]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20] & t[11]);
  assign t[17] = ~(t[38] & t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[38] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[41] & t[42]);
  assign t[25] = ~(t[43] & t[44]);
  assign t[26] = ~(t[37] & t[28]);
  assign t[27] = ~(t[20] & t[29]);
  assign t[28] = ~(t[39] | t[30]);
  assign t[29] = t[31] & t[40];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[38] | t[37]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = t[58] ^ x[3];
  assign t[46] = t[59] ^ x[6];
  assign t[47] = t[60] ^ x[9];
  assign t[48] = t[61] ^ x[12];
  assign t[49] = t[62] ^ x[15];
  assign t[4] = ~(t[9] | t[10]);
  assign t[50] = t[63] ^ x[18];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[24];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[30];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[36];
  assign t[57] = t[70] ^ x[39];
  assign t[58] = (~t[71] & t[72]);
  assign t[59] = (~t[73] & t[74]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[60] = (~t[75] & t[76]);
  assign t[61] = (~t[77] & t[78]);
  assign t[62] = (~t[79] & t[80]);
  assign t[63] = (~t[81] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[85] & t[86]);
  assign t[66] = (~t[87] & t[88]);
  assign t[67] = (~t[89] & t[90]);
  assign t[68] = (~t[91] & t[92]);
  assign t[69] = (~t[93] & t[94]);
  assign t[6] = ~(x[0]);
  assign t[70] = (~t[95] & t[96]);
  assign t[71] = t[97] ^ x[2];
  assign t[72] = t[98] ^ x[3];
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[6];
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[9];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[12];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[32] & t[33]);
  assign t[80] = t[106] ^ x[15];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[18];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[21];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[24];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[27];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = ~(t[34] & t[35]);
  assign t[90] = t[116] ^ x[30];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[33];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[36];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[39];
  assign t[97] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[1]);
  assign t[99] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [39:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[4]);
  assign t[101] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[7]);
  assign t[103] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[10]);
  assign t[105] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[13]);
  assign t[107] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[16]);
  assign t[109] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[36] & t[6]);
  assign t[110] = (x[19]);
  assign t[111] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[22]);
  assign t[113] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[25]);
  assign t[115] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[28]);
  assign t[117] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[31]);
  assign t[119] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[37]);
  assign t[120] = (x[34]);
  assign t[121] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[37]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20] & t[11]);
  assign t[17] = ~(t[38] & t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[38] | t[26]);
  assign t[23] = ~(t[27]);
  assign t[24] = ~(t[41] & t[42]);
  assign t[25] = ~(t[43] & t[44]);
  assign t[26] = ~(t[37] & t[28]);
  assign t[27] = ~(t[20] & t[29]);
  assign t[28] = ~(t[39] | t[30]);
  assign t[29] = t[31] & t[40];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[38] | t[37]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = t[58] ^ x[3];
  assign t[46] = t[59] ^ x[6];
  assign t[47] = t[60] ^ x[9];
  assign t[48] = t[61] ^ x[12];
  assign t[49] = t[62] ^ x[15];
  assign t[4] = ~(t[9] | t[10]);
  assign t[50] = t[63] ^ x[18];
  assign t[51] = t[64] ^ x[21];
  assign t[52] = t[65] ^ x[24];
  assign t[53] = t[66] ^ x[27];
  assign t[54] = t[67] ^ x[30];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[36];
  assign t[57] = t[70] ^ x[39];
  assign t[58] = (~t[71] & t[72]);
  assign t[59] = (~t[73] & t[74]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[60] = (~t[75] & t[76]);
  assign t[61] = (~t[77] & t[78]);
  assign t[62] = (~t[79] & t[80]);
  assign t[63] = (~t[81] & t[82]);
  assign t[64] = (~t[83] & t[84]);
  assign t[65] = (~t[85] & t[86]);
  assign t[66] = (~t[87] & t[88]);
  assign t[67] = (~t[89] & t[90]);
  assign t[68] = (~t[91] & t[92]);
  assign t[69] = (~t[93] & t[94]);
  assign t[6] = ~(x[0]);
  assign t[70] = (~t[95] & t[96]);
  assign t[71] = t[97] ^ x[2];
  assign t[72] = t[98] ^ x[3];
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[6];
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[9];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[12];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[32] & t[33]);
  assign t[80] = t[106] ^ x[15];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[18];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[21];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[24];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[27];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = ~(t[34] & t[35]);
  assign t[90] = t[116] ^ x[30];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[33];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[36];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[39];
  assign t[97] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[1]);
  assign t[99] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [24:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[13]);
  assign t[11] = ~(t[20] & t[21]);
  assign t[12] = ~(t[22] & t[23]);
  assign t[13] = ~(t[19] | t[14]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(x[0]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = t[32] ^ x[3];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = t[36] ^ x[15];
  assign t[29] = t[37] ^ x[18];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = t[38] ^ x[21];
  assign t[31] = t[39] ^ x[24];
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[42] & t[43]);
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[2];
  assign t[41] = t[57] ^ x[3];
  assign t[42] = t[58] ^ x[5];
  assign t[43] = t[59] ^ x[6];
  assign t[44] = t[60] ^ x[8];
  assign t[45] = t[61] ^ x[9];
  assign t[46] = t[62] ^ x[11];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[14];
  assign t[49] = t[65] ^ x[15];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[66] ^ x[17];
  assign t[51] = t[67] ^ x[18];
  assign t[52] = t[68] ^ x[20];
  assign t[53] = t[69] ^ x[21];
  assign t[54] = t[70] ^ x[23];
  assign t[55] = t[71] ^ x[24];
  assign t[56] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[1]);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[16] | t[17]);
  assign t[60] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[7]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[13]);
  assign t[66] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[16]);
  assign t[68] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[9] | t[18]);
  assign t[70] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[22]);
  assign t[7] = ~(t[16] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [24:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[13]);
  assign t[11] = ~(t[20] & t[21]);
  assign t[12] = ~(t[22] & t[23]);
  assign t[13] = ~(t[19] | t[14]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(x[0]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = t[32] ^ x[3];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[9];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = t[36] ^ x[15];
  assign t[29] = t[37] ^ x[18];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = t[38] ^ x[21];
  assign t[31] = t[39] ^ x[24];
  assign t[32] = (~t[40] & t[41]);
  assign t[33] = (~t[42] & t[43]);
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[2];
  assign t[41] = t[57] ^ x[3];
  assign t[42] = t[58] ^ x[5];
  assign t[43] = t[59] ^ x[6];
  assign t[44] = t[60] ^ x[8];
  assign t[45] = t[61] ^ x[9];
  assign t[46] = t[62] ^ x[11];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[14];
  assign t[49] = t[65] ^ x[15];
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = t[66] ^ x[17];
  assign t[51] = t[67] ^ x[18];
  assign t[52] = t[68] ^ x[20];
  assign t[53] = t[69] ^ x[21];
  assign t[54] = t[70] ^ x[23];
  assign t[55] = t[71] ^ x[24];
  assign t[56] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[1]);
  assign t[58] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[16] | t[17]);
  assign t[60] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[7]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[13]);
  assign t[66] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[16]);
  assign t[68] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[9] | t[18]);
  assign t[70] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[22]);
  assign t[7] = ~(t[16] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[19]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [39:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[1]);
  assign t[101] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[4]);
  assign t[103] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[7]);
  assign t[105] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[10]);
  assign t[107] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[13]);
  assign t[109] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = (x[16]);
  assign t[111] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[19]);
  assign t[113] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[22]);
  assign t[115] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[25]);
  assign t[117] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[28]);
  assign t[119] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[34]);
  assign t[120] = (x[31]);
  assign t[121] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[34]);
  assign t[123] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[37]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[21] | t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[35] & t[36]);
  assign t[16] = ~(t[37] & t[38]);
  assign t[17] = ~(t[25]);
  assign t[18] = ~(t[39] & t[8]);
  assign t[19] = ~(t[40] & t[41]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[42] & t[43]);
  assign t[21] = ~(t[44] | t[26]);
  assign t[22] = ~(t[27]);
  assign t[23] = ~(t[44] | t[45]);
  assign t[24] = ~(t[28] | t[34]);
  assign t[25] = ~(t[29] | t[30]);
  assign t[26] = ~(t[45] & t[31]);
  assign t[27] = ~(t[28] & t[32]);
  assign t[28] = ~(t[46]);
  assign t[29] = ~(t[28] & t[33]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[44] & t[11]);
  assign t[31] = ~(t[46] | t[5]);
  assign t[32] = t[23] & t[34];
  assign t[33] = ~(t[45]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[3];
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[9];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[63] ^ x[12];
  assign t[51] = t[64] ^ x[15];
  assign t[52] = t[65] ^ x[18];
  assign t[53] = t[66] ^ x[21];
  assign t[54] = t[67] ^ x[24];
  assign t[55] = t[68] ^ x[27];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[33];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[39];
  assign t[5] = ~(t[11]);
  assign t[60] = (~t[73] & t[74]);
  assign t[61] = (~t[75] & t[76]);
  assign t[62] = (~t[77] & t[78]);
  assign t[63] = (~t[79] & t[80]);
  assign t[64] = (~t[81] & t[82]);
  assign t[65] = (~t[83] & t[84]);
  assign t[66] = (~t[85] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[89] & t[90]);
  assign t[69] = (~t[91] & t[92]);
  assign t[6] = ~(t[12]);
  assign t[70] = (~t[93] & t[94]);
  assign t[71] = (~t[95] & t[96]);
  assign t[72] = (~t[97] & t[98]);
  assign t[73] = t[99] ^ x[2];
  assign t[74] = t[100] ^ x[3];
  assign t[75] = t[101] ^ x[5];
  assign t[76] = t[102] ^ x[6];
  assign t[77] = t[103] ^ x[8];
  assign t[78] = t[104] ^ x[9];
  assign t[79] = t[105] ^ x[11];
  assign t[7] = ~(t[13] & t[14]);
  assign t[80] = t[106] ^ x[12];
  assign t[81] = t[107] ^ x[14];
  assign t[82] = t[108] ^ x[15];
  assign t[83] = t[109] ^ x[17];
  assign t[84] = t[110] ^ x[18];
  assign t[85] = t[111] ^ x[20];
  assign t[86] = t[112] ^ x[21];
  assign t[87] = t[113] ^ x[23];
  assign t[88] = t[114] ^ x[24];
  assign t[89] = t[115] ^ x[26];
  assign t[8] = ~(x[0]);
  assign t[90] = t[116] ^ x[27];
  assign t[91] = t[117] ^ x[29];
  assign t[92] = t[118] ^ x[30];
  assign t[93] = t[119] ^ x[32];
  assign t[94] = t[120] ^ x[33];
  assign t[95] = t[121] ^ x[35];
  assign t[96] = t[122] ^ x[36];
  assign t[97] = t[123] ^ x[38];
  assign t[98] = t[124] ^ x[39];
  assign t[99] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[15] | t[16]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [39:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[1]);
  assign t[101] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[4]);
  assign t[103] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[7]);
  assign t[105] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[10]);
  assign t[107] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[13]);
  assign t[109] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = (x[16]);
  assign t[111] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[19]);
  assign t[113] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[22]);
  assign t[115] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[25]);
  assign t[117] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[28]);
  assign t[119] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(t[34]);
  assign t[120] = (x[31]);
  assign t[121] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[34]);
  assign t[123] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[37]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[21] | t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[35] & t[36]);
  assign t[16] = ~(t[37] & t[38]);
  assign t[17] = ~(t[25]);
  assign t[18] = ~(t[39] & t[8]);
  assign t[19] = ~(t[40] & t[41]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[42] & t[43]);
  assign t[21] = ~(t[44] | t[26]);
  assign t[22] = ~(t[27]);
  assign t[23] = ~(t[44] | t[45]);
  assign t[24] = ~(t[28] | t[34]);
  assign t[25] = ~(t[29] | t[30]);
  assign t[26] = ~(t[45] & t[31]);
  assign t[27] = ~(t[28] & t[32]);
  assign t[28] = ~(t[46]);
  assign t[29] = ~(t[28] & t[33]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[44] & t[11]);
  assign t[31] = ~(t[46] | t[5]);
  assign t[32] = t[23] & t[34];
  assign t[33] = ~(t[45]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[3];
  assign t[48] = t[61] ^ x[6];
  assign t[49] = t[62] ^ x[9];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[63] ^ x[12];
  assign t[51] = t[64] ^ x[15];
  assign t[52] = t[65] ^ x[18];
  assign t[53] = t[66] ^ x[21];
  assign t[54] = t[67] ^ x[24];
  assign t[55] = t[68] ^ x[27];
  assign t[56] = t[69] ^ x[30];
  assign t[57] = t[70] ^ x[33];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[39];
  assign t[5] = ~(t[11]);
  assign t[60] = (~t[73] & t[74]);
  assign t[61] = (~t[75] & t[76]);
  assign t[62] = (~t[77] & t[78]);
  assign t[63] = (~t[79] & t[80]);
  assign t[64] = (~t[81] & t[82]);
  assign t[65] = (~t[83] & t[84]);
  assign t[66] = (~t[85] & t[86]);
  assign t[67] = (~t[87] & t[88]);
  assign t[68] = (~t[89] & t[90]);
  assign t[69] = (~t[91] & t[92]);
  assign t[6] = ~(t[12]);
  assign t[70] = (~t[93] & t[94]);
  assign t[71] = (~t[95] & t[96]);
  assign t[72] = (~t[97] & t[98]);
  assign t[73] = t[99] ^ x[2];
  assign t[74] = t[100] ^ x[3];
  assign t[75] = t[101] ^ x[5];
  assign t[76] = t[102] ^ x[6];
  assign t[77] = t[103] ^ x[8];
  assign t[78] = t[104] ^ x[9];
  assign t[79] = t[105] ^ x[11];
  assign t[7] = ~(t[13] & t[14]);
  assign t[80] = t[106] ^ x[12];
  assign t[81] = t[107] ^ x[14];
  assign t[82] = t[108] ^ x[15];
  assign t[83] = t[109] ^ x[17];
  assign t[84] = t[110] ^ x[18];
  assign t[85] = t[111] ^ x[20];
  assign t[86] = t[112] ^ x[21];
  assign t[87] = t[113] ^ x[23];
  assign t[88] = t[114] ^ x[24];
  assign t[89] = t[115] ^ x[26];
  assign t[8] = ~(x[0]);
  assign t[90] = t[116] ^ x[27];
  assign t[91] = t[117] ^ x[29];
  assign t[92] = t[118] ^ x[30];
  assign t[93] = t[119] ^ x[32];
  assign t[94] = t[120] ^ x[33];
  assign t[95] = t[121] ^ x[35];
  assign t[96] = t[122] ^ x[36];
  assign t[97] = t[123] ^ x[38];
  assign t[98] = t[124] ^ x[39];
  assign t[99] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[15] | t[16]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [39:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[22]);
  assign t[103] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[25]);
  assign t[105] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[28]);
  assign t[107] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[31]);
  assign t[109] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[24]);
  assign t[110] = (x[34]);
  assign t[111] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[37]);
  assign t[11] = ~(t[12] & t[25]);
  assign t[12] = t[26] & t[13];
  assign t[13] = ~(t[14] | t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[27]);
  assign t[17] = t[19] & t[28];
  assign t[18] = ~(t[20] | t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[31] & t[32]);
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = (t[35]);
  assign t[23] = (t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = t[22] ? t[5] : t[4];
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = t[48] ^ x[2];
  assign t[36] = t[49] ^ x[6];
  assign t[37] = t[50] ^ x[9];
  assign t[38] = t[51] ^ x[12];
  assign t[39] = t[52] ^ x[15];
  assign t[3] = ~(x[3]);
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[24];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[30];
  assign t[45] = t[58] ^ x[33];
  assign t[46] = t[59] ^ x[36];
  assign t[47] = t[60] ^ x[39];
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[63] & t[64]);
  assign t[4] = t[6] | t[7];
  assign t[50] = (~t[65] & t[66]);
  assign t[51] = (~t[67] & t[68]);
  assign t[52] = (~t[69] & t[70]);
  assign t[53] = (~t[71] & t[72]);
  assign t[54] = (~t[73] & t[74]);
  assign t[55] = (~t[75] & t[76]);
  assign t[56] = (~t[77] & t[78]);
  assign t[57] = (~t[79] & t[80]);
  assign t[58] = (~t[81] & t[82]);
  assign t[59] = (~t[83] & t[84]);
  assign t[5] = ~(t[6] | t[8]);
  assign t[60] = (~t[85] & t[86]);
  assign t[61] = t[87] ^ x[1];
  assign t[62] = t[88] ^ x[2];
  assign t[63] = t[89] ^ x[5];
  assign t[64] = t[90] ^ x[6];
  assign t[65] = t[91] ^ x[8];
  assign t[66] = t[92] ^ x[9];
  assign t[67] = t[93] ^ x[11];
  assign t[68] = t[94] ^ x[12];
  assign t[69] = t[95] ^ x[14];
  assign t[6] = ~(t[23]);
  assign t[70] = t[96] ^ x[15];
  assign t[71] = t[97] ^ x[17];
  assign t[72] = t[98] ^ x[18];
  assign t[73] = t[99] ^ x[20];
  assign t[74] = t[100] ^ x[21];
  assign t[75] = t[101] ^ x[23];
  assign t[76] = t[102] ^ x[24];
  assign t[77] = t[103] ^ x[26];
  assign t[78] = t[104] ^ x[27];
  assign t[79] = t[105] ^ x[29];
  assign t[7] = ~(t[9] & t[24]);
  assign t[80] = t[106] ^ x[30];
  assign t[81] = t[107] ^ x[32];
  assign t[82] = t[108] ^ x[33];
  assign t[83] = t[109] ^ x[35];
  assign t[84] = t[110] ^ x[36];
  assign t[85] = t[111] ^ x[38];
  assign t[86] = t[112] ^ x[39];
  assign t[87] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[0]);
  assign t[89] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = t[10] | t[11];
  assign t[90] = (x[4]);
  assign t[91] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[7]);
  assign t[93] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[10]);
  assign t[95] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[13]);
  assign t[97] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[16]);
  assign t[99] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind31(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind34(x, y);
 input [39:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[102] = (x[22]);
  assign t[103] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[104] = (x[25]);
  assign t[105] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[106] = (x[28]);
  assign t[107] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[31]);
  assign t[109] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[24]);
  assign t[110] = (x[34]);
  assign t[111] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[37]);
  assign t[11] = ~(t[12] & t[25]);
  assign t[12] = t[26] & t[13];
  assign t[13] = ~(t[14] | t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[27]);
  assign t[17] = t[19] & t[28];
  assign t[18] = ~(t[20] | t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[31] & t[32]);
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = (t[35]);
  assign t[23] = (t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = t[22] ? t[5] : t[4];
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = t[48] ^ x[2];
  assign t[36] = t[49] ^ x[6];
  assign t[37] = t[50] ^ x[9];
  assign t[38] = t[51] ^ x[12];
  assign t[39] = t[52] ^ x[15];
  assign t[3] = ~(x[3]);
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[24];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[30];
  assign t[45] = t[58] ^ x[33];
  assign t[46] = t[59] ^ x[36];
  assign t[47] = t[60] ^ x[39];
  assign t[48] = (~t[61] & t[62]);
  assign t[49] = (~t[63] & t[64]);
  assign t[4] = t[6] | t[7];
  assign t[50] = (~t[65] & t[66]);
  assign t[51] = (~t[67] & t[68]);
  assign t[52] = (~t[69] & t[70]);
  assign t[53] = (~t[71] & t[72]);
  assign t[54] = (~t[73] & t[74]);
  assign t[55] = (~t[75] & t[76]);
  assign t[56] = (~t[77] & t[78]);
  assign t[57] = (~t[79] & t[80]);
  assign t[58] = (~t[81] & t[82]);
  assign t[59] = (~t[83] & t[84]);
  assign t[5] = ~(t[6] | t[8]);
  assign t[60] = (~t[85] & t[86]);
  assign t[61] = t[87] ^ x[1];
  assign t[62] = t[88] ^ x[2];
  assign t[63] = t[89] ^ x[5];
  assign t[64] = t[90] ^ x[6];
  assign t[65] = t[91] ^ x[8];
  assign t[66] = t[92] ^ x[9];
  assign t[67] = t[93] ^ x[11];
  assign t[68] = t[94] ^ x[12];
  assign t[69] = t[95] ^ x[14];
  assign t[6] = ~(t[23]);
  assign t[70] = t[96] ^ x[15];
  assign t[71] = t[97] ^ x[17];
  assign t[72] = t[98] ^ x[18];
  assign t[73] = t[99] ^ x[20];
  assign t[74] = t[100] ^ x[21];
  assign t[75] = t[101] ^ x[23];
  assign t[76] = t[102] ^ x[24];
  assign t[77] = t[103] ^ x[26];
  assign t[78] = t[104] ^ x[27];
  assign t[79] = t[105] ^ x[29];
  assign t[7] = ~(t[9] & t[24]);
  assign t[80] = t[106] ^ x[30];
  assign t[81] = t[107] ^ x[32];
  assign t[82] = t[108] ^ x[33];
  assign t[83] = t[109] ^ x[35];
  assign t[84] = t[110] ^ x[36];
  assign t[85] = t[111] ^ x[38];
  assign t[86] = t[112] ^ x[39];
  assign t[87] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[0]);
  assign t[89] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = t[10] | t[11];
  assign t[90] = (x[4]);
  assign t[91] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[7]);
  assign t[93] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[10]);
  assign t[95] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[13]);
  assign t[97] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[16]);
  assign t[99] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [33:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[12] & t[19];
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = (t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = t[3] ^ t[15];
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[9];
  assign t[29] = t[40] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] ^ x[15];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[24];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[30];
  assign t[36] = t[47] ^ x[33];
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[5] & t[16]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = (~t[58] & t[59]);
  assign t[43] = (~t[60] & t[61]);
  assign t[44] = (~t[62] & t[63]);
  assign t[45] = (~t[64] & t[65]);
  assign t[46] = (~t[66] & t[67]);
  assign t[47] = (~t[68] & t[69]);
  assign t[48] = t[70] ^ x[1];
  assign t[49] = t[71] ^ x[2];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[4];
  assign t[51] = t[73] ^ x[5];
  assign t[52] = t[74] ^ x[8];
  assign t[53] = t[75] ^ x[9];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[12];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[15];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[18];
  assign t[5] = t[17] & t[6];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[21];
  assign t[62] = t[84] ^ x[23];
  assign t[63] = t[85] ^ x[24];
  assign t[64] = t[86] ^ x[26];
  assign t[65] = t[87] ^ x[27];
  assign t[66] = t[88] ^ x[29];
  assign t[67] = t[89] ^ x[30];
  assign t[68] = t[90] ^ x[32];
  assign t[69] = t[91] ^ x[33];
  assign t[6] = ~(t[7] | t[8]);
  assign t[70] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[0]);
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[7]);
  assign t[76] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[10]);
  assign t[78] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[16]);
  assign t[82] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[19]);
  assign t[84] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[22]);
  assign t[86] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[25]);
  assign t[88] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[28]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[31]);
  assign t[9] = ~(t[18]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind36(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind37(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind38(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind39(x, y);
 input [33:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[12] & t[19];
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = (t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = t[3] ^ t[15];
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[9];
  assign t[29] = t[40] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] ^ x[15];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[24];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[30];
  assign t[36] = t[47] ^ x[33];
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[5] & t[16]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = (~t[58] & t[59]);
  assign t[43] = (~t[60] & t[61]);
  assign t[44] = (~t[62] & t[63]);
  assign t[45] = (~t[64] & t[65]);
  assign t[46] = (~t[66] & t[67]);
  assign t[47] = (~t[68] & t[69]);
  assign t[48] = t[70] ^ x[1];
  assign t[49] = t[71] ^ x[2];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[4];
  assign t[51] = t[73] ^ x[5];
  assign t[52] = t[74] ^ x[8];
  assign t[53] = t[75] ^ x[9];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[12];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[15];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[18];
  assign t[5] = t[17] & t[6];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[21];
  assign t[62] = t[84] ^ x[23];
  assign t[63] = t[85] ^ x[24];
  assign t[64] = t[86] ^ x[26];
  assign t[65] = t[87] ^ x[27];
  assign t[66] = t[88] ^ x[29];
  assign t[67] = t[89] ^ x[30];
  assign t[68] = t[90] ^ x[32];
  assign t[69] = t[91] ^ x[33];
  assign t[6] = ~(t[7] | t[8]);
  assign t[70] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[0]);
  assign t[72] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[3]);
  assign t[74] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[7]);
  assign t[76] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[10]);
  assign t[78] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[16]);
  assign t[82] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[19]);
  assign t[84] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[22]);
  assign t[86] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[25]);
  assign t[88] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[28]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[31]);
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [30:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = (t[24]);
  assign t[15] = (t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[12];
  assign t[28] = t[38] ^ x[15];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[24];
  assign t[32] = t[42] ^ x[27];
  assign t[33] = t[43] ^ x[30];
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = t[15] & t[5];
  assign t[40] = (~t[56] & t[57]);
  assign t[41] = (~t[58] & t[59]);
  assign t[42] = (~t[60] & t[61]);
  assign t[43] = (~t[62] & t[63]);
  assign t[44] = t[64] ^ x[1];
  assign t[45] = t[65] ^ x[2];
  assign t[46] = t[66] ^ x[4];
  assign t[47] = t[67] ^ x[5];
  assign t[48] = t[68] ^ x[8];
  assign t[49] = t[69] ^ x[9];
  assign t[4] = ~(x[6]);
  assign t[50] = t[70] ^ x[11];
  assign t[51] = t[71] ^ x[12];
  assign t[52] = t[72] ^ x[14];
  assign t[53] = t[73] ^ x[15];
  assign t[54] = t[74] ^ x[17];
  assign t[55] = t[75] ^ x[18];
  assign t[56] = t[76] ^ x[20];
  assign t[57] = t[77] ^ x[21];
  assign t[58] = t[78] ^ x[23];
  assign t[59] = t[79] ^ x[24];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[80] ^ x[26];
  assign t[61] = t[81] ^ x[27];
  assign t[62] = t[82] ^ x[29];
  assign t[63] = t[83] ^ x[30];
  assign t[64] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[0]);
  assign t[66] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[3]);
  assign t[68] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[10]);
  assign t[72] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[13]);
  assign t[74] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[16]);
  assign t[76] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[19]);
  assign t[78] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[22]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[25]);
  assign t[82] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[28]);
  assign t[8] = ~(t[16]);
  assign t[9] = t[11] & t[17];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind41(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind42(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind43(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind44(x, y);
 input [30:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = (t[24]);
  assign t[15] = (t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[12];
  assign t[28] = t[38] ^ x[15];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[24];
  assign t[32] = t[42] ^ x[27];
  assign t[33] = t[43] ^ x[30];
  assign t[34] = (~t[44] & t[45]);
  assign t[35] = (~t[46] & t[47]);
  assign t[36] = (~t[48] & t[49]);
  assign t[37] = (~t[50] & t[51]);
  assign t[38] = (~t[52] & t[53]);
  assign t[39] = (~t[54] & t[55]);
  assign t[3] = t[15] & t[5];
  assign t[40] = (~t[56] & t[57]);
  assign t[41] = (~t[58] & t[59]);
  assign t[42] = (~t[60] & t[61]);
  assign t[43] = (~t[62] & t[63]);
  assign t[44] = t[64] ^ x[1];
  assign t[45] = t[65] ^ x[2];
  assign t[46] = t[66] ^ x[4];
  assign t[47] = t[67] ^ x[5];
  assign t[48] = t[68] ^ x[8];
  assign t[49] = t[69] ^ x[9];
  assign t[4] = ~(x[6]);
  assign t[50] = t[70] ^ x[11];
  assign t[51] = t[71] ^ x[12];
  assign t[52] = t[72] ^ x[14];
  assign t[53] = t[73] ^ x[15];
  assign t[54] = t[74] ^ x[17];
  assign t[55] = t[75] ^ x[18];
  assign t[56] = t[76] ^ x[20];
  assign t[57] = t[77] ^ x[21];
  assign t[58] = t[78] ^ x[23];
  assign t[59] = t[79] ^ x[24];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[80] ^ x[26];
  assign t[61] = t[81] ^ x[27];
  assign t[62] = t[82] ^ x[29];
  assign t[63] = t[83] ^ x[30];
  assign t[64] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[0]);
  assign t[66] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[3]);
  assign t[68] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[10]);
  assign t[72] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[13]);
  assign t[74] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[16]);
  assign t[76] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[19]);
  assign t[78] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[22]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[25]);
  assign t[82] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[28]);
  assign t[8] = ~(t[16]);
  assign t[9] = t[11] & t[17];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [27:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[13] ^ t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = t[31] ^ x[2];
  assign t[23] = t[32] ^ x[6];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[18];
  assign t[28] = t[37] ^ x[21];
  assign t[29] = t[38] ^ x[24];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[27];
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = (~t[54] & t[55]);
  assign t[39] = (~t[56] & t[57]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[1];
  assign t[41] = t[59] ^ x[2];
  assign t[42] = t[60] ^ x[5];
  assign t[43] = t[61] ^ x[6];
  assign t[44] = t[62] ^ x[8];
  assign t[45] = t[63] ^ x[9];
  assign t[46] = t[64] ^ x[11];
  assign t[47] = t[65] ^ x[12];
  assign t[48] = t[66] ^ x[14];
  assign t[49] = t[67] ^ x[15];
  assign t[4] = ~(x[3]);
  assign t[50] = t[68] ^ x[17];
  assign t[51] = t[69] ^ x[18];
  assign t[52] = t[70] ^ x[20];
  assign t[53] = t[71] ^ x[21];
  assign t[54] = t[72] ^ x[23];
  assign t[55] = t[73] ^ x[24];
  assign t[56] = t[74] ^ x[26];
  assign t[57] = t[75] ^ x[27];
  assign t[58] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[0]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[4]);
  assign t[62] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[7]);
  assign t[64] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[10]);
  assign t[66] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[13]);
  assign t[68] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[19]);
  assign t[72] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[22]);
  assign t[74] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[25]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[10] & t[15];
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind46(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind47(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind48(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind49(x, y);
 input [27:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[13] ^ t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = t[31] ^ x[2];
  assign t[23] = t[32] ^ x[6];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[18];
  assign t[28] = t[37] ^ x[21];
  assign t[29] = t[38] ^ x[24];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[27];
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = (~t[54] & t[55]);
  assign t[39] = (~t[56] & t[57]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[1];
  assign t[41] = t[59] ^ x[2];
  assign t[42] = t[60] ^ x[5];
  assign t[43] = t[61] ^ x[6];
  assign t[44] = t[62] ^ x[8];
  assign t[45] = t[63] ^ x[9];
  assign t[46] = t[64] ^ x[11];
  assign t[47] = t[65] ^ x[12];
  assign t[48] = t[66] ^ x[14];
  assign t[49] = t[67] ^ x[15];
  assign t[4] = ~(x[3]);
  assign t[50] = t[68] ^ x[17];
  assign t[51] = t[69] ^ x[18];
  assign t[52] = t[70] ^ x[20];
  assign t[53] = t[71] ^ x[21];
  assign t[54] = t[72] ^ x[23];
  assign t[55] = t[73] ^ x[24];
  assign t[56] = t[74] ^ x[26];
  assign t[57] = t[75] ^ x[27];
  assign t[58] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[0]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[4]);
  assign t[62] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[7]);
  assign t[64] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[10]);
  assign t[66] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[13]);
  assign t[68] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[19]);
  assign t[72] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[22]);
  assign t[74] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[25]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[10] & t[15];
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[34]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[21]);
  assign t[12] = t[14] & t[22];
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[23] | t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[3] ^ t[17];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[4]);
  assign t[30] = t[42] ^ x[6];
  assign t[31] = t[43] ^ x[9];
  assign t[32] = t[44] ^ x[12];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[18];
  assign t[35] = t[47] ^ x[21];
  assign t[36] = t[48] ^ x[24];
  assign t[37] = t[49] ^ x[27];
  assign t[38] = t[50] ^ x[30];
  assign t[39] = t[51] ^ x[33];
  assign t[3] = t[5] | t[6];
  assign t[40] = t[52] ^ x[36];
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = (~t[73] & t[74]);
  assign t[52] = (~t[75] & t[76]);
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[5];
  assign t[56] = t[80] ^ x[6];
  assign t[57] = t[81] ^ x[8];
  assign t[58] = t[82] ^ x[9];
  assign t[59] = t[83] ^ x[11];
  assign t[5] = ~(t[18]);
  assign t[60] = t[84] ^ x[12];
  assign t[61] = t[85] ^ x[14];
  assign t[62] = t[86] ^ x[15];
  assign t[63] = t[87] ^ x[17];
  assign t[64] = t[88] ^ x[18];
  assign t[65] = t[89] ^ x[20];
  assign t[66] = t[90] ^ x[21];
  assign t[67] = t[91] ^ x[23];
  assign t[68] = t[92] ^ x[24];
  assign t[69] = t[93] ^ x[26];
  assign t[6] = ~(t[7] & t[19]);
  assign t[70] = t[94] ^ x[27];
  assign t[71] = t[95] ^ x[29];
  assign t[72] = t[96] ^ x[30];
  assign t[73] = t[97] ^ x[32];
  assign t[74] = t[98] ^ x[33];
  assign t[75] = t[99] ^ x[35];
  assign t[76] = t[100] ^ x[36];
  assign t[77] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[0]);
  assign t[79] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[20] & t[8];
  assign t[80] = (x[4]);
  assign t[81] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[7]);
  assign t[83] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[10]);
  assign t[85] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[13]);
  assign t[87] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[16]);
  assign t[89] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] | t[10]);
  assign t[90] = (x[19]);
  assign t[91] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[22]);
  assign t[93] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[25]);
  assign t[95] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[28]);
  assign t[97] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[31]);
  assign t[99] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11] & t[12]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind51(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind52(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind53(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind54(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[34]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[21]);
  assign t[12] = t[14] & t[22];
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[23] | t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[3] ^ t[17];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[4]);
  assign t[30] = t[42] ^ x[6];
  assign t[31] = t[43] ^ x[9];
  assign t[32] = t[44] ^ x[12];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[18];
  assign t[35] = t[47] ^ x[21];
  assign t[36] = t[48] ^ x[24];
  assign t[37] = t[49] ^ x[27];
  assign t[38] = t[50] ^ x[30];
  assign t[39] = t[51] ^ x[33];
  assign t[3] = t[5] | t[6];
  assign t[40] = t[52] ^ x[36];
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = (~t[73] & t[74]);
  assign t[52] = (~t[75] & t[76]);
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[5];
  assign t[56] = t[80] ^ x[6];
  assign t[57] = t[81] ^ x[8];
  assign t[58] = t[82] ^ x[9];
  assign t[59] = t[83] ^ x[11];
  assign t[5] = ~(t[18]);
  assign t[60] = t[84] ^ x[12];
  assign t[61] = t[85] ^ x[14];
  assign t[62] = t[86] ^ x[15];
  assign t[63] = t[87] ^ x[17];
  assign t[64] = t[88] ^ x[18];
  assign t[65] = t[89] ^ x[20];
  assign t[66] = t[90] ^ x[21];
  assign t[67] = t[91] ^ x[23];
  assign t[68] = t[92] ^ x[24];
  assign t[69] = t[93] ^ x[26];
  assign t[6] = ~(t[7] & t[19]);
  assign t[70] = t[94] ^ x[27];
  assign t[71] = t[95] ^ x[29];
  assign t[72] = t[96] ^ x[30];
  assign t[73] = t[97] ^ x[32];
  assign t[74] = t[98] ^ x[33];
  assign t[75] = t[99] ^ x[35];
  assign t[76] = t[100] ^ x[36];
  assign t[77] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[0]);
  assign t[79] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = t[20] & t[8];
  assign t[80] = (x[4]);
  assign t[81] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[7]);
  assign t[83] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[10]);
  assign t[85] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[13]);
  assign t[87] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[16]);
  assign t[89] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[9] | t[10]);
  assign t[90] = (x[19]);
  assign t[91] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[22]);
  assign t[93] = (x[25] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0 & ~1'b0) | (x[25] & 1'b0 & ~1'b0 & 1'b0) | (x[25] & ~1'b0 & 1'b0 & 1'b0) | (~x[25] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[25]);
  assign t[95] = (x[28] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[28] & 1'b0 & ~1'b0 & ~1'b0) | (~x[28] & ~1'b0 & 1'b0 & ~1'b0) | (~x[28] & ~1'b0 & ~1'b0 & 1'b0) | (x[28] & 1'b0 & 1'b0 & ~1'b0) | (x[28] & 1'b0 & ~1'b0 & 1'b0) | (x[28] & ~1'b0 & 1'b0 & 1'b0) | (~x[28] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[28]);
  assign t[97] = (x[31] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[31] & 1'b0 & ~1'b0 & ~1'b0) | (~x[31] & ~1'b0 & 1'b0 & ~1'b0) | (~x[31] & ~1'b0 & ~1'b0 & 1'b0) | (x[31] & 1'b0 & 1'b0 & ~1'b0) | (x[31] & 1'b0 & ~1'b0 & 1'b0) | (x[31] & ~1'b0 & 1'b0 & 1'b0) | (~x[31] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[31]);
  assign t[99] = (x[34] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[34] & 1'b0 & ~1'b0 & ~1'b0) | (~x[34] & ~1'b0 & 1'b0 & ~1'b0) | (~x[34] & ~1'b0 & ~1'b0 & 1'b0) | (x[34] & 1'b0 & 1'b0 & ~1'b0) | (x[34] & 1'b0 & ~1'b0 & 1'b0) | (x[34] & ~1'b0 & 1'b0 & 1'b0) | (~x[34] & 1'b0 & 1'b0 & 1'b0);
  assign t[9] = ~(t[11] & t[12]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [21:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[30] & t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[32]);
  assign t[18] = ~(t[33]);
  assign t[19] = ~(t[30] | t[21]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[32] & t[23]);
  assign t[22] = ~(t[16] & t[24]);
  assign t[23] = ~(t[31] | t[25]);
  assign t[24] = t[26] & t[33];
  assign t[25] = ~(t[18]);
  assign t[26] = ~(t[30] | t[32]);
  assign t[27] = (t[34]);
  assign t[28] = (t[35]);
  assign t[29] = (t[36]);
  assign t[2] = t[27] ^ t[4];
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = t[41] ^ x[2];
  assign t[35] = t[42] ^ x[5];
  assign t[36] = t[43] ^ x[9];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[15];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[5]);
  assign t[40] = t[47] ^ x[21];
  assign t[41] = (~t[48] & t[49]);
  assign t[42] = (~t[50] & t[51]);
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[56] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[60] & t[61]);
  assign t[48] = t[62] ^ x[1];
  assign t[49] = t[63] ^ x[2];
  assign t[4] = ~(t[6] & t[28]);
  assign t[50] = t[64] ^ x[4];
  assign t[51] = t[65] ^ x[5];
  assign t[52] = t[66] ^ x[8];
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[12];
  assign t[56] = t[70] ^ x[14];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = t[74] ^ x[20];
  assign t[61] = t[75] ^ x[21];
  assign t[62] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[0]);
  assign t[64] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[3]);
  assign t[66] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[7]);
  assign t[68] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[10]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[13]);
  assign t[72] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[16]);
  assign t[74] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[19]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(x[6]);
  assign t[9] = ~(t[29]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind56(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind57(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind58(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind59(x, y);
 input [21:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[30] & t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[32]);
  assign t[18] = ~(t[33]);
  assign t[19] = ~(t[30] | t[21]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[32] & t[23]);
  assign t[22] = ~(t[16] & t[24]);
  assign t[23] = ~(t[31] | t[25]);
  assign t[24] = t[26] & t[33];
  assign t[25] = ~(t[18]);
  assign t[26] = ~(t[30] | t[32]);
  assign t[27] = (t[34]);
  assign t[28] = (t[35]);
  assign t[29] = (t[36]);
  assign t[2] = t[27] ^ t[4];
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = t[41] ^ x[2];
  assign t[35] = t[42] ^ x[5];
  assign t[36] = t[43] ^ x[9];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[15];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[5]);
  assign t[40] = t[47] ^ x[21];
  assign t[41] = (~t[48] & t[49]);
  assign t[42] = (~t[50] & t[51]);
  assign t[43] = (~t[52] & t[53]);
  assign t[44] = (~t[54] & t[55]);
  assign t[45] = (~t[56] & t[57]);
  assign t[46] = (~t[58] & t[59]);
  assign t[47] = (~t[60] & t[61]);
  assign t[48] = t[62] ^ x[1];
  assign t[49] = t[63] ^ x[2];
  assign t[4] = ~(t[6] & t[28]);
  assign t[50] = t[64] ^ x[4];
  assign t[51] = t[65] ^ x[5];
  assign t[52] = t[66] ^ x[8];
  assign t[53] = t[67] ^ x[9];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[12];
  assign t[56] = t[70] ^ x[14];
  assign t[57] = t[71] ^ x[15];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = t[74] ^ x[20];
  assign t[61] = t[75] ^ x[21];
  assign t[62] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[0]);
  assign t[64] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[3]);
  assign t[66] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[7]);
  assign t[68] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[10]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[13]);
  assign t[72] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[16]);
  assign t[74] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[19]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(x[6]);
  assign t[9] = ~(t[29]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [24:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(x[9]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[33] & t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~(t[29] ^ t[3]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[33] | t[23]);
  assign t[22] = ~(t[24]);
  assign t[23] = ~(t[35] & t[25]);
  assign t[24] = ~(t[18] & t[26]);
  assign t[25] = ~(t[34] | t[27]);
  assign t[26] = t[28] & t[36];
  assign t[27] = ~(t[20]);
  assign t[28] = ~(t[33] | t[35]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = t[45] ^ x[2];
  assign t[38] = t[46] ^ x[5];
  assign t[39] = t[47] ^ x[8];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[48] ^ x[12];
  assign t[41] = t[49] ^ x[15];
  assign t[42] = t[50] ^ x[18];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[24];
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = (~t[65] & t[66]);
  assign t[52] = (~t[67] & t[68]);
  assign t[53] = t[69] ^ x[1];
  assign t[54] = t[70] ^ x[2];
  assign t[55] = t[71] ^ x[4];
  assign t[56] = t[72] ^ x[5];
  assign t[57] = t[73] ^ x[7];
  assign t[58] = t[74] ^ x[8];
  assign t[59] = t[75] ^ x[11];
  assign t[5] = ~(t[30]);
  assign t[60] = t[76] ^ x[12];
  assign t[61] = t[77] ^ x[14];
  assign t[62] = t[78] ^ x[15];
  assign t[63] = t[79] ^ x[17];
  assign t[64] = t[80] ^ x[18];
  assign t[65] = t[81] ^ x[20];
  assign t[66] = t[82] ^ x[21];
  assign t[67] = t[83] ^ x[23];
  assign t[68] = t[84] ^ x[24];
  assign t[69] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[8] & t[31]);
  assign t[70] = (x[0]);
  assign t[71] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[3]);
  assign t[73] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[6]);
  assign t[75] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[10]);
  assign t[77] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[13]);
  assign t[79] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16]);
  assign t[81] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[19]);
  assign t[83] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[22]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind61(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind62(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind63(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind64(x, y);
 input [24:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(x[9]);
  assign t[11] = ~(t[32]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[33] & t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~(t[29] ^ t[3]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[33] | t[23]);
  assign t[22] = ~(t[24]);
  assign t[23] = ~(t[35] & t[25]);
  assign t[24] = ~(t[18] & t[26]);
  assign t[25] = ~(t[34] | t[27]);
  assign t[26] = t[28] & t[36];
  assign t[27] = ~(t[20]);
  assign t[28] = ~(t[33] | t[35]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = t[45] ^ x[2];
  assign t[38] = t[46] ^ x[5];
  assign t[39] = t[47] ^ x[8];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[48] ^ x[12];
  assign t[41] = t[49] ^ x[15];
  assign t[42] = t[50] ^ x[18];
  assign t[43] = t[51] ^ x[21];
  assign t[44] = t[52] ^ x[24];
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = (~t[65] & t[66]);
  assign t[52] = (~t[67] & t[68]);
  assign t[53] = t[69] ^ x[1];
  assign t[54] = t[70] ^ x[2];
  assign t[55] = t[71] ^ x[4];
  assign t[56] = t[72] ^ x[5];
  assign t[57] = t[73] ^ x[7];
  assign t[58] = t[74] ^ x[8];
  assign t[59] = t[75] ^ x[11];
  assign t[5] = ~(t[30]);
  assign t[60] = t[76] ^ x[12];
  assign t[61] = t[77] ^ x[14];
  assign t[62] = t[78] ^ x[15];
  assign t[63] = t[79] ^ x[17];
  assign t[64] = t[80] ^ x[18];
  assign t[65] = t[81] ^ x[20];
  assign t[66] = t[82] ^ x[21];
  assign t[67] = t[83] ^ x[23];
  assign t[68] = t[84] ^ x[24];
  assign t[69] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[8] & t[31]);
  assign t[70] = (x[0]);
  assign t[71] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[3]);
  assign t[73] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[6]);
  assign t[75] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[10]);
  assign t[77] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[13]);
  assign t[79] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16]);
  assign t[81] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[19]);
  assign t[83] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[22]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [18:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(x[6]);
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[28] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[28] & t[21]);
  assign t[17] = ~(t[29] & t[22]);
  assign t[18] = ~(t[19] & t[23]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[26]);
  assign t[20] = ~(t[29]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[30] | t[24]);
  assign t[23] = t[25] & t[31];
  assign t[24] = ~(t[21]);
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = (t[32]);
  assign t[27] = (t[33]);
  assign t[28] = (t[34]);
  assign t[29] = (t[35]);
  assign t[2] = ~(t[4]);
  assign t[30] = (t[36]);
  assign t[31] = (t[37]);
  assign t[32] = t[38] ^ x[2];
  assign t[33] = t[39] ^ x[5];
  assign t[34] = t[40] ^ x[9];
  assign t[35] = t[41] ^ x[12];
  assign t[36] = t[42] ^ x[15];
  assign t[37] = t[43] ^ x[18];
  assign t[38] = (~t[44] & t[45]);
  assign t[39] = (~t[46] & t[47]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (~t[48] & t[49]);
  assign t[41] = (~t[50] & t[51]);
  assign t[42] = (~t[52] & t[53]);
  assign t[43] = (~t[54] & t[55]);
  assign t[44] = t[56] ^ x[1];
  assign t[45] = t[57] ^ x[2];
  assign t[46] = t[58] ^ x[4];
  assign t[47] = t[59] ^ x[5];
  assign t[48] = t[60] ^ x[8];
  assign t[49] = t[61] ^ x[9];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ x[11];
  assign t[51] = t[63] ^ x[12];
  assign t[52] = t[64] ^ x[14];
  assign t[53] = t[65] ^ x[15];
  assign t[54] = t[66] ^ x[17];
  assign t[55] = t[67] ^ x[18];
  assign t[56] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[0]);
  assign t[58] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[3]);
  assign t[5] = ~(t[27]);
  assign t[60] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[7]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[13]);
  assign t[66] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[16]);
  assign t[6] = ~(t[8]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind66(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind67(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind68(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind69(x, y);
 input [18:0] x;
 output y;

 wire [67:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(x[6]);
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[28] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[28] & t[21]);
  assign t[17] = ~(t[29] & t[22]);
  assign t[18] = ~(t[19] & t[23]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[26]);
  assign t[20] = ~(t[29]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[30] | t[24]);
  assign t[23] = t[25] & t[31];
  assign t[24] = ~(t[21]);
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = (t[32]);
  assign t[27] = (t[33]);
  assign t[28] = (t[34]);
  assign t[29] = (t[35]);
  assign t[2] = ~(t[4]);
  assign t[30] = (t[36]);
  assign t[31] = (t[37]);
  assign t[32] = t[38] ^ x[2];
  assign t[33] = t[39] ^ x[5];
  assign t[34] = t[40] ^ x[9];
  assign t[35] = t[41] ^ x[12];
  assign t[36] = t[42] ^ x[15];
  assign t[37] = t[43] ^ x[18];
  assign t[38] = (~t[44] & t[45]);
  assign t[39] = (~t[46] & t[47]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (~t[48] & t[49]);
  assign t[41] = (~t[50] & t[51]);
  assign t[42] = (~t[52] & t[53]);
  assign t[43] = (~t[54] & t[55]);
  assign t[44] = t[56] ^ x[1];
  assign t[45] = t[57] ^ x[2];
  assign t[46] = t[58] ^ x[4];
  assign t[47] = t[59] ^ x[5];
  assign t[48] = t[60] ^ x[8];
  assign t[49] = t[61] ^ x[9];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ x[11];
  assign t[51] = t[63] ^ x[12];
  assign t[52] = t[64] ^ x[14];
  assign t[53] = t[65] ^ x[15];
  assign t[54] = t[66] ^ x[17];
  assign t[55] = t[67] ^ x[18];
  assign t[56] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[0]);
  assign t[58] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[3]);
  assign t[5] = ~(t[27]);
  assign t[60] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[7]);
  assign t[62] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[10]);
  assign t[64] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[13]);
  assign t[66] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[16]);
  assign t[6] = ~(t[8]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[12]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [15:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[25] | t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[26] & t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[18] & t[20]);
  assign t[16] = ~(t[25] & t[21]);
  assign t[17] = ~(t[27] | t[22]);
  assign t[18] = ~(t[27]);
  assign t[19] = t[23] & t[28];
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[26]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[21]);
  assign t[23] = ~(t[25] | t[26]);
  assign t[24] = (t[29]);
  assign t[25] = (t[30]);
  assign t[26] = (t[31]);
  assign t[27] = (t[32]);
  assign t[28] = (t[33]);
  assign t[29] = t[34] ^ x[2];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[9];
  assign t[32] = t[37] ^ x[12];
  assign t[33] = t[38] ^ x[15];
  assign t[34] = (~t[39] & t[40]);
  assign t[35] = (~t[41] & t[42]);
  assign t[36] = (~t[43] & t[44]);
  assign t[37] = (~t[45] & t[46]);
  assign t[38] = (~t[47] & t[48]);
  assign t[39] = t[49] ^ x[1];
  assign t[3] = ~(t[6]);
  assign t[40] = t[50] ^ x[2];
  assign t[41] = t[51] ^ x[5];
  assign t[42] = t[52] ^ x[6];
  assign t[43] = t[53] ^ x[8];
  assign t[44] = t[54] ^ x[9];
  assign t[45] = t[55] ^ x[11];
  assign t[46] = t[56] ^ x[12];
  assign t[47] = t[57] ^ x[14];
  assign t[48] = t[58] ^ x[15];
  assign t[49] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[24]);
  assign t[50] = (x[0]);
  assign t[51] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[4]);
  assign t[53] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[7]);
  assign t[55] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[10]);
  assign t[57] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[13]);
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(x[3]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind71(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind72(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind73(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind74(x, y);
 input [15:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[25] | t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[26] & t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[18] & t[20]);
  assign t[16] = ~(t[25] & t[21]);
  assign t[17] = ~(t[27] | t[22]);
  assign t[18] = ~(t[27]);
  assign t[19] = t[23] & t[28];
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[26]);
  assign t[21] = ~(t[28]);
  assign t[22] = ~(t[21]);
  assign t[23] = ~(t[25] | t[26]);
  assign t[24] = (t[29]);
  assign t[25] = (t[30]);
  assign t[26] = (t[31]);
  assign t[27] = (t[32]);
  assign t[28] = (t[33]);
  assign t[29] = t[34] ^ x[2];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[9];
  assign t[32] = t[37] ^ x[12];
  assign t[33] = t[38] ^ x[15];
  assign t[34] = (~t[39] & t[40]);
  assign t[35] = (~t[41] & t[42]);
  assign t[36] = (~t[43] & t[44]);
  assign t[37] = (~t[45] & t[46]);
  assign t[38] = (~t[47] & t[48]);
  assign t[39] = t[49] ^ x[1];
  assign t[3] = ~(t[6]);
  assign t[40] = t[50] ^ x[2];
  assign t[41] = t[51] ^ x[5];
  assign t[42] = t[52] ^ x[6];
  assign t[43] = t[53] ^ x[8];
  assign t[44] = t[54] ^ x[9];
  assign t[45] = t[55] ^ x[11];
  assign t[46] = t[56] ^ x[12];
  assign t[47] = t[57] ^ x[14];
  assign t[48] = t[58] ^ x[15];
  assign t[49] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[24]);
  assign t[50] = (x[0]);
  assign t[51] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[52] = (x[4]);
  assign t[53] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[54] = (x[7]);
  assign t[55] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[56] = (x[10]);
  assign t[57] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[13]);
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(x[3]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [69:0] x;
 output y;

 wire [216:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (t[122]);
  assign t[101] = (t[123]);
  assign t[102] = (t[124]);
  assign t[103] = (t[125]);
  assign t[104] = (t[126]);
  assign t[105] = (t[127]);
  assign t[106] = (t[128]);
  assign t[107] = t[129] ^ x[5];
  assign t[108] = t[130] ^ x[9];
  assign t[109] = t[131] ^ x[15];
  assign t[10] = ~(t[17] & t[18]);
  assign t[110] = t[132] ^ x[21];
  assign t[111] = t[133] ^ x[25];
  assign t[112] = t[134] ^ x[28];
  assign t[113] = t[135] ^ x[34];
  assign t[114] = t[136] ^ x[35];
  assign t[115] = t[137] ^ x[36];
  assign t[116] = t[138] ^ x[39];
  assign t[117] = t[139] ^ x[40];
  assign t[118] = t[140] ^ x[41];
  assign t[119] = t[141] ^ x[42];
  assign t[11] = t[19] ? x[6] : t[85];
  assign t[120] = t[142] ^ x[43];
  assign t[121] = t[143] ^ x[44];
  assign t[122] = t[144] ^ x[45];
  assign t[123] = t[145] ^ x[46];
  assign t[124] = t[146] ^ x[52];
  assign t[125] = t[147] ^ x[54];
  assign t[126] = t[148] ^ x[60];
  assign t[127] = t[149] ^ x[62];
  assign t[128] = t[150] ^ x[68];
  assign t[129] = (~t[151] & t[152]);
  assign t[12] = ~(t[3]);
  assign t[130] = (~t[153] & t[154]);
  assign t[131] = (~t[155] & t[156]);
  assign t[132] = (~t[157] & t[158]);
  assign t[133] = (~t[159] & t[160]);
  assign t[134] = (~t[161] & t[162]);
  assign t[135] = (~t[163] & t[164]);
  assign t[136] = (~t[163] & t[165]);
  assign t[137] = (~t[155] & t[166]);
  assign t[138] = (~t[167] & t[168]);
  assign t[139] = (~t[163] & t[169]);
  assign t[13] = ~(t[86] | t[20]);
  assign t[140] = (~t[155] & t[170]);
  assign t[141] = (~t[157] & t[171]);
  assign t[142] = (~t[157] & t[172]);
  assign t[143] = (~t[155] & t[173]);
  assign t[144] = (~t[157] & t[174]);
  assign t[145] = (~t[151] & t[175]);
  assign t[146] = (~t[176] & t[177]);
  assign t[147] = (~t[151] & t[178]);
  assign t[148] = (~t[179] & t[180]);
  assign t[149] = (~t[151] & t[181]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = (~t[182] & t[183]);
  assign t[151] = t[184] ^ x[4];
  assign t[152] = t[185] ^ x[5];
  assign t[153] = t[186] ^ x[8];
  assign t[154] = t[187] ^ x[9];
  assign t[155] = t[188] ^ x[14];
  assign t[156] = t[189] ^ x[15];
  assign t[157] = t[190] ^ x[20];
  assign t[158] = t[191] ^ x[21];
  assign t[159] = t[192] ^ x[24];
  assign t[15] = t[87] ^ t[88];
  assign t[160] = t[193] ^ x[25];
  assign t[161] = t[194] ^ x[27];
  assign t[162] = t[195] ^ x[28];
  assign t[163] = t[196] ^ x[33];
  assign t[164] = t[197] ^ x[34];
  assign t[165] = t[198] ^ x[35];
  assign t[166] = t[199] ^ x[36];
  assign t[167] = t[200] ^ x[38];
  assign t[168] = t[201] ^ x[39];
  assign t[169] = t[202] ^ x[40];
  assign t[16] = ~(t[23]);
  assign t[170] = t[203] ^ x[41];
  assign t[171] = t[204] ^ x[42];
  assign t[172] = t[205] ^ x[43];
  assign t[173] = t[206] ^ x[44];
  assign t[174] = t[207] ^ x[45];
  assign t[175] = t[208] ^ x[46];
  assign t[176] = t[209] ^ x[51];
  assign t[177] = t[210] ^ x[52];
  assign t[178] = t[211] ^ x[54];
  assign t[179] = t[212] ^ x[59];
  assign t[17] = ~(t[24]);
  assign t[180] = t[213] ^ x[60];
  assign t[181] = t[214] ^ x[62];
  assign t[182] = t[215] ^ x[67];
  assign t[183] = t[216] ^ x[68];
  assign t[184] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[185] = (x[0]);
  assign t[186] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[187] = (x[7]);
  assign t[188] = (x[10] & ~x[11] & ~x[12] & ~x[13]) | (~x[10] & x[11] & ~x[12] & ~x[13]) | (~x[10] & ~x[11] & x[12] & ~x[13]) | (~x[10] & ~x[11] & ~x[12] & x[13]) | (x[10] & x[11] & x[12] & ~x[13]) | (x[10] & x[11] & ~x[12] & x[13]) | (x[10] & ~x[11] & x[12] & x[13]) | (~x[10] & x[11] & x[12] & x[13]);
  assign t[189] = (x[13]);
  assign t[18] = ~(x[22]);
  assign t[190] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[191] = (x[19]);
  assign t[192] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[193] = (x[23]);
  assign t[194] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[195] = (x[26]);
  assign t[196] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[197] = (x[32]);
  assign t[198] = (x[30]);
  assign t[199] = (x[10]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[201] = (x[37]);
  assign t[202] = (x[31]);
  assign t[203] = (x[12]);
  assign t[204] = (x[18]);
  assign t[205] = (x[16]);
  assign t[206] = (x[11]);
  assign t[207] = (x[17]);
  assign t[208] = (x[1]);
  assign t[209] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[20] = ~(t[89] & t[26]);
  assign t[210] = (x[50]);
  assign t[211] = (x[2]);
  assign t[212] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[213] = (x[58]);
  assign t[214] = (x[3]);
  assign t[215] = (x[63] & ~x[64] & ~x[65] & ~x[66]) | (~x[63] & x[64] & ~x[65] & ~x[66]) | (~x[63] & ~x[64] & x[65] & ~x[66]) | (~x[63] & ~x[64] & ~x[65] & x[66]) | (x[63] & x[64] & x[65] & ~x[66]) | (x[63] & x[64] & ~x[65] & x[66]) | (x[63] & ~x[64] & x[65] & x[66]) | (~x[63] & x[64] & x[65] & x[66]);
  assign t[216] = (x[66]);
  assign t[21] = ~(t[27] | t[28]);
  assign t[22] = ~(t[29] ^ t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = ~(t[33] | t[34]);
  assign t[25] = ~(x[22]);
  assign t[26] = ~(t[90] | t[35]);
  assign t[27] = ~(t[36]);
  assign t[28] = t[24] ? t[91] : t[37];
  assign t[29] = t[24] ? t[92] : t[38];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[24] ? t[93] : t[15];
  assign t[31] = ~(t[90]);
  assign t[32] = t[39] & t[94];
  assign t[33] = ~(t[31] & t[40]);
  assign t[34] = ~(t[86] & t[41]);
  assign t[35] = ~(t[41]);
  assign t[36] = t[24] ? t[95] : t[42];
  assign t[37] = t[96] ^ t[97];
  assign t[38] = t[93] ^ t[98];
  assign t[39] = ~(t[86] | t[89]);
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = ~(t[89]);
  assign t[41] = ~(t[94]);
  assign t[42] = t[99] ^ t[100];
  assign t[43] = ~(t[44] & t[45]);
  assign t[44] = t[3] ? t[47] : t[46];
  assign t[45] = ~(t[6] & t[48]);
  assign t[46] = ~(t[101]);
  assign t[47] = ~(t[10] & t[49]);
  assign t[48] = t[13] ? t[37] : t[50];
  assign t[49] = t[19] ? x[53] : t[102];
  assign t[4] = ~(t[85]);
  assign t[50] = ~(t[51] | t[52]);
  assign t[51] = ~(t[53] | t[54]);
  assign t[52] = ~(t[27] | t[22]);
  assign t[53] = ~(t[55] | t[27]);
  assign t[54] = t[29] ? t[56] : t[28];
  assign t[55] = ~(t[29] | t[30]);
  assign t[56] = ~(t[28] & t[57]);
  assign t[57] = ~(t[58] & t[27]);
  assign t[58] = ~(t[30]);
  assign t[59] = ~(t[60] & t[61]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = t[3] ? t[63] : t[62];
  assign t[61] = ~(t[6] & t[64]);
  assign t[62] = ~(t[103]);
  assign t[63] = ~(t[10] & t[65]);
  assign t[64] = t[13] ? t[42] : t[66];
  assign t[65] = t[19] ? x[61] : t[104];
  assign t[66] = ~(t[67] & t[68]);
  assign t[67] = ~(t[69] & t[56]);
  assign t[68] = ~(t[53] & t[54]);
  assign t[69] = ~(t[36] | t[70]);
  assign t[6] = ~(t[10] | t[12]);
  assign t[70] = ~(t[71] | t[72]);
  assign t[71] = ~(t[29]);
  assign t[72] = ~(t[58] & t[73]);
  assign t[73] = ~(t[28]);
  assign t[74] = ~(t[75] & t[76]);
  assign t[75] = t[3] ? t[78] : t[77];
  assign t[76] = ~(t[6] & t[79]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[10] & t[80]);
  assign t[79] = t[13] ? t[38] : t[81];
  assign t[7] = t[13] ? t[15] : t[14];
  assign t[80] = t[19] ? x[69] : t[106];
  assign t[81] = ~(t[82] & t[83]);
  assign t[82] = t[29] ? t[84] : t[56];
  assign t[83] = ~(t[55] & t[73]);
  assign t[84] = ~(t[27] & t[72]);
  assign t[85] = (t[107]);
  assign t[86] = (t[108]);
  assign t[87] = (t[109]);
  assign t[88] = (t[110]);
  assign t[89] = (t[111]);
  assign t[8] = ~(t[13] | t[16]);
  assign t[90] = (t[112]);
  assign t[91] = (t[113]);
  assign t[92] = (t[114]);
  assign t[93] = (t[115]);
  assign t[94] = (t[116]);
  assign t[95] = (t[117]);
  assign t[96] = (t[118]);
  assign t[97] = (t[119]);
  assign t[98] = (t[120]);
  assign t[99] = (t[121]);
  assign t[9] = ~(t[10]);
  assign y = (t[0] & ~t[43] & ~t[59] & ~t[74]) | (~t[0] & t[43] & ~t[59] & ~t[74]) | (~t[0] & ~t[43] & t[59] & ~t[74]) | (~t[0] & ~t[43] & ~t[59] & t[74]) | (t[0] & t[43] & t[59] & ~t[74]) | (t[0] & t[43] & ~t[59] & t[74]) | (t[0] & ~t[43] & t[59] & t[74]) | (~t[0] & t[43] & t[59] & t[74]);
endmodule

module R2ind76(x, y);
 input [51:0] x;
 output y;

 wire [152:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (~t[109] & t[126]);
  assign t[101] = t[127] ^ x[4];
  assign t[102] = t[128] ^ x[5];
  assign t[103] = t[129] ^ x[10];
  assign t[104] = t[130] ^ x[11];
  assign t[105] = t[131] ^ x[14];
  assign t[106] = t[132] ^ x[15];
  assign t[107] = t[133] ^ x[20];
  assign t[108] = t[134] ^ x[21];
  assign t[109] = t[135] ^ x[26];
  assign t[10] = ~(t[17] & t[18]);
  assign t[110] = t[136] ^ x[27];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[33];
  assign t[114] = t[140] ^ x[34];
  assign t[115] = t[141] ^ x[39];
  assign t[116] = t[142] ^ x[40];
  assign t[117] = t[143] ^ x[42];
  assign t[118] = t[144] ^ x[43];
  assign t[119] = t[145] ^ x[44];
  assign t[11] = t[19] ? x[12] : t[51];
  assign t[120] = t[146] ^ x[45];
  assign t[121] = t[147] ^ x[46];
  assign t[122] = t[148] ^ x[47];
  assign t[123] = t[149] ^ x[48];
  assign t[124] = t[150] ^ x[49];
  assign t[125] = t[151] ^ x[50];
  assign t[126] = t[152] ^ x[51];
  assign t[127] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[128] = (x[3]);
  assign t[129] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[12] = ~(t[3]);
  assign t[130] = (x[9]);
  assign t[131] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[13]);
  assign t[133] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[134] = (x[16]);
  assign t[135] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[136] = (x[22]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[13] = ~(t[52] | t[20]);
  assign t[140] = (x[32]);
  assign t[141] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[142] = (x[36]);
  assign t[143] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[144] = (x[41]);
  assign t[145] = (x[38]);
  assign t[146] = (x[18]);
  assign t[147] = (x[24]);
  assign t[148] = (x[37]);
  assign t[149] = (x[19]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[150] = (x[25]);
  assign t[151] = (x[17]);
  assign t[152] = (x[23]);
  assign t[15] = t[53] ^ t[54];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(x[28]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[55] & t[26]);
  assign t[21] = t[27] ? t[29] : t[28];
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(x[28]);
  assign t[26] = ~(t[56] | t[36]);
  assign t[27] = t[24] ? t[57] : t[15];
  assign t[28] = ~(t[37] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[27] | t[41]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[56]);
  assign t[33] = t[42] & t[58];
  assign t[34] = ~(t[32] & t[43]);
  assign t[35] = ~(t[52] & t[44]);
  assign t[36] = ~(t[44]);
  assign t[37] = t[24] ? t[59] : t[45];
  assign t[38] = ~(t[46] & t[39]);
  assign t[39] = ~(t[47]);
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = ~(t[46] & t[31]);
  assign t[41] = t[24] ? t[53] : t[48];
  assign t[42] = ~(t[52] | t[55]);
  assign t[43] = ~(t[55]);
  assign t[44] = ~(t[58]);
  assign t[45] = t[60] ^ t[61];
  assign t[46] = ~(t[41]);
  assign t[47] = t[24] ? t[62] : t[49];
  assign t[48] = t[63] ^ t[64];
  assign t[49] = t[65] ^ t[66];
  assign t[4] = ~(t[50]);
  assign t[50] = (t[67]);
  assign t[51] = (t[68]);
  assign t[52] = (t[69]);
  assign t[53] = (t[70]);
  assign t[54] = (t[71]);
  assign t[55] = (t[72]);
  assign t[56] = (t[73]);
  assign t[57] = (t[74]);
  assign t[58] = (t[75]);
  assign t[59] = (t[76]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (t[77]);
  assign t[61] = (t[78]);
  assign t[62] = (t[79]);
  assign t[63] = (t[80]);
  assign t[64] = (t[81]);
  assign t[65] = (t[82]);
  assign t[66] = (t[83]);
  assign t[67] = t[84] ^ x[5];
  assign t[68] = t[85] ^ x[11];
  assign t[69] = t[86] ^ x[15];
  assign t[6] = ~(t[10] | t[12]);
  assign t[70] = t[87] ^ x[21];
  assign t[71] = t[88] ^ x[27];
  assign t[72] = t[89] ^ x[31];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[40];
  assign t[75] = t[92] ^ x[43];
  assign t[76] = t[93] ^ x[44];
  assign t[77] = t[94] ^ x[45];
  assign t[78] = t[95] ^ x[46];
  assign t[79] = t[96] ^ x[47];
  assign t[7] = t[13] ? t[15] : t[14];
  assign t[80] = t[97] ^ x[48];
  assign t[81] = t[98] ^ x[49];
  assign t[82] = t[99] ^ x[50];
  assign t[83] = t[100] ^ x[51];
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[13] | t[16]);
  assign t[90] = (~t[113] & t[114]);
  assign t[91] = (~t[115] & t[116]);
  assign t[92] = (~t[117] & t[118]);
  assign t[93] = (~t[115] & t[119]);
  assign t[94] = (~t[107] & t[120]);
  assign t[95] = (~t[109] & t[121]);
  assign t[96] = (~t[115] & t[122]);
  assign t[97] = (~t[107] & t[123]);
  assign t[98] = (~t[109] & t[124]);
  assign t[99] = (~t[107] & t[125]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [51:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (~t[113] & t[126]);
  assign t[101] = (~t[111] & t[127]);
  assign t[102] = (~t[113] & t[128]);
  assign t[103] = (~t[111] & t[129]);
  assign t[104] = (~t[113] & t[130]);
  assign t[105] = t[131] ^ x[4];
  assign t[106] = t[132] ^ x[5];
  assign t[107] = t[133] ^ x[10];
  assign t[108] = t[134] ^ x[11];
  assign t[109] = t[135] ^ x[14];
  assign t[10] = ~(t[17] & t[18]);
  assign t[110] = t[136] ^ x[15];
  assign t[111] = t[137] ^ x[20];
  assign t[112] = t[138] ^ x[21];
  assign t[113] = t[139] ^ x[26];
  assign t[114] = t[140] ^ x[27];
  assign t[115] = t[141] ^ x[30];
  assign t[116] = t[142] ^ x[31];
  assign t[117] = t[143] ^ x[33];
  assign t[118] = t[144] ^ x[34];
  assign t[119] = t[145] ^ x[36];
  assign t[11] = t[19] ? x[12] : t[55];
  assign t[120] = t[146] ^ x[37];
  assign t[121] = t[147] ^ x[42];
  assign t[122] = t[148] ^ x[43];
  assign t[123] = t[149] ^ x[44];
  assign t[124] = t[150] ^ x[45];
  assign t[125] = t[151] ^ x[46];
  assign t[126] = t[152] ^ x[47];
  assign t[127] = t[153] ^ x[48];
  assign t[128] = t[154] ^ x[49];
  assign t[129] = t[155] ^ x[50];
  assign t[12] = ~(t[3]);
  assign t[130] = t[156] ^ x[51];
  assign t[131] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[132] = (x[2]);
  assign t[133] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[134] = (x[9]);
  assign t[135] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[13]);
  assign t[137] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[138] = (x[17]);
  assign t[139] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[13] = ~(t[56] | t[20]);
  assign t[140] = (x[23]);
  assign t[141] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[142] = (x[29]);
  assign t[143] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[144] = (x[32]);
  assign t[145] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[146] = (x[35]);
  assign t[147] = (x[38] & ~x[39] & ~x[40] & ~x[41]) | (~x[38] & x[39] & ~x[40] & ~x[41]) | (~x[38] & ~x[39] & x[40] & ~x[41]) | (~x[38] & ~x[39] & ~x[40] & x[41]) | (x[38] & x[39] & x[40] & ~x[41]) | (x[38] & x[39] & ~x[40] & x[41]) | (x[38] & ~x[39] & x[40] & x[41]) | (~x[38] & x[39] & x[40] & x[41]);
  assign t[148] = (x[40]);
  assign t[149] = (x[41]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[150] = (x[39]);
  assign t[151] = (x[18]);
  assign t[152] = (x[24]);
  assign t[153] = (x[16]);
  assign t[154] = (x[22]);
  assign t[155] = (x[19]);
  assign t[156] = (x[25]);
  assign t[15] = t[57] ^ t[58];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(x[28]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[59] & t[26]);
  assign t[21] = ~(t[27] & t[28]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = ~(t[33] | t[34]);
  assign t[25] = ~(x[28]);
  assign t[26] = ~(t[60] | t[35]);
  assign t[27] = ~(t[36] | t[37]);
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = ~(t[40] | t[41]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[42] ? t[28] : t[38];
  assign t[31] = ~(t[60]);
  assign t[32] = t[43] & t[61];
  assign t[33] = ~(t[31] & t[44]);
  assign t[34] = ~(t[56] & t[45]);
  assign t[35] = ~(t[45]);
  assign t[36] = t[24] ? t[62] : t[15];
  assign t[37] = ~(t[46] | t[47]);
  assign t[38] = t[24] ? t[63] : t[48];
  assign t[39] = ~(t[49] & t[41]);
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = ~(t[42] | t[50]);
  assign t[41] = ~(t[36]);
  assign t[42] = t[24] ? t[64] : t[51];
  assign t[43] = ~(t[56] | t[59]);
  assign t[44] = ~(t[59]);
  assign t[45] = ~(t[61]);
  assign t[46] = ~(t[42]);
  assign t[47] = ~(t[49] & t[52]);
  assign t[48] = t[65] ^ t[66];
  assign t[49] = ~(t[50]);
  assign t[4] = ~(t[54]);
  assign t[50] = t[24] ? t[67] : t[53];
  assign t[51] = t[67] ^ t[68];
  assign t[52] = ~(t[38]);
  assign t[53] = t[69] ^ t[70];
  assign t[54] = (t[71]);
  assign t[55] = (t[72]);
  assign t[56] = (t[73]);
  assign t[57] = (t[74]);
  assign t[58] = (t[75]);
  assign t[59] = (t[76]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (t[77]);
  assign t[61] = (t[78]);
  assign t[62] = (t[79]);
  assign t[63] = (t[80]);
  assign t[64] = (t[81]);
  assign t[65] = (t[82]);
  assign t[66] = (t[83]);
  assign t[67] = (t[84]);
  assign t[68] = (t[85]);
  assign t[69] = (t[86]);
  assign t[6] = ~(t[10] | t[12]);
  assign t[70] = (t[87]);
  assign t[71] = t[88] ^ x[5];
  assign t[72] = t[89] ^ x[11];
  assign t[73] = t[90] ^ x[15];
  assign t[74] = t[91] ^ x[21];
  assign t[75] = t[92] ^ x[27];
  assign t[76] = t[93] ^ x[31];
  assign t[77] = t[94] ^ x[34];
  assign t[78] = t[95] ^ x[37];
  assign t[79] = t[96] ^ x[43];
  assign t[7] = t[13] ? t[15] : t[14];
  assign t[80] = t[97] ^ x[44];
  assign t[81] = t[98] ^ x[45];
  assign t[82] = t[99] ^ x[46];
  assign t[83] = t[100] ^ x[47];
  assign t[84] = t[101] ^ x[48];
  assign t[85] = t[102] ^ x[49];
  assign t[86] = t[103] ^ x[50];
  assign t[87] = t[104] ^ x[51];
  assign t[88] = (~t[105] & t[106]);
  assign t[89] = (~t[107] & t[108]);
  assign t[8] = ~(t[13] | t[16]);
  assign t[90] = (~t[109] & t[110]);
  assign t[91] = (~t[111] & t[112]);
  assign t[92] = (~t[113] & t[114]);
  assign t[93] = (~t[115] & t[116]);
  assign t[94] = (~t[117] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[121] & t[122]);
  assign t[97] = (~t[121] & t[123]);
  assign t[98] = (~t[121] & t[124]);
  assign t[99] = (~t[111] & t[125]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [51:0] x;
 output y;

 wire [152:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (~t[109] & t[126]);
  assign t[101] = t[127] ^ x[4];
  assign t[102] = t[128] ^ x[5];
  assign t[103] = t[129] ^ x[10];
  assign t[104] = t[130] ^ x[11];
  assign t[105] = t[131] ^ x[14];
  assign t[106] = t[132] ^ x[15];
  assign t[107] = t[133] ^ x[20];
  assign t[108] = t[134] ^ x[21];
  assign t[109] = t[135] ^ x[26];
  assign t[10] = ~(t[17] & t[18]);
  assign t[110] = t[136] ^ x[27];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[33];
  assign t[114] = t[140] ^ x[34];
  assign t[115] = t[141] ^ x[36];
  assign t[116] = t[142] ^ x[37];
  assign t[117] = t[143] ^ x[42];
  assign t[118] = t[144] ^ x[43];
  assign t[119] = t[145] ^ x[44];
  assign t[11] = t[19] ? x[12] : t[51];
  assign t[120] = t[146] ^ x[45];
  assign t[121] = t[147] ^ x[46];
  assign t[122] = t[148] ^ x[47];
  assign t[123] = t[149] ^ x[48];
  assign t[124] = t[150] ^ x[49];
  assign t[125] = t[151] ^ x[50];
  assign t[126] = t[152] ^ x[51];
  assign t[127] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[128] = (x[1]);
  assign t[129] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[12] = ~(t[3]);
  assign t[130] = (x[9]);
  assign t[131] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[13]);
  assign t[133] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[134] = (x[18]);
  assign t[135] = (x[22] & ~x[23] & ~x[24] & ~x[25]) | (~x[22] & x[23] & ~x[24] & ~x[25]) | (~x[22] & ~x[23] & x[24] & ~x[25]) | (~x[22] & ~x[23] & ~x[24] & x[25]) | (x[22] & x[23] & x[24] & ~x[25]) | (x[22] & x[23] & ~x[24] & x[25]) | (x[22] & ~x[23] & x[24] & x[25]) | (~x[22] & x[23] & x[24] & x[25]);
  assign t[136] = (x[24]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[13] = ~(t[52] | t[20]);
  assign t[140] = (x[32]);
  assign t[141] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[142] = (x[35]);
  assign t[143] = (x[38] & ~x[39] & ~x[40] & ~x[41]) | (~x[38] & x[39] & ~x[40] & ~x[41]) | (~x[38] & ~x[39] & x[40] & ~x[41]) | (~x[38] & ~x[39] & ~x[40] & x[41]) | (x[38] & x[39] & x[40] & ~x[41]) | (x[38] & x[39] & ~x[40] & x[41]) | (x[38] & ~x[39] & x[40] & x[41]) | (~x[38] & x[39] & x[40] & x[41]);
  assign t[144] = (x[39]);
  assign t[145] = (x[41]);
  assign t[146] = (x[40]);
  assign t[147] = (x[16]);
  assign t[148] = (x[22]);
  assign t[149] = (x[17]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[150] = (x[23]);
  assign t[151] = (x[19]);
  assign t[152] = (x[25]);
  assign t[15] = t[53] ^ t[54];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(x[28]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[55] & t[26]);
  assign t[21] = ~(t[27] | t[28]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = ~(t[33] | t[34]);
  assign t[25] = ~(x[28]);
  assign t[26] = ~(t[56] | t[35]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[37] ? t[39] : t[38];
  assign t[29] = ~(t[40]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = ~(t[37] ^ t[41]);
  assign t[31] = ~(t[56]);
  assign t[32] = t[42] & t[57];
  assign t[33] = ~(t[31] & t[43]);
  assign t[34] = ~(t[52] & t[44]);
  assign t[35] = ~(t[44]);
  assign t[36] = ~(t[37] | t[41]);
  assign t[37] = t[24] ? t[58] : t[45];
  assign t[38] = t[24] ? t[59] : t[15];
  assign t[39] = ~(t[38] & t[46]);
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = t[24] ? t[60] : t[47];
  assign t[41] = t[24] ? t[61] : t[48];
  assign t[42] = ~(t[52] | t[55]);
  assign t[43] = ~(t[55]);
  assign t[44] = ~(t[57]);
  assign t[45] = t[61] ^ t[62];
  assign t[46] = ~(t[49] & t[29]);
  assign t[47] = t[63] ^ t[64];
  assign t[48] = t[65] ^ t[66];
  assign t[49] = ~(t[41]);
  assign t[4] = ~(t[50]);
  assign t[50] = (t[67]);
  assign t[51] = (t[68]);
  assign t[52] = (t[69]);
  assign t[53] = (t[70]);
  assign t[54] = (t[71]);
  assign t[55] = (t[72]);
  assign t[56] = (t[73]);
  assign t[57] = (t[74]);
  assign t[58] = (t[75]);
  assign t[59] = (t[76]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = (t[77]);
  assign t[61] = (t[78]);
  assign t[62] = (t[79]);
  assign t[63] = (t[80]);
  assign t[64] = (t[81]);
  assign t[65] = (t[82]);
  assign t[66] = (t[83]);
  assign t[67] = t[84] ^ x[5];
  assign t[68] = t[85] ^ x[11];
  assign t[69] = t[86] ^ x[15];
  assign t[6] = ~(t[10] | t[12]);
  assign t[70] = t[87] ^ x[21];
  assign t[71] = t[88] ^ x[27];
  assign t[72] = t[89] ^ x[31];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[37];
  assign t[75] = t[92] ^ x[43];
  assign t[76] = t[93] ^ x[44];
  assign t[77] = t[94] ^ x[45];
  assign t[78] = t[95] ^ x[46];
  assign t[79] = t[96] ^ x[47];
  assign t[7] = t[13] ? t[15] : t[14];
  assign t[80] = t[97] ^ x[48];
  assign t[81] = t[98] ^ x[49];
  assign t[82] = t[99] ^ x[50];
  assign t[83] = t[100] ^ x[51];
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[13] | t[16]);
  assign t[90] = (~t[113] & t[114]);
  assign t[91] = (~t[115] & t[116]);
  assign t[92] = (~t[117] & t[118]);
  assign t[93] = (~t[117] & t[119]);
  assign t[94] = (~t[117] & t[120]);
  assign t[95] = (~t[107] & t[121]);
  assign t[96] = (~t[109] & t[122]);
  assign t[97] = (~t[107] & t[123]);
  assign t[98] = (~t[109] & t[124]);
  assign t[99] = (~t[107] & t[125]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [45:0] x;
 output y;

 wire [138:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[124] ^ x[25];
  assign t[101] = t[125] ^ x[27];
  assign t[102] = t[126] ^ x[28];
  assign t[103] = t[127] ^ x[33];
  assign t[104] = t[128] ^ x[34];
  assign t[105] = t[129] ^ x[35];
  assign t[106] = t[130] ^ x[36];
  assign t[107] = t[131] ^ x[38];
  assign t[108] = t[132] ^ x[39];
  assign t[109] = t[133] ^ x[40];
  assign t[10] = ~(t[17] & t[18]);
  assign t[110] = t[134] ^ x[41];
  assign t[111] = t[135] ^ x[42];
  assign t[112] = t[136] ^ x[43];
  assign t[113] = t[137] ^ x[44];
  assign t[114] = t[138] ^ x[45];
  assign t[115] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[116] = (x[0]);
  assign t[117] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[7]);
  assign t[119] = (x[10] & ~x[11] & ~x[12] & ~x[13]) | (~x[10] & x[11] & ~x[12] & ~x[13]) | (~x[10] & ~x[11] & x[12] & ~x[13]) | (~x[10] & ~x[11] & ~x[12] & x[13]) | (x[10] & x[11] & x[12] & ~x[13]) | (x[10] & x[11] & ~x[12] & x[13]) | (x[10] & ~x[11] & x[12] & x[13]) | (~x[10] & x[11] & x[12] & x[13]);
  assign t[11] = t[19] ? x[6] : t[43];
  assign t[120] = (x[13]);
  assign t[121] = (x[16] & ~x[17] & ~x[18] & ~x[19]) | (~x[16] & x[17] & ~x[18] & ~x[19]) | (~x[16] & ~x[17] & x[18] & ~x[19]) | (~x[16] & ~x[17] & ~x[18] & x[19]) | (x[16] & x[17] & x[18] & ~x[19]) | (x[16] & x[17] & ~x[18] & x[19]) | (x[16] & ~x[17] & x[18] & x[19]) | (~x[16] & x[17] & x[18] & x[19]);
  assign t[122] = (x[19]);
  assign t[123] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[23]);
  assign t[125] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[26]);
  assign t[127] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[128] = (x[32]);
  assign t[129] = (x[30]);
  assign t[12] = ~(t[3]);
  assign t[130] = (x[10]);
  assign t[131] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[37]);
  assign t[133] = (x[31]);
  assign t[134] = (x[12]);
  assign t[135] = (x[18]);
  assign t[136] = (x[16]);
  assign t[137] = (x[11]);
  assign t[138] = (x[17]);
  assign t[13] = ~(t[44] | t[20]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = t[45] ^ t[46];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(x[22]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[47] & t[26]);
  assign t[21] = ~(t[27] | t[28]);
  assign t[22] = ~(t[29] ^ t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = ~(t[33] | t[34]);
  assign t[25] = ~(x[22]);
  assign t[26] = ~(t[48] | t[35]);
  assign t[27] = ~(t[36]);
  assign t[28] = t[24] ? t[49] : t[37];
  assign t[29] = t[24] ? t[50] : t[38];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[24] ? t[51] : t[15];
  assign t[31] = ~(t[48]);
  assign t[32] = t[39] & t[52];
  assign t[33] = ~(t[31] & t[40]);
  assign t[34] = ~(t[44] & t[41]);
  assign t[35] = ~(t[41]);
  assign t[36] = t[24] ? t[53] : t[42];
  assign t[37] = t[54] ^ t[55];
  assign t[38] = t[51] ^ t[56];
  assign t[39] = ~(t[44] | t[47]);
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = ~(t[47]);
  assign t[41] = ~(t[52]);
  assign t[42] = t[57] ^ t[58];
  assign t[43] = (t[59]);
  assign t[44] = (t[60]);
  assign t[45] = (t[61]);
  assign t[46] = (t[62]);
  assign t[47] = (t[63]);
  assign t[48] = (t[64]);
  assign t[49] = (t[65]);
  assign t[4] = ~(t[43]);
  assign t[50] = (t[66]);
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = t[75] ^ x[5];
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = t[76] ^ x[9];
  assign t[61] = t[77] ^ x[15];
  assign t[62] = t[78] ^ x[21];
  assign t[63] = t[79] ^ x[25];
  assign t[64] = t[80] ^ x[28];
  assign t[65] = t[81] ^ x[34];
  assign t[66] = t[82] ^ x[35];
  assign t[67] = t[83] ^ x[36];
  assign t[68] = t[84] ^ x[39];
  assign t[69] = t[85] ^ x[40];
  assign t[6] = ~(t[10] | t[12]);
  assign t[70] = t[86] ^ x[41];
  assign t[71] = t[87] ^ x[42];
  assign t[72] = t[88] ^ x[43];
  assign t[73] = t[89] ^ x[44];
  assign t[74] = t[90] ^ x[45];
  assign t[75] = (~t[91] & t[92]);
  assign t[76] = (~t[93] & t[94]);
  assign t[77] = (~t[95] & t[96]);
  assign t[78] = (~t[97] & t[98]);
  assign t[79] = (~t[99] & t[100]);
  assign t[7] = t[13] ? t[15] : t[14];
  assign t[80] = (~t[101] & t[102]);
  assign t[81] = (~t[103] & t[104]);
  assign t[82] = (~t[103] & t[105]);
  assign t[83] = (~t[95] & t[106]);
  assign t[84] = (~t[107] & t[108]);
  assign t[85] = (~t[103] & t[109]);
  assign t[86] = (~t[95] & t[110]);
  assign t[87] = (~t[97] & t[111]);
  assign t[88] = (~t[97] & t[112]);
  assign t[89] = (~t[95] & t[113]);
  assign t[8] = ~(t[13] | t[16]);
  assign t[90] = (~t[97] & t[114]);
  assign t[91] = t[115] ^ x[4];
  assign t[92] = t[116] ^ x[5];
  assign t[93] = t[117] ^ x[8];
  assign t[94] = t[118] ^ x[9];
  assign t[95] = t[119] ^ x[14];
  assign t[96] = t[120] ^ x[15];
  assign t[97] = t[121] ^ x[20];
  assign t[98] = t[122] ^ x[21];
  assign t[99] = t[123] ^ x[24];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [58:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[11];
  assign t[101] = t[127] ^ x[16];
  assign t[102] = t[128] ^ x[17];
  assign t[103] = t[129] ^ x[21];
  assign t[104] = t[130] ^ x[22];
  assign t[105] = t[131] ^ x[24];
  assign t[106] = t[132] ^ x[25];
  assign t[107] = t[133] ^ x[27];
  assign t[108] = t[134] ^ x[28];
  assign t[109] = t[135] ^ x[30];
  assign t[10] = ~(t[14] & t[15]);
  assign t[110] = t[136] ^ x[31];
  assign t[111] = t[137] ^ x[32];
  assign t[112] = t[138] ^ x[33];
  assign t[113] = t[139] ^ x[38];
  assign t[114] = t[140] ^ x[39];
  assign t[115] = t[141] ^ x[41];
  assign t[116] = t[142] ^ x[42];
  assign t[117] = t[143] ^ x[47];
  assign t[118] = t[144] ^ x[48];
  assign t[119] = t[145] ^ x[50];
  assign t[11] = ~(t[16]);
  assign t[120] = t[146] ^ x[51];
  assign t[121] = t[147] ^ x[56];
  assign t[122] = t[148] ^ x[57];
  assign t[123] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[124] = (x[3]);
  assign t[125] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[126] = (x[6]);
  assign t[127] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[128] = (x[15]);
  assign t[129] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(x[19]);
  assign t[130] = (x[20]);
  assign t[131] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[23]);
  assign t[133] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[26]);
  assign t[135] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[29]);
  assign t[137] = (x[2]);
  assign t[138] = (x[7]);
  assign t[139] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[37]);
  assign t[141] = (x[1]);
  assign t[142] = (x[8]);
  assign t[143] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[144] = (x[46]);
  assign t[145] = (x[0]);
  assign t[146] = (x[9]);
  assign t[147] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[148] = (x[55]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[8]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(x[19]);
  assign t[18] = ~(t[52] | t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[52] & t[26]);
  assign t[22] = ~(t[53] & t[27]);
  assign t[23] = ~(t[24] & t[28]);
  assign t[24] = ~(t[54]);
  assign t[25] = ~(t[53]);
  assign t[26] = ~(t[55]);
  assign t[27] = ~(t[54] | t[29]);
  assign t[28] = t[30] & t[55];
  assign t[29] = ~(t[26]);
  assign t[2] = ~(t[6] & t[49]);
  assign t[30] = ~(t[52] | t[53]);
  assign t[31] = ~(t[32] & t[33]);
  assign t[32] = t[3] ? t[35] : t[34];
  assign t[33] = ~(t[6] & t[56]);
  assign t[34] = ~(t[57]);
  assign t[35] = ~(t[8] & t[36]);
  assign t[36] = t[13] ? x[40] : t[58];
  assign t[37] = ~(t[38] & t[39]);
  assign t[38] = t[3] ? t[41] : t[40];
  assign t[39] = ~(t[6] & t[59]);
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[8] & t[42]);
  assign t[42] = t[13] ? x[49] : t[61];
  assign t[43] = ~(t[44] & t[45]);
  assign t[44] = t[3] ? t[47] : t[46];
  assign t[45] = ~(t[6] & t[62]);
  assign t[46] = ~(t[63]);
  assign t[47] = ~(t[8] & t[48]);
  assign t[48] = t[13] ? x[58] : t[64];
  assign t[49] = (t[65]);
  assign t[4] = ~(t[50]);
  assign t[50] = (t[66]);
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = t[81] ^ x[5];
  assign t[66] = t[82] ^ x[11];
  assign t[67] = t[83] ^ x[17];
  assign t[68] = t[84] ^ x[22];
  assign t[69] = t[85] ^ x[25];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[28];
  assign t[71] = t[87] ^ x[31];
  assign t[72] = t[88] ^ x[32];
  assign t[73] = t[89] ^ x[33];
  assign t[74] = t[90] ^ x[39];
  assign t[75] = t[91] ^ x[41];
  assign t[76] = t[92] ^ x[42];
  assign t[77] = t[93] ^ x[48];
  assign t[78] = t[94] ^ x[50];
  assign t[79] = t[95] ^ x[51];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[57];
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[109] & t[110]);
  assign t[88] = (~t[97] & t[111]);
  assign t[89] = (~t[99] & t[112]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[90] = (~t[113] & t[114]);
  assign t[91] = (~t[97] & t[115]);
  assign t[92] = (~t[99] & t[116]);
  assign t[93] = (~t[117] & t[118]);
  assign t[94] = (~t[97] & t[119]);
  assign t[95] = (~t[99] & t[120]);
  assign t[96] = (~t[121] & t[122]);
  assign t[97] = t[123] ^ x[4];
  assign t[98] = t[124] ^ x[5];
  assign t[99] = t[125] ^ x[10];
  assign t[9] = t[13] ? x[18] : t[51];
  assign y = (t[0] & ~t[31] & ~t[37] & ~t[43]) | (~t[0] & t[31] & ~t[37] & ~t[43]) | (~t[0] & ~t[31] & t[37] & ~t[43]) | (~t[0] & ~t[31] & ~t[37] & t[43]) | (t[0] & t[31] & t[37] & ~t[43]) | (t[0] & t[31] & ~t[37] & t[43]) | (t[0] & ~t[31] & t[37] & t[43]) | (~t[0] & t[31] & t[37] & t[43]);
endmodule

module R2ind81(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = ~(x[19]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[8]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(x[19]);
  assign t[18] = ~(t[34] | t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[24] & t[28]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[35]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[26]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[35]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[17];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[71] = (x[15]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[13] ? x[18] : t[33];
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = ~(x[19]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[8]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(x[19]);
  assign t[18] = ~(t[34] | t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[24] & t[28]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[35]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[26]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[35]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[17];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[1]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[8]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[71] = (x[15]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[13] ? x[18] : t[33];
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = ~(x[19]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[8]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(x[19]);
  assign t[18] = ~(t[34] | t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[24] & t[28]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[35]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[26]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[35]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[17];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[2]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[71] = (x[15]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[13] ? x[18] : t[33];
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = ~(x[19]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[8]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(x[19]);
  assign t[18] = ~(t[34] | t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34] & t[26]);
  assign t[22] = ~(t[35] & t[27]);
  assign t[23] = ~(t[24] & t[28]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[35]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[36] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[26]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[35]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[17];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[16];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[71] = (x[15]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[13] ? x[18] : t[33];
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [58:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[11];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[21];
  assign t[106] = t[132] ^ x[22];
  assign t[107] = t[133] ^ x[24];
  assign t[108] = t[134] ^ x[25];
  assign t[109] = t[135] ^ x[27];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[136] ^ x[28];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[32];
  assign t[114] = t[140] ^ x[33];
  assign t[115] = t[141] ^ x[38];
  assign t[116] = t[142] ^ x[39];
  assign t[117] = t[143] ^ x[41];
  assign t[118] = t[144] ^ x[42];
  assign t[119] = t[145] ^ x[47];
  assign t[11] = ~(t[15]);
  assign t[120] = t[146] ^ x[48];
  assign t[121] = t[147] ^ x[50];
  assign t[122] = t[148] ^ x[51];
  assign t[123] = t[149] ^ x[56];
  assign t[124] = t[150] ^ x[57];
  assign t[125] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[126] = (x[0]);
  assign t[127] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[128] = (x[6]);
  assign t[129] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[15]);
  assign t[131] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[20]);
  assign t[133] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[23]);
  assign t[135] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[26]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[1]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (x[7]);
  assign t[141] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[142] = (x[37]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[146] = (x[46]);
  assign t[147] = (x[3]);
  assign t[148] = (x[9]);
  assign t[149] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[14] = ~(t[15]);
  assign t[150] = (x[55]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = t[12] ? x[40] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[49] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = t[12] ? x[58] : t[66];
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = t[83] ^ x[5];
  assign t[68] = t[84] ^ x[11];
  assign t[69] = t[85] ^ x[17];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[22];
  assign t[71] = t[87] ^ x[25];
  assign t[72] = t[88] ^ x[28];
  assign t[73] = t[89] ^ x[31];
  assign t[74] = t[90] ^ x[32];
  assign t[75] = t[91] ^ x[33];
  assign t[76] = t[92] ^ x[39];
  assign t[77] = t[93] ^ x[41];
  assign t[78] = t[94] ^ x[42];
  assign t[79] = t[95] ^ x[48];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[50];
  assign t[81] = t[97] ^ x[51];
  assign t[82] = t[98] ^ x[57];
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[99] & t[113]);
  assign t[91] = (~t[101] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = (~t[99] & t[117]);
  assign t[94] = (~t[101] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[99] & t[121]);
  assign t[97] = (~t[101] & t[122]);
  assign t[98] = (~t[123] & t[124]);
  assign t[99] = t[125] ^ x[4];
  assign t[9] = t[12] ? x[18] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind86(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [58:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[11];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[21];
  assign t[106] = t[132] ^ x[22];
  assign t[107] = t[133] ^ x[24];
  assign t[108] = t[134] ^ x[25];
  assign t[109] = t[135] ^ x[27];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[136] ^ x[28];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[32];
  assign t[114] = t[140] ^ x[33];
  assign t[115] = t[141] ^ x[38];
  assign t[116] = t[142] ^ x[39];
  assign t[117] = t[143] ^ x[41];
  assign t[118] = t[144] ^ x[42];
  assign t[119] = t[145] ^ x[47];
  assign t[11] = ~(t[15]);
  assign t[120] = t[146] ^ x[48];
  assign t[121] = t[147] ^ x[50];
  assign t[122] = t[148] ^ x[51];
  assign t[123] = t[149] ^ x[56];
  assign t[124] = t[150] ^ x[57];
  assign t[125] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[126] = (x[0]);
  assign t[127] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[128] = (x[6]);
  assign t[129] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[15]);
  assign t[131] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[20]);
  assign t[133] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[23]);
  assign t[135] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[26]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[1]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (x[7]);
  assign t[141] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[142] = (x[37]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[146] = (x[46]);
  assign t[147] = (x[3]);
  assign t[148] = (x[9]);
  assign t[149] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[14] = ~(t[15]);
  assign t[150] = (x[55]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = t[12] ? x[40] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[49] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = t[12] ? x[58] : t[66];
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = t[83] ^ x[5];
  assign t[68] = t[84] ^ x[11];
  assign t[69] = t[85] ^ x[17];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[22];
  assign t[71] = t[87] ^ x[25];
  assign t[72] = t[88] ^ x[28];
  assign t[73] = t[89] ^ x[31];
  assign t[74] = t[90] ^ x[32];
  assign t[75] = t[91] ^ x[33];
  assign t[76] = t[92] ^ x[39];
  assign t[77] = t[93] ^ x[41];
  assign t[78] = t[94] ^ x[42];
  assign t[79] = t[95] ^ x[48];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[50];
  assign t[81] = t[97] ^ x[51];
  assign t[82] = t[98] ^ x[57];
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[99] & t[113]);
  assign t[91] = (~t[101] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = (~t[99] & t[117]);
  assign t[94] = (~t[101] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[99] & t[121]);
  assign t[97] = (~t[101] & t[122]);
  assign t[98] = (~t[123] & t[124]);
  assign t[99] = t[125] ^ x[4];
  assign t[9] = t[12] ? x[18] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind91(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [52:0] x;
 output y;

 wire [142:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[124] ^ x[15];
  assign t[101] = t[125] ^ x[16];
  assign t[102] = t[126] ^ x[18];
  assign t[103] = t[127] ^ x[19];
  assign t[104] = t[128] ^ x[22];
  assign t[105] = t[129] ^ x[23];
  assign t[106] = t[130] ^ x[25];
  assign t[107] = t[131] ^ x[26];
  assign t[108] = t[132] ^ x[27];
  assign t[109] = t[133] ^ x[28];
  assign t[10] = t[16] ? x[13] : t[52];
  assign t[110] = t[134] ^ x[33];
  assign t[111] = t[135] ^ x[34];
  assign t[112] = t[136] ^ x[36];
  assign t[113] = t[137] ^ x[41];
  assign t[114] = t[138] ^ x[42];
  assign t[115] = t[139] ^ x[44];
  assign t[116] = t[140] ^ x[45];
  assign t[117] = t[141] ^ x[50];
  assign t[118] = t[142] ^ x[51];
  assign t[119] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[11] = ~(t[3]);
  assign t[120] = (x[0]);
  assign t[121] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[122] = (x[6]);
  assign t[123] = (x[2]);
  assign t[124] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[14]);
  assign t[126] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[17]);
  assign t[128] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[21]);
  assign t[12] = ~(t[53] | t[17]);
  assign t[130] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[24]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[135] = (x[31]);
  assign t[136] = (x[8]);
  assign t[137] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[138] = (x[39]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[18]);
  assign t[140] = (x[9]);
  assign t[141] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[142] = (x[47]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[54] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[20]);
  assign t[21] = ~(x[20]);
  assign t[22] = ~(t[55] | t[26]);
  assign t[23] = ~(t[55]);
  assign t[24] = t[27] & t[56];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[53] | t[54]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[53] & t[30]);
  assign t[2] = ~(t[6] & t[50]);
  assign t[30] = ~(t[56]);
  assign t[31] = ~(t[54]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[57]);
  assign t[35] = ~(t[58]);
  assign t[36] = ~(t[9] & t[37]);
  assign t[37] = t[16] ? x[35] : t[59];
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = ~(t[6] & t[52]);
  assign t[41] = ~(t[60]);
  assign t[42] = ~(t[9] & t[43]);
  assign t[43] = t[16] ? x[43] : t[61];
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[62]);
  assign t[47] = ~(t[63]);
  assign t[48] = ~(t[9] & t[49]);
  assign t[49] = t[16] ? x[52] : t[64];
  assign t[4] = ~(t[51]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = t[80] ^ x[5];
  assign t[66] = t[81] ^ x[11];
  assign t[67] = t[82] ^ x[12];
  assign t[68] = t[83] ^ x[16];
  assign t[69] = t[84] ^ x[19];
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = t[85] ^ x[23];
  assign t[71] = t[86] ^ x[26];
  assign t[72] = t[87] ^ x[27];
  assign t[73] = t[88] ^ x[28];
  assign t[74] = t[89] ^ x[34];
  assign t[75] = t[90] ^ x[36];
  assign t[76] = t[91] ^ x[42];
  assign t[77] = t[92] ^ x[44];
  assign t[78] = t[93] ^ x[45];
  assign t[79] = t[94] ^ x[51];
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[95] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[95] & t[108]);
  assign t[88] = (~t[97] & t[109]);
  assign t[89] = (~t[110] & t[111]);
  assign t[8] = ~(t[14]);
  assign t[90] = (~t[97] & t[112]);
  assign t[91] = (~t[113] & t[114]);
  assign t[92] = (~t[95] & t[115]);
  assign t[93] = (~t[97] & t[116]);
  assign t[94] = (~t[117] & t[118]);
  assign t[95] = t[119] ^ x[4];
  assign t[96] = t[120] ^ x[5];
  assign t[97] = t[121] ^ x[10];
  assign t[98] = t[122] ^ x[11];
  assign t[99] = t[123] ^ x[12];
  assign t[9] = ~(t[15]);
  assign y = (t[0] & ~t[32] & ~t[38] & ~t[44]) | (~t[0] & t[32] & ~t[38] & ~t[44]) | (~t[0] & ~t[32] & t[38] & ~t[44]) | (~t[0] & ~t[32] & ~t[38] & t[44]) | (t[0] & t[32] & t[38] & ~t[44]) | (t[0] & t[32] & ~t[38] & t[44]) | (t[0] & ~t[32] & t[38] & t[44]) | (~t[0] & t[32] & t[38] & t[44]);
endmodule

module R2ind96(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[9]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[13]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[8]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[14]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[7]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[14]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[13] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[20]);
  assign t[21] = ~(x[20]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[12];
  assign t[42] = t[49] ^ x[16];
  assign t[43] = t[50] ^ x[19];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[53] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[12];
  assign t[58] = t[71] ^ x[15];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[73] ^ x[18];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[2]);
  assign t[71] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[14]);
  assign t[73] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[17]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[22];
  assign t[101] = t[123] ^ x[24];
  assign t[102] = t[124] ^ x[25];
  assign t[103] = t[125] ^ x[27];
  assign t[104] = t[126] ^ x[28];
  assign t[105] = t[127] ^ x[30];
  assign t[106] = t[128] ^ x[31];
  assign t[107] = t[129] ^ x[32];
  assign t[108] = t[130] ^ x[33];
  assign t[109] = t[131] ^ x[38];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[132] ^ x[39];
  assign t[111] = t[133] ^ x[41];
  assign t[112] = t[134] ^ x[42];
  assign t[113] = t[135] ^ x[44];
  assign t[114] = t[136] ^ x[45];
  assign t[115] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[116] = (x[0]);
  assign t[117] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[118] = (x[6]);
  assign t[119] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[11] = ~(t[15]);
  assign t[120] = (x[14]);
  assign t[121] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[20]);
  assign t[123] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[23]);
  assign t[125] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[26]);
  assign t[127] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[29]);
  assign t[129] = (x[1]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[7]);
  assign t[131] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[132] = (x[36]);
  assign t[133] = (x[2]);
  assign t[134] = (x[8]);
  assign t[135] = (x[3]);
  assign t[136] = (x[9]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = t[12] ? x[40] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[43] : t[62];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[63]);
  assign t[48] = ~(t[64]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = t[12] ? x[46] : t[61];
  assign t[51] = (t[65]);
  assign t[52] = (t[66]);
  assign t[53] = (t[67]);
  assign t[54] = (t[68]);
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = t[79] ^ x[5];
  assign t[66] = t[80] ^ x[11];
  assign t[67] = t[81] ^ x[17];
  assign t[68] = t[82] ^ x[22];
  assign t[69] = t[83] ^ x[25];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[84] ^ x[28];
  assign t[71] = t[85] ^ x[31];
  assign t[72] = t[86] ^ x[32];
  assign t[73] = t[87] ^ x[33];
  assign t[74] = t[88] ^ x[39];
  assign t[75] = t[89] ^ x[41];
  assign t[76] = t[90] ^ x[42];
  assign t[77] = t[91] ^ x[44];
  assign t[78] = t[92] ^ x[45];
  assign t[79] = (~t[93] & t[94]);
  assign t[7] = ~(t[10]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[93] & t[107]);
  assign t[87] = (~t[95] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[93] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[95] & t[112]);
  assign t[91] = (~t[93] & t[113]);
  assign t[92] = (~t[95] & t[114]);
  assign t[93] = t[115] ^ x[4];
  assign t[94] = t[116] ^ x[5];
  assign t[95] = t[117] ^ x[10];
  assign t[96] = t[118] ^ x[11];
  assign t[97] = t[119] ^ x[16];
  assign t[98] = t[120] ^ x[17];
  assign t[99] = t[121] ^ x[21];
  assign t[9] = t[12] ? x[18] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind101(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[14]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[14]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[12];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[54] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[12];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[2]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[13] : t[35];
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [25:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[13]);
  assign t[17] = ~(t[35] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[13]);
  assign t[21] = ~(t[36] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[37] | t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = t[30] & t[38];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[35] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[35] | t[36]);
  assign t[31] = ~(t[36]);
  assign t[32] = ~(t[38]);
  assign t[33] = (t[39]);
  assign t[34] = (t[40]);
  assign t[35] = (t[41]);
  assign t[36] = (t[42]);
  assign t[37] = (t[43]);
  assign t[38] = (t[44]);
  assign t[39] = t[45] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[46] ^ x[11];
  assign t[41] = t[47] ^ x[16];
  assign t[42] = t[48] ^ x[19];
  assign t[43] = t[49] ^ x[22];
  assign t[44] = t[50] ^ x[25];
  assign t[45] = (~t[51] & t[52]);
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = t[63] ^ x[4];
  assign t[52] = t[64] ^ x[5];
  assign t[53] = t[65] ^ x[10];
  assign t[54] = t[66] ^ x[11];
  assign t[55] = t[67] ^ x[15];
  assign t[56] = t[68] ^ x[16];
  assign t[57] = t[69] ^ x[18];
  assign t[58] = t[70] ^ x[19];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[24];
  assign t[62] = t[74] ^ x[25];
  assign t[63] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[64] = (x[2]);
  assign t[65] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[66] = (x[8]);
  assign t[67] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[14]);
  assign t[69] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[17]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[12] : t[34];
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [58:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[11];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[21];
  assign t[106] = t[132] ^ x[22];
  assign t[107] = t[133] ^ x[24];
  assign t[108] = t[134] ^ x[25];
  assign t[109] = t[135] ^ x[27];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[136] ^ x[28];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[32];
  assign t[114] = t[140] ^ x[33];
  assign t[115] = t[141] ^ x[38];
  assign t[116] = t[142] ^ x[39];
  assign t[117] = t[143] ^ x[41];
  assign t[118] = t[144] ^ x[42];
  assign t[119] = t[145] ^ x[47];
  assign t[11] = ~(t[15]);
  assign t[120] = t[146] ^ x[48];
  assign t[121] = t[147] ^ x[50];
  assign t[122] = t[148] ^ x[51];
  assign t[123] = t[149] ^ x[56];
  assign t[124] = t[150] ^ x[57];
  assign t[125] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[126] = (x[0]);
  assign t[127] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[128] = (x[6]);
  assign t[129] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[14]);
  assign t[131] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[20]);
  assign t[133] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[23]);
  assign t[135] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[26]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[1]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (x[7]);
  assign t[141] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[142] = (x[36]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[146] = (x[45]);
  assign t[147] = (x[3]);
  assign t[148] = (x[9]);
  assign t[149] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[14] = ~(t[15]);
  assign t[150] = (x[54]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = t[12] ? x[40] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[49] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = t[12] ? x[58] : t[66];
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = t[83] ^ x[5];
  assign t[68] = t[84] ^ x[11];
  assign t[69] = t[85] ^ x[17];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[22];
  assign t[71] = t[87] ^ x[25];
  assign t[72] = t[88] ^ x[28];
  assign t[73] = t[89] ^ x[31];
  assign t[74] = t[90] ^ x[32];
  assign t[75] = t[91] ^ x[33];
  assign t[76] = t[92] ^ x[39];
  assign t[77] = t[93] ^ x[41];
  assign t[78] = t[94] ^ x[42];
  assign t[79] = t[95] ^ x[48];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[50];
  assign t[81] = t[97] ^ x[51];
  assign t[82] = t[98] ^ x[57];
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[99] & t[113]);
  assign t[91] = (~t[101] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = (~t[99] & t[117]);
  assign t[94] = (~t[101] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[99] & t[121]);
  assign t[97] = (~t[101] & t[122]);
  assign t[98] = (~t[123] & t[124]);
  assign t[99] = t[125] ^ x[4];
  assign t[9] = t[12] ? x[18] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind106(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [58:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[11];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[21];
  assign t[106] = t[132] ^ x[22];
  assign t[107] = t[133] ^ x[24];
  assign t[108] = t[134] ^ x[25];
  assign t[109] = t[135] ^ x[27];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[136] ^ x[28];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[32];
  assign t[114] = t[140] ^ x[33];
  assign t[115] = t[141] ^ x[38];
  assign t[116] = t[142] ^ x[39];
  assign t[117] = t[143] ^ x[41];
  assign t[118] = t[144] ^ x[42];
  assign t[119] = t[145] ^ x[47];
  assign t[11] = ~(t[15]);
  assign t[120] = t[146] ^ x[48];
  assign t[121] = t[147] ^ x[50];
  assign t[122] = t[148] ^ x[51];
  assign t[123] = t[149] ^ x[56];
  assign t[124] = t[150] ^ x[57];
  assign t[125] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[126] = (x[0]);
  assign t[127] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[128] = (x[6]);
  assign t[129] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[14]);
  assign t[131] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[20]);
  assign t[133] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[23]);
  assign t[135] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[26]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[1]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (x[7]);
  assign t[141] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[142] = (x[36]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[146] = (x[45]);
  assign t[147] = (x[3]);
  assign t[148] = (x[9]);
  assign t[149] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[14] = ~(t[15]);
  assign t[150] = (x[54]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = t[12] ? x[40] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[49] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = t[12] ? x[58] : t[66];
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = t[83] ^ x[5];
  assign t[68] = t[84] ^ x[11];
  assign t[69] = t[85] ^ x[17];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[22];
  assign t[71] = t[87] ^ x[25];
  assign t[72] = t[88] ^ x[28];
  assign t[73] = t[89] ^ x[31];
  assign t[74] = t[90] ^ x[32];
  assign t[75] = t[91] ^ x[33];
  assign t[76] = t[92] ^ x[39];
  assign t[77] = t[93] ^ x[41];
  assign t[78] = t[94] ^ x[42];
  assign t[79] = t[95] ^ x[48];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[50];
  assign t[81] = t[97] ^ x[51];
  assign t[82] = t[98] ^ x[57];
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[99] & t[113]);
  assign t[91] = (~t[101] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = (~t[99] & t[117]);
  assign t[94] = (~t[101] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[99] & t[121]);
  assign t[97] = (~t[101] & t[122]);
  assign t[98] = (~t[123] & t[124]);
  assign t[99] = t[125] ^ x[4];
  assign t[9] = t[12] ? x[18] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind111(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [58:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[11];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[21];
  assign t[106] = t[132] ^ x[22];
  assign t[107] = t[133] ^ x[24];
  assign t[108] = t[134] ^ x[25];
  assign t[109] = t[135] ^ x[27];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[136] ^ x[28];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[32];
  assign t[114] = t[140] ^ x[33];
  assign t[115] = t[141] ^ x[38];
  assign t[116] = t[142] ^ x[39];
  assign t[117] = t[143] ^ x[41];
  assign t[118] = t[144] ^ x[42];
  assign t[119] = t[145] ^ x[47];
  assign t[11] = ~(t[15]);
  assign t[120] = t[146] ^ x[48];
  assign t[121] = t[147] ^ x[50];
  assign t[122] = t[148] ^ x[51];
  assign t[123] = t[149] ^ x[56];
  assign t[124] = t[150] ^ x[57];
  assign t[125] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[126] = (x[0]);
  assign t[127] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[128] = (x[6]);
  assign t[129] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[13]);
  assign t[131] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[20]);
  assign t[133] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[23]);
  assign t[135] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[26]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[1]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[140] = (x[7]);
  assign t[141] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[142] = (x[35]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[146] = (x[44]);
  assign t[147] = (x[3]);
  assign t[148] = (x[9]);
  assign t[149] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[14] = ~(t[15]);
  assign t[150] = (x[54]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = t[12] ? x[40] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[49] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = t[12] ? x[58] : t[66];
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = t[83] ^ x[5];
  assign t[68] = t[84] ^ x[11];
  assign t[69] = t[85] ^ x[17];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[22];
  assign t[71] = t[87] ^ x[25];
  assign t[72] = t[88] ^ x[28];
  assign t[73] = t[89] ^ x[31];
  assign t[74] = t[90] ^ x[32];
  assign t[75] = t[91] ^ x[33];
  assign t[76] = t[92] ^ x[39];
  assign t[77] = t[93] ^ x[41];
  assign t[78] = t[94] ^ x[42];
  assign t[79] = t[95] ^ x[48];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[50];
  assign t[81] = t[97] ^ x[51];
  assign t[82] = t[98] ^ x[57];
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[99] & t[113]);
  assign t[91] = (~t[101] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = (~t[99] & t[117]);
  assign t[94] = (~t[101] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[99] & t[121]);
  assign t[97] = (~t[101] & t[122]);
  assign t[98] = (~t[123] & t[124]);
  assign t[99] = t[125] ^ x[4];
  assign t[9] = t[12] ? x[18] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind116(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[13]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[13]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[13]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [58:0] x;
 output y;

 wire [151:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[4];
  assign t[101] = t[127] ^ x[5];
  assign t[102] = t[128] ^ x[10];
  assign t[103] = t[129] ^ x[11];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[18];
  assign t[106] = t[132] ^ x[21];
  assign t[107] = t[133] ^ x[22];
  assign t[108] = t[134] ^ x[24];
  assign t[109] = t[135] ^ x[25];
  assign t[10] = x[12] ? x[19] : t[54];
  assign t[110] = t[136] ^ x[27];
  assign t[111] = t[137] ^ x[28];
  assign t[112] = t[138] ^ x[30];
  assign t[113] = t[139] ^ x[31];
  assign t[114] = t[140] ^ x[32];
  assign t[115] = t[141] ^ x[33];
  assign t[116] = t[142] ^ x[38];
  assign t[117] = t[143] ^ x[39];
  assign t[118] = t[144] ^ x[41];
  assign t[119] = t[145] ^ x[42];
  assign t[11] = ~(t[3]);
  assign t[120] = t[146] ^ x[47];
  assign t[121] = t[147] ^ x[48];
  assign t[122] = t[148] ^ x[50];
  assign t[123] = t[149] ^ x[51];
  assign t[124] = t[150] ^ x[56];
  assign t[125] = t[151] ^ x[57];
  assign t[126] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[127] = (x[0]);
  assign t[128] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[129] = (x[6]);
  assign t[12] = ~(t[55] | t[16]);
  assign t[130] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[131] = (x[14]);
  assign t[132] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[133] = (x[20]);
  assign t[134] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[135] = (x[23]);
  assign t[136] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[137] = (x[26]);
  assign t[138] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[139] = (x[29]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[1]);
  assign t[141] = (x[7]);
  assign t[142] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[143] = (x[35]);
  assign t[144] = (x[2]);
  assign t[145] = (x[8]);
  assign t[146] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[147] = (x[44]);
  assign t[148] = (x[3]);
  assign t[149] = (x[9]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[150] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[151] = (x[53]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[56] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[57] | t[24]);
  assign t[21] = ~(t[57]);
  assign t[22] = t[25] & t[58];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[55] | t[56]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[55] & t[28]);
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[56]);
  assign t[2] = ~(t[6] & t[52]);
  assign t[30] = ~(t[31] & t[32]);
  assign t[31] = t[3] ? t[34] : t[33];
  assign t[32] = ~(t[6] & t[59]);
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[9] & t[35]);
  assign t[35] = t[36] ? x[40] : t[61];
  assign t[36] = ~(t[37]);
  assign t[37] = ~(x[12]);
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = ~(t[6] & t[62]);
  assign t[41] = ~(t[63]);
  assign t[42] = ~(t[9] & t[43]);
  assign t[43] = t[44] ? x[49] : t[64];
  assign t[44] = ~(t[37]);
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[65]);
  assign t[48] = ~(t[66]);
  assign t[49] = ~(t[9] & t[50]);
  assign t[4] = ~(t[53]);
  assign t[50] = t[51] ? x[58] : t[67];
  assign t[51] = ~(t[37]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = (t[83]);
  assign t[68] = t[84] ^ x[5];
  assign t[69] = t[85] ^ x[11];
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = t[86] ^ x[18];
  assign t[71] = t[87] ^ x[22];
  assign t[72] = t[88] ^ x[25];
  assign t[73] = t[89] ^ x[28];
  assign t[74] = t[90] ^ x[31];
  assign t[75] = t[91] ^ x[32];
  assign t[76] = t[92] ^ x[33];
  assign t[77] = t[93] ^ x[39];
  assign t[78] = t[94] ^ x[41];
  assign t[79] = t[95] ^ x[42];
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = t[96] ^ x[48];
  assign t[81] = t[97] ^ x[50];
  assign t[82] = t[98] ^ x[51];
  assign t[83] = t[99] ^ x[57];
  assign t[84] = (~t[100] & t[101]);
  assign t[85] = (~t[102] & t[103]);
  assign t[86] = (~t[104] & t[105]);
  assign t[87] = (~t[106] & t[107]);
  assign t[88] = (~t[108] & t[109]);
  assign t[89] = (~t[110] & t[111]);
  assign t[8] = ~(t[14]);
  assign t[90] = (~t[112] & t[113]);
  assign t[91] = (~t[100] & t[114]);
  assign t[92] = (~t[102] & t[115]);
  assign t[93] = (~t[116] & t[117]);
  assign t[94] = (~t[100] & t[118]);
  assign t[95] = (~t[102] & t[119]);
  assign t[96] = (~t[120] & t[121]);
  assign t[97] = (~t[100] & t[122]);
  assign t[98] = (~t[102] & t[123]);
  assign t[99] = (~t[124] & t[125]);
  assign t[9] = ~(t[15]);
  assign y = (t[0] & ~t[30] & ~t[38] & ~t[45]) | (~t[0] & t[30] & ~t[38] & ~t[45]) | (~t[0] & ~t[30] & t[38] & ~t[45]) | (~t[0] & ~t[30] & ~t[38] & t[45]) | (t[0] & t[30] & t[38] & ~t[45]) | (t[0] & t[30] & ~t[38] & t[45]) | (t[0] & ~t[30] & t[38] & t[45]) | (~t[0] & t[30] & t[38] & t[45]);
endmodule

module R2ind121(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[9]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[13]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[8]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[13]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[7]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[13]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [31:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = x[12] ? x[19] : t[32];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[33] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[34] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35] | t[24]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[25] & t[36];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[33] | t[34]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[33] & t[28]);
  assign t[28] = ~(t[36]);
  assign t[29] = ~(t[34]);
  assign t[2] = ~(t[6] & t[30]);
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = t[44] ^ x[5];
  assign t[38] = t[45] ^ x[11];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[22];
  assign t[41] = t[48] ^ x[25];
  assign t[42] = t[49] ^ x[28];
  assign t[43] = t[50] ^ x[31];
  assign t[44] = (~t[51] & t[52]);
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[31]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = t[65] ^ x[4];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[25];
  assign t[61] = t[75] ^ x[27];
  assign t[62] = t[76] ^ x[28];
  assign t[63] = t[77] ^ x[30];
  assign t[64] = t[78] ^ x[31];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[0]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[6]);
  assign t[69] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[14]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[75] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[26]);
  assign t[77] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[29]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [42:0] x;
 output y;

 wire [138:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[18];
  assign t[101] = t[123] ^ x[21];
  assign t[102] = t[124] ^ x[22];
  assign t[103] = t[125] ^ x[24];
  assign t[104] = t[126] ^ x[25];
  assign t[105] = t[127] ^ x[27];
  assign t[106] = t[128] ^ x[28];
  assign t[107] = t[129] ^ x[30];
  assign t[108] = t[130] ^ x[31];
  assign t[109] = t[131] ^ x[32];
  assign t[10] = ~(t[3]);
  assign t[110] = t[132] ^ x[33];
  assign t[111] = t[133] ^ x[34];
  assign t[112] = t[134] ^ x[36];
  assign t[113] = t[135] ^ x[37];
  assign t[114] = t[136] ^ x[38];
  assign t[115] = t[137] ^ x[40];
  assign t[116] = t[138] ^ x[41];
  assign t[117] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[118] = (x[0]);
  assign t[119] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[120] = (x[6]);
  assign t[121] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[122] = (x[14]);
  assign t[123] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[20]);
  assign t[125] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[23]);
  assign t[127] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[26]);
  assign t[129] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15]);
  assign t[130] = (x[29]);
  assign t[131] = (x[1]);
  assign t[132] = (x[7]);
  assign t[133] = (x[15]);
  assign t[134] = (x[2]);
  assign t[135] = (x[8]);
  assign t[136] = (x[16]);
  assign t[137] = (x[3]);
  assign t[138] = (x[9]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[53] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[55] | t[28]);
  assign t[24] = ~(t[55]);
  assign t[25] = t[29] & t[56];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[53] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[53] | t[54]);
  assign t[2] = ~(t[6] & t[50]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[56]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[57]);
  assign t[35] = ~(t[58]);
  assign t[36] = ~(t[8] & t[37]);
  assign t[37] = x[12] ? x[35] : t[59];
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[6] & t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = ~(t[8] & t[43]);
  assign t[43] = x[12] ? x[39] : t[62];
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[63]);
  assign t[47] = ~(t[64]);
  assign t[48] = ~(t[8] & t[49]);
  assign t[49] = x[12] ? x[42] : t[51];
  assign t[4] = ~(t[51]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = t[80] ^ x[5];
  assign t[66] = t[81] ^ x[11];
  assign t[67] = t[82] ^ x[18];
  assign t[68] = t[83] ^ x[22];
  assign t[69] = t[84] ^ x[25];
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = t[85] ^ x[28];
  assign t[71] = t[86] ^ x[31];
  assign t[72] = t[87] ^ x[32];
  assign t[73] = t[88] ^ x[33];
  assign t[74] = t[89] ^ x[34];
  assign t[75] = t[90] ^ x[36];
  assign t[76] = t[91] ^ x[37];
  assign t[77] = t[92] ^ x[38];
  assign t[78] = t[93] ^ x[40];
  assign t[79] = t[94] ^ x[41];
  assign t[7] = ~(t[11]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[95] & t[109]);
  assign t[88] = (~t[97] & t[110]);
  assign t[89] = (~t[99] & t[111]);
  assign t[8] = ~(t[12]);
  assign t[90] = (~t[95] & t[112]);
  assign t[91] = (~t[97] & t[113]);
  assign t[92] = (~t[99] & t[114]);
  assign t[93] = (~t[95] & t[115]);
  assign t[94] = (~t[97] & t[116]);
  assign t[95] = t[117] ^ x[4];
  assign t[96] = t[118] ^ x[5];
  assign t[97] = t[119] ^ x[10];
  assign t[98] = t[120] ^ x[11];
  assign t[99] = t[121] ^ x[17];
  assign t[9] = x[12] ? x[19] : t[52];
  assign y = (t[0] & ~t[32] & ~t[38] & ~t[44]) | (~t[0] & t[32] & ~t[38] & ~t[44]) | (~t[0] & ~t[32] & t[38] & ~t[44]) | (~t[0] & ~t[32] & ~t[38] & t[44]) | (t[0] & t[32] & t[38] & ~t[44]) | (t[0] & t[32] & ~t[38] & t[44]) | (t[0] & ~t[32] & t[38] & t[44]) | (~t[0] & t[32] & t[38] & t[44]);
endmodule

module R2ind126(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[13];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[20];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[55] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[13];
  assign t[58] = t[71] ^ x[16];
  assign t[59] = t[72] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[19];
  assign t[61] = t[74] ^ x[20];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[15]);
  assign t[73] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[18]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[14] : t[34];
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[8]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[16]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[7]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[15]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[14]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [42:0] x;
 output y;

 wire [138:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[18];
  assign t[101] = t[123] ^ x[21];
  assign t[102] = t[124] ^ x[22];
  assign t[103] = t[125] ^ x[24];
  assign t[104] = t[126] ^ x[25];
  assign t[105] = t[127] ^ x[27];
  assign t[106] = t[128] ^ x[28];
  assign t[107] = t[129] ^ x[30];
  assign t[108] = t[130] ^ x[31];
  assign t[109] = t[131] ^ x[32];
  assign t[10] = ~(t[3]);
  assign t[110] = t[132] ^ x[33];
  assign t[111] = t[133] ^ x[34];
  assign t[112] = t[134] ^ x[36];
  assign t[113] = t[135] ^ x[37];
  assign t[114] = t[136] ^ x[38];
  assign t[115] = t[137] ^ x[40];
  assign t[116] = t[138] ^ x[41];
  assign t[117] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[118] = (x[0]);
  assign t[119] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[120] = (x[6]);
  assign t[121] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[122] = (x[14]);
  assign t[123] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[20]);
  assign t[125] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[23]);
  assign t[127] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[26]);
  assign t[129] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15]);
  assign t[130] = (x[29]);
  assign t[131] = (x[1]);
  assign t[132] = (x[7]);
  assign t[133] = (x[15]);
  assign t[134] = (x[2]);
  assign t[135] = (x[8]);
  assign t[136] = (x[16]);
  assign t[137] = (x[3]);
  assign t[138] = (x[9]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[53] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[55] | t[28]);
  assign t[24] = ~(t[55]);
  assign t[25] = t[29] & t[56];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[53] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[53] | t[54]);
  assign t[2] = ~(t[6] & t[50]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[56]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[57]);
  assign t[35] = ~(t[58]);
  assign t[36] = ~(t[8] & t[37]);
  assign t[37] = x[12] ? x[35] : t[59];
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[6] & t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = ~(t[8] & t[43]);
  assign t[43] = x[12] ? x[39] : t[62];
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[63]);
  assign t[47] = ~(t[64]);
  assign t[48] = ~(t[8] & t[49]);
  assign t[49] = x[12] ? x[42] : t[51];
  assign t[4] = ~(t[51]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = t[80] ^ x[5];
  assign t[66] = t[81] ^ x[11];
  assign t[67] = t[82] ^ x[18];
  assign t[68] = t[83] ^ x[22];
  assign t[69] = t[84] ^ x[25];
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = t[85] ^ x[28];
  assign t[71] = t[86] ^ x[31];
  assign t[72] = t[87] ^ x[32];
  assign t[73] = t[88] ^ x[33];
  assign t[74] = t[89] ^ x[34];
  assign t[75] = t[90] ^ x[36];
  assign t[76] = t[91] ^ x[37];
  assign t[77] = t[92] ^ x[38];
  assign t[78] = t[93] ^ x[40];
  assign t[79] = t[94] ^ x[41];
  assign t[7] = ~(t[11]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[95] & t[109]);
  assign t[88] = (~t[97] & t[110]);
  assign t[89] = (~t[99] & t[111]);
  assign t[8] = ~(t[12]);
  assign t[90] = (~t[95] & t[112]);
  assign t[91] = (~t[97] & t[113]);
  assign t[92] = (~t[99] & t[114]);
  assign t[93] = (~t[95] & t[115]);
  assign t[94] = (~t[97] & t[116]);
  assign t[95] = t[117] ^ x[4];
  assign t[96] = t[118] ^ x[5];
  assign t[97] = t[119] ^ x[10];
  assign t[98] = t[120] ^ x[11];
  assign t[99] = t[121] ^ x[17];
  assign t[9] = x[12] ? x[19] : t[52];
  assign y = (t[0] & ~t[32] & ~t[38] & ~t[44]) | (~t[0] & t[32] & ~t[38] & ~t[44]) | (~t[0] & ~t[32] & t[38] & ~t[44]) | (~t[0] & ~t[32] & ~t[38] & t[44]) | (t[0] & t[32] & t[38] & ~t[44]) | (t[0] & t[32] & ~t[38] & t[44]) | (t[0] & ~t[32] & t[38] & t[44]) | (~t[0] & t[32] & t[38] & t[44]);
endmodule

module R2ind131(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[13];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[20];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[55] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[13];
  assign t[58] = t[71] ^ x[16];
  assign t[59] = t[72] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[19];
  assign t[61] = t[74] ^ x[20];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[15]);
  assign t[73] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[18]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[14] : t[34];
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[8]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[16]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[7]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[15]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[14]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind136(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [45:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[124] ^ x[4];
  assign t[101] = t[125] ^ x[5];
  assign t[102] = t[126] ^ x[10];
  assign t[103] = t[127] ^ x[11];
  assign t[104] = t[128] ^ x[15];
  assign t[105] = t[129] ^ x[16];
  assign t[106] = t[130] ^ x[21];
  assign t[107] = t[131] ^ x[22];
  assign t[108] = t[132] ^ x[24];
  assign t[109] = t[133] ^ x[25];
  assign t[10] = ~(t[13]);
  assign t[110] = t[134] ^ x[27];
  assign t[111] = t[135] ^ x[28];
  assign t[112] = t[136] ^ x[30];
  assign t[113] = t[137] ^ x[31];
  assign t[114] = t[138] ^ x[33];
  assign t[115] = t[139] ^ x[34];
  assign t[116] = t[140] ^ x[35];
  assign t[117] = t[141] ^ x[36];
  assign t[118] = t[142] ^ x[37];
  assign t[119] = t[143] ^ x[39];
  assign t[11] = ~(t[14]);
  assign t[120] = t[144] ^ x[40];
  assign t[121] = t[145] ^ x[41];
  assign t[122] = t[146] ^ x[43];
  assign t[123] = t[147] ^ x[44];
  assign t[124] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[125] = (x[0]);
  assign t[126] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[127] = (x[6]);
  assign t[128] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[14]);
  assign t[12] = t[54] ^ t[55];
  assign t[130] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[131] = (x[18]);
  assign t[132] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[133] = (x[23]);
  assign t[134] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[135] = (x[26]);
  assign t[136] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[137] = (x[29]);
  assign t[138] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[139] = (x[32]);
  assign t[13] = ~(t[15]);
  assign t[140] = (x[1]);
  assign t[141] = (x[7]);
  assign t[142] = (x[19]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[20]);
  assign t[146] = (x[3]);
  assign t[147] = (x[9]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[14]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[56] | t[25]);
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[27] & t[28]);
  assign t[24] = ~(t[56] & t[29]);
  assign t[25] = ~(t[57] & t[30]);
  assign t[26] = ~(t[27] & t[31]);
  assign t[27] = ~(t[58]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[59]);
  assign t[2] = ~(t[6] & t[52]);
  assign t[30] = ~(t[58] | t[32]);
  assign t[31] = t[33] & t[59];
  assign t[32] = ~(t[29]);
  assign t[33] = ~(t[56] | t[57]);
  assign t[34] = ~(t[35] & t[36]);
  assign t[35] = t[3] ? t[38] : t[37];
  assign t[36] = ~(t[6] & t[60]);
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[8] & t[39]);
  assign t[39] = x[12] ? x[38] : t[62];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[41] & t[42]);
  assign t[41] = t[3] ? t[44] : t[43];
  assign t[42] = ~(t[6] & t[63]);
  assign t[43] = ~(t[64]);
  assign t[44] = ~(t[8] & t[45]);
  assign t[45] = x[12] ? x[42] : t[65];
  assign t[46] = ~(t[47] & t[48]);
  assign t[47] = t[3] ? t[50] : t[49];
  assign t[48] = ~(t[6] & t[66]);
  assign t[49] = ~(t[67]);
  assign t[4] = ~(t[53]);
  assign t[50] = ~(t[8] & t[51]);
  assign t[51] = x[12] ? x[45] : t[53];
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = (t[83]);
  assign t[68] = t[84] ^ x[5];
  assign t[69] = t[85] ^ x[11];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[16];
  assign t[71] = t[87] ^ x[22];
  assign t[72] = t[88] ^ x[25];
  assign t[73] = t[89] ^ x[28];
  assign t[74] = t[90] ^ x[31];
  assign t[75] = t[91] ^ x[34];
  assign t[76] = t[92] ^ x[35];
  assign t[77] = t[93] ^ x[36];
  assign t[78] = t[94] ^ x[37];
  assign t[79] = t[95] ^ x[39];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[40];
  assign t[81] = t[97] ^ x[41];
  assign t[82] = t[98] ^ x[43];
  assign t[83] = t[99] ^ x[44];
  assign t[84] = (~t[100] & t[101]);
  assign t[85] = (~t[102] & t[103]);
  assign t[86] = (~t[104] & t[105]);
  assign t[87] = (~t[106] & t[107]);
  assign t[88] = (~t[108] & t[109]);
  assign t[89] = (~t[110] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[112] & t[113]);
  assign t[91] = (~t[114] & t[115]);
  assign t[92] = (~t[100] & t[116]);
  assign t[93] = (~t[102] & t[117]);
  assign t[94] = (~t[106] & t[118]);
  assign t[95] = (~t[100] & t[119]);
  assign t[96] = (~t[102] & t[120]);
  assign t[97] = (~t[106] & t[121]);
  assign t[98] = (~t[100] & t[122]);
  assign t[99] = (~t[102] & t[123]);
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0] & ~t[34] & ~t[40] & ~t[46]) | (~t[0] & t[34] & ~t[40] & ~t[46]) | (~t[0] & ~t[34] & t[40] & ~t[46]) | (~t[0] & ~t[34] & ~t[40] & t[46]) | (t[0] & t[34] & t[40] & ~t[46]) | (t[0] & t[34] & ~t[40] & t[46]) | (t[0] & ~t[34] & t[40] & t[46]) | (~t[0] & t[34] & t[40] & t[46]);
endmodule

module R2ind141(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [34:0] x;
 output y;

 wire [89:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = t[36] ^ t[37];
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(x[12]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[14]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[38] | t[25]);
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[27] & t[28]);
  assign t[24] = ~(t[38] & t[29]);
  assign t[25] = ~(t[39] & t[30]);
  assign t[26] = ~(t[27] & t[31]);
  assign t[27] = ~(t[40]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[41]);
  assign t[2] = ~(t[6] & t[34]);
  assign t[30] = ~(t[40] | t[32]);
  assign t[31] = t[33] & t[41];
  assign t[32] = ~(t[29]);
  assign t[33] = ~(t[38] | t[39]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[48]);
  assign t[41] = (t[49]);
  assign t[42] = t[50] ^ x[5];
  assign t[43] = t[51] ^ x[11];
  assign t[44] = t[52] ^ x[16];
  assign t[45] = t[53] ^ x[22];
  assign t[46] = t[54] ^ x[25];
  assign t[47] = t[55] ^ x[28];
  assign t[48] = t[56] ^ x[31];
  assign t[49] = t[57] ^ x[34];
  assign t[4] = ~(t[35]);
  assign t[50] = (~t[58] & t[59]);
  assign t[51] = (~t[60] & t[61]);
  assign t[52] = (~t[62] & t[63]);
  assign t[53] = (~t[64] & t[65]);
  assign t[54] = (~t[66] & t[67]);
  assign t[55] = (~t[68] & t[69]);
  assign t[56] = (~t[70] & t[71]);
  assign t[57] = (~t[72] & t[73]);
  assign t[58] = t[74] ^ x[4];
  assign t[59] = t[75] ^ x[5];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[76] ^ x[10];
  assign t[61] = t[77] ^ x[11];
  assign t[62] = t[78] ^ x[15];
  assign t[63] = t[79] ^ x[16];
  assign t[64] = t[80] ^ x[21];
  assign t[65] = t[81] ^ x[22];
  assign t[66] = t[82] ^ x[24];
  assign t[67] = t[83] ^ x[25];
  assign t[68] = t[84] ^ x[27];
  assign t[69] = t[85] ^ x[28];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[30];
  assign t[71] = t[87] ^ x[31];
  assign t[72] = t[88] ^ x[33];
  assign t[73] = t[89] ^ x[34];
  assign t[74] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[75] = (x[0]);
  assign t[76] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[77] = (x[6]);
  assign t[78] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[14]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[81] = (x[18]);
  assign t[82] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[23]);
  assign t[84] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[26]);
  assign t[86] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[29]);
  assign t[88] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[32]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [54:0] x;
 output y;

 wire [169:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (~t[112] & t[127]);
  assign t[101] = (~t[128] & t[129]);
  assign t[102] = (~t[116] & t[130]);
  assign t[103] = (~t[110] & t[131]);
  assign t[104] = (~t[112] & t[132]);
  assign t[105] = (~t[133] & t[134]);
  assign t[106] = (~t[116] & t[135]);
  assign t[107] = (~t[110] & t[136]);
  assign t[108] = (~t[112] & t[137]);
  assign t[109] = (~t[138] & t[139]);
  assign t[10] = ~(t[14]);
  assign t[110] = t[140] ^ x[4];
  assign t[111] = t[141] ^ x[5];
  assign t[112] = t[142] ^ x[10];
  assign t[113] = t[143] ^ x[11];
  assign t[114] = t[144] ^ x[15];
  assign t[115] = t[145] ^ x[16];
  assign t[116] = t[146] ^ x[21];
  assign t[117] = t[147] ^ x[22];
  assign t[118] = t[148] ^ x[24];
  assign t[119] = t[149] ^ x[25];
  assign t[11] = ~(t[15]);
  assign t[120] = t[150] ^ x[27];
  assign t[121] = t[151] ^ x[28];
  assign t[122] = t[152] ^ x[30];
  assign t[123] = t[153] ^ x[31];
  assign t[124] = t[154] ^ x[33];
  assign t[125] = t[155] ^ x[34];
  assign t[126] = t[156] ^ x[35];
  assign t[127] = t[157] ^ x[36];
  assign t[128] = t[158] ^ x[39];
  assign t[129] = t[159] ^ x[40];
  assign t[12] = ~(x[12]);
  assign t[130] = t[160] ^ x[41];
  assign t[131] = t[161] ^ x[42];
  assign t[132] = t[162] ^ x[43];
  assign t[133] = t[163] ^ x[46];
  assign t[134] = t[164] ^ x[47];
  assign t[135] = t[165] ^ x[48];
  assign t[136] = t[166] ^ x[49];
  assign t[137] = t[167] ^ x[50];
  assign t[138] = t[168] ^ x[53];
  assign t[139] = t[169] ^ x[54];
  assign t[13] = t[55] ^ t[56];
  assign t[140] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[141] = (x[0]);
  assign t[142] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[143] = (x[6]);
  assign t[144] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[145] = (x[14]);
  assign t[146] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[147] = (x[18]);
  assign t[148] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[149] = (x[23]);
  assign t[14] = ~(t[16]);
  assign t[150] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[151] = (x[26]);
  assign t[152] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[153] = (x[29]);
  assign t[154] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[155] = (x[32]);
  assign t[156] = (x[1]);
  assign t[157] = (x[7]);
  assign t[158] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[159] = (x[38]);
  assign t[15] = ~(t[17] | t[18]);
  assign t[160] = (x[19]);
  assign t[161] = (x[2]);
  assign t[162] = (x[8]);
  assign t[163] = (x[45] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[45] & 1'b0 & ~1'b0 & ~1'b0) | (~x[45] & ~1'b0 & 1'b0 & ~1'b0) | (~x[45] & ~1'b0 & ~1'b0 & 1'b0) | (x[45] & 1'b0 & 1'b0 & ~1'b0) | (x[45] & 1'b0 & ~1'b0 & 1'b0) | (x[45] & ~1'b0 & 1'b0 & 1'b0) | (~x[45] & 1'b0 & 1'b0 & 1'b0);
  assign t[164] = (x[45]);
  assign t[165] = (x[20]);
  assign t[166] = (x[3]);
  assign t[167] = (x[9]);
  assign t[168] = (x[52] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[52] & 1'b0 & ~1'b0 & ~1'b0) | (~x[52] & ~1'b0 & 1'b0 & ~1'b0) | (~x[52] & ~1'b0 & ~1'b0 & 1'b0) | (x[52] & 1'b0 & 1'b0 & ~1'b0) | (x[52] & 1'b0 & ~1'b0 & 1'b0) | (x[52] & ~1'b0 & 1'b0 & 1'b0) | (~x[52] & 1'b0 & 1'b0 & 1'b0);
  assign t[169] = (x[52]);
  assign t[16] = ~(t[19] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[57] & t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[8]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[60]);
  assign t[24] = ~(t[57] | t[26]);
  assign t[25] = ~(t[27]);
  assign t[26] = ~(t[59] & t[28]);
  assign t[27] = ~(t[21] & t[29]);
  assign t[28] = ~(t[58] | t[30]);
  assign t[29] = t[31] & t[60];
  assign t[2] = ~(t[6] & t[53]);
  assign t[30] = ~(t[23]);
  assign t[31] = ~(t[57] | t[59]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[61]);
  assign t[35] = ~(t[62]);
  assign t[36] = ~(t[8] & t[37]);
  assign t[37] = x[12] ? x[37] : t[38];
  assign t[38] = t[63] ^ t[64];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[65]);
  assign t[42] = ~(t[66]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[44] : t[45];
  assign t[45] = t[67] ^ t[68];
  assign t[46] = ~(t[47] & t[48]);
  assign t[47] = t[3] ? t[50] : t[49];
  assign t[48] = ~(t[6] & t[69]);
  assign t[49] = ~(t[70]);
  assign t[4] = ~(t[54]);
  assign t[50] = ~(t[8] & t[51]);
  assign t[51] = x[12] ? x[51] : t[52];
  assign t[52] = t[71] ^ t[54];
  assign t[53] = (t[72]);
  assign t[54] = (t[73]);
  assign t[55] = (t[74]);
  assign t[56] = (t[75]);
  assign t[57] = (t[76]);
  assign t[58] = (t[77]);
  assign t[59] = (t[78]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[79]);
  assign t[61] = (t[80]);
  assign t[62] = (t[81]);
  assign t[63] = (t[82]);
  assign t[64] = (t[83]);
  assign t[65] = (t[84]);
  assign t[66] = (t[85]);
  assign t[67] = (t[86]);
  assign t[68] = (t[87]);
  assign t[69] = (t[88]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (t[89]);
  assign t[71] = (t[90]);
  assign t[72] = t[91] ^ x[5];
  assign t[73] = t[92] ^ x[11];
  assign t[74] = t[93] ^ x[16];
  assign t[75] = t[94] ^ x[22];
  assign t[76] = t[95] ^ x[25];
  assign t[77] = t[96] ^ x[28];
  assign t[78] = t[97] ^ x[31];
  assign t[79] = t[98] ^ x[34];
  assign t[7] = ~(t[10]);
  assign t[80] = t[99] ^ x[35];
  assign t[81] = t[100] ^ x[36];
  assign t[82] = t[101] ^ x[40];
  assign t[83] = t[102] ^ x[41];
  assign t[84] = t[103] ^ x[42];
  assign t[85] = t[104] ^ x[43];
  assign t[86] = t[105] ^ x[47];
  assign t[87] = t[106] ^ x[48];
  assign t[88] = t[107] ^ x[49];
  assign t[89] = t[108] ^ x[50];
  assign t[8] = ~(t[11] & t[12]);
  assign t[90] = t[109] ^ x[54];
  assign t[91] = (~t[110] & t[111]);
  assign t[92] = (~t[112] & t[113]);
  assign t[93] = (~t[114] & t[115]);
  assign t[94] = (~t[116] & t[117]);
  assign t[95] = (~t[118] & t[119]);
  assign t[96] = (~t[120] & t[121]);
  assign t[97] = (~t[122] & t[123]);
  assign t[98] = (~t[124] & t[125]);
  assign t[99] = (~t[110] & t[126]);
  assign t[9] = x[12] ? x[13] : t[13];
  assign y = (t[0] & ~t[32] & ~t[39] & ~t[46]) | (~t[0] & t[32] & ~t[39] & ~t[46]) | (~t[0] & ~t[32] & t[39] & ~t[46]) | (~t[0] & ~t[32] & ~t[39] & t[46]) | (t[0] & t[32] & t[39] & ~t[46]) | (t[0] & t[32] & ~t[39] & t[46]) | (t[0] & ~t[32] & t[39] & t[46]) | (~t[0] & t[32] & t[39] & t[46]);
endmodule

module R2ind146(x, y);
 input [29:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(x[12]);
  assign t[13] = t[34] ^ t[35];
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[17] | t[18]);
  assign t[16] = ~(t[19] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[36] & t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[8]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[39]);
  assign t[24] = ~(t[36] | t[26]);
  assign t[25] = ~(t[27]);
  assign t[26] = ~(t[38] & t[28]);
  assign t[27] = ~(t[21] & t[29]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[39];
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[23]);
  assign t[31] = ~(t[36] | t[38]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[16];
  assign t[43] = t[51] ^ x[17];
  assign t[44] = t[52] ^ x[20];
  assign t[45] = t[53] ^ x[23];
  assign t[46] = t[54] ^ x[26];
  assign t[47] = t[55] ^ x[29];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[58] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = (~t[67] & t[68]);
  assign t[55] = (~t[69] & t[70]);
  assign t[56] = t[71] ^ x[4];
  assign t[57] = t[72] ^ x[5];
  assign t[58] = t[73] ^ x[10];
  assign t[59] = t[74] ^ x[11];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[75] ^ x[15];
  assign t[61] = t[76] ^ x[16];
  assign t[62] = t[77] ^ x[17];
  assign t[63] = t[78] ^ x[19];
  assign t[64] = t[79] ^ x[20];
  assign t[65] = t[80] ^ x[22];
  assign t[66] = t[81] ^ x[23];
  assign t[67] = t[82] ^ x[25];
  assign t[68] = t[83] ^ x[26];
  assign t[69] = t[84] ^ x[28];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[29];
  assign t[71] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[72] = (x[3]);
  assign t[73] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[74] = (x[9]);
  assign t[75] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[14]);
  assign t[77] = (x[6]);
  assign t[78] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[18]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[21]);
  assign t[82] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[24]);
  assign t[84] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[27]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[13] : t[13];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [34:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(x[12]);
  assign t[13] = t[34] ^ t[35];
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[17] | t[18]);
  assign t[16] = ~(t[19] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[36] & t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[8]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[39]);
  assign t[24] = ~(t[36] | t[26]);
  assign t[25] = ~(t[27]);
  assign t[26] = ~(t[38] & t[28]);
  assign t[27] = ~(t[21] & t[29]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[39];
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[23]);
  assign t[31] = ~(t[36] | t[38]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[16];
  assign t[43] = t[51] ^ x[22];
  assign t[44] = t[52] ^ x[25];
  assign t[45] = t[53] ^ x[28];
  assign t[46] = t[54] ^ x[31];
  assign t[47] = t[55] ^ x[34];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = t[72] ^ x[4];
  assign t[57] = t[73] ^ x[5];
  assign t[58] = t[74] ^ x[10];
  assign t[59] = t[75] ^ x[11];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[76] ^ x[15];
  assign t[61] = t[77] ^ x[16];
  assign t[62] = t[78] ^ x[21];
  assign t[63] = t[79] ^ x[22];
  assign t[64] = t[80] ^ x[24];
  assign t[65] = t[81] ^ x[25];
  assign t[66] = t[82] ^ x[27];
  assign t[67] = t[83] ^ x[28];
  assign t[68] = t[84] ^ x[30];
  assign t[69] = t[85] ^ x[31];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[33];
  assign t[71] = t[87] ^ x[34];
  assign t[72] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[73] = (x[2]);
  assign t[74] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[75] = (x[8]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[20]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[23]);
  assign t[82] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[26]);
  assign t[84] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[29]);
  assign t[86] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[32]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[13] : t[13];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [34:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(x[12]);
  assign t[13] = t[34] ^ t[35];
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[17] | t[18]);
  assign t[16] = ~(t[19] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[36] & t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[8]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[39]);
  assign t[24] = ~(t[36] | t[26]);
  assign t[25] = ~(t[27]);
  assign t[26] = ~(t[38] & t[28]);
  assign t[27] = ~(t[21] & t[29]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[39];
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[23]);
  assign t[31] = ~(t[36] | t[38]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[16];
  assign t[43] = t[51] ^ x[22];
  assign t[44] = t[52] ^ x[25];
  assign t[45] = t[53] ^ x[28];
  assign t[46] = t[54] ^ x[31];
  assign t[47] = t[55] ^ x[34];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = t[72] ^ x[4];
  assign t[57] = t[73] ^ x[5];
  assign t[58] = t[74] ^ x[10];
  assign t[59] = t[75] ^ x[11];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[76] ^ x[15];
  assign t[61] = t[77] ^ x[16];
  assign t[62] = t[78] ^ x[21];
  assign t[63] = t[79] ^ x[22];
  assign t[64] = t[80] ^ x[24];
  assign t[65] = t[81] ^ x[25];
  assign t[66] = t[82] ^ x[27];
  assign t[67] = t[83] ^ x[28];
  assign t[68] = t[84] ^ x[30];
  assign t[69] = t[85] ^ x[31];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[33];
  assign t[71] = t[87] ^ x[34];
  assign t[72] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[73] = (x[1]);
  assign t[74] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[75] = (x[7]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[19]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[23]);
  assign t[82] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[26]);
  assign t[84] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[29]);
  assign t[86] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[32]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[13] : t[13];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [34:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(x[12]);
  assign t[13] = t[34] ^ t[35];
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[17] | t[18]);
  assign t[16] = ~(t[19] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[36] & t[23]);
  assign t[19] = ~(t[24] | t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[8]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[39]);
  assign t[24] = ~(t[36] | t[26]);
  assign t[25] = ~(t[27]);
  assign t[26] = ~(t[38] & t[28]);
  assign t[27] = ~(t[21] & t[29]);
  assign t[28] = ~(t[37] | t[30]);
  assign t[29] = t[31] & t[39];
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[23]);
  assign t[31] = ~(t[36] | t[38]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[16];
  assign t[43] = t[51] ^ x[22];
  assign t[44] = t[52] ^ x[25];
  assign t[45] = t[53] ^ x[28];
  assign t[46] = t[54] ^ x[31];
  assign t[47] = t[55] ^ x[34];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = (~t[68] & t[69]);
  assign t[55] = (~t[70] & t[71]);
  assign t[56] = t[72] ^ x[4];
  assign t[57] = t[73] ^ x[5];
  assign t[58] = t[74] ^ x[10];
  assign t[59] = t[75] ^ x[11];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[76] ^ x[15];
  assign t[61] = t[77] ^ x[16];
  assign t[62] = t[78] ^ x[21];
  assign t[63] = t[79] ^ x[22];
  assign t[64] = t[80] ^ x[24];
  assign t[65] = t[81] ^ x[25];
  assign t[66] = t[82] ^ x[27];
  assign t[67] = t[83] ^ x[28];
  assign t[68] = t[84] ^ x[30];
  assign t[69] = t[85] ^ x[31];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[33];
  assign t[71] = t[87] ^ x[34];
  assign t[72] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[73] = (x[0]);
  assign t[74] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[75] = (x[6]);
  assign t[76] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[14]);
  assign t[78] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[79] = (x[18]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[23]);
  assign t[82] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[26]);
  assign t[84] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[29]);
  assign t[86] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[32]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[13] : t[13];
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [42:0] x;
 output y;

 wire [137:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[21];
  assign t[101] = t[123] ^ x[22];
  assign t[102] = t[124] ^ x[24];
  assign t[103] = t[125] ^ x[25];
  assign t[104] = t[126] ^ x[27];
  assign t[105] = t[127] ^ x[28];
  assign t[106] = t[128] ^ x[30];
  assign t[107] = t[129] ^ x[31];
  assign t[108] = t[130] ^ x[32];
  assign t[109] = t[131] ^ x[33];
  assign t[10] = ~(t[13]);
  assign t[110] = t[132] ^ x[34];
  assign t[111] = t[133] ^ x[36];
  assign t[112] = t[134] ^ x[37];
  assign t[113] = t[135] ^ x[38];
  assign t[114] = t[136] ^ x[40];
  assign t[115] = t[137] ^ x[41];
  assign t[116] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[117] = (x[0]);
  assign t[118] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[119] = (x[6]);
  assign t[11] = ~(t[14]);
  assign t[120] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[121] = (x[14]);
  assign t[122] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[20]);
  assign t[124] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[23]);
  assign t[126] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[26]);
  assign t[128] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[29]);
  assign t[12] = ~(x[12]);
  assign t[130] = (x[1]);
  assign t[131] = (x[7]);
  assign t[132] = (x[15]);
  assign t[133] = (x[2]);
  assign t[134] = (x[8]);
  assign t[135] = (x[16]);
  assign t[136] = (x[3]);
  assign t[137] = (x[9]);
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[52] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[8]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[53]);
  assign t[21] = ~(t[54]);
  assign t[22] = ~(t[55]);
  assign t[23] = ~(t[52] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[54] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[53] | t[29]);
  assign t[28] = t[30] & t[55];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6] & t[49]);
  assign t[30] = ~(t[52] | t[54]);
  assign t[31] = ~(t[32] & t[33]);
  assign t[32] = t[3] ? t[35] : t[34];
  assign t[33] = ~(t[6] & t[56]);
  assign t[34] = ~(t[57]);
  assign t[35] = ~(t[8] & t[36]);
  assign t[36] = x[12] ? x[35] : t[58];
  assign t[37] = ~(t[38] & t[39]);
  assign t[38] = t[3] ? t[41] : t[40];
  assign t[39] = ~(t[6] & t[59]);
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[8] & t[42]);
  assign t[42] = x[12] ? x[39] : t[61];
  assign t[43] = ~(t[44] & t[45]);
  assign t[44] = t[3] ? t[47] : t[46];
  assign t[45] = ~(t[6] & t[62]);
  assign t[46] = ~(t[63]);
  assign t[47] = ~(t[8] & t[48]);
  assign t[48] = x[12] ? x[42] : t[50];
  assign t[49] = (t[64]);
  assign t[4] = ~(t[50]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = t[79] ^ x[5];
  assign t[65] = t[80] ^ x[11];
  assign t[66] = t[81] ^ x[18];
  assign t[67] = t[82] ^ x[22];
  assign t[68] = t[83] ^ x[25];
  assign t[69] = t[84] ^ x[28];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[31];
  assign t[71] = t[86] ^ x[32];
  assign t[72] = t[87] ^ x[33];
  assign t[73] = t[88] ^ x[34];
  assign t[74] = t[89] ^ x[36];
  assign t[75] = t[90] ^ x[37];
  assign t[76] = t[91] ^ x[38];
  assign t[77] = t[92] ^ x[40];
  assign t[78] = t[93] ^ x[41];
  assign t[79] = (~t[94] & t[95]);
  assign t[7] = ~(t[10]);
  assign t[80] = (~t[96] & t[97]);
  assign t[81] = (~t[98] & t[99]);
  assign t[82] = (~t[100] & t[101]);
  assign t[83] = (~t[102] & t[103]);
  assign t[84] = (~t[104] & t[105]);
  assign t[85] = (~t[106] & t[107]);
  assign t[86] = (~t[94] & t[108]);
  assign t[87] = (~t[96] & t[109]);
  assign t[88] = (~t[98] & t[110]);
  assign t[89] = (~t[94] & t[111]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[90] = (~t[96] & t[112]);
  assign t[91] = (~t[98] & t[113]);
  assign t[92] = (~t[94] & t[114]);
  assign t[93] = (~t[96] & t[115]);
  assign t[94] = t[116] ^ x[4];
  assign t[95] = t[117] ^ x[5];
  assign t[96] = t[118] ^ x[10];
  assign t[97] = t[119] ^ x[11];
  assign t[98] = t[120] ^ x[17];
  assign t[99] = t[121] ^ x[18];
  assign t[9] = x[12] ? x[19] : t[51];
  assign y = (t[0] & ~t[31] & ~t[37] & ~t[43]) | (~t[0] & t[31] & ~t[37] & ~t[43]) | (~t[0] & ~t[31] & t[37] & ~t[43]) | (~t[0] & ~t[31] & ~t[37] & t[43]) | (t[0] & t[31] & t[37] & ~t[43]) | (t[0] & t[31] & ~t[37] & t[43]) | (t[0] & ~t[31] & t[37] & t[43]) | (~t[0] & t[31] & t[37] & t[43]);
endmodule

module R2ind151(x, y);
 input [26:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(x[12]);
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[34] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[8]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[34] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[36] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[35] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[36]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[13];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[20];
  assign t[43] = t[50] ^ x[23];
  assign t[44] = t[51] ^ x[26];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[54] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[5];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[11];
  assign t[56] = t[69] ^ x[13];
  assign t[57] = t[70] ^ x[16];
  assign t[58] = t[71] ^ x[17];
  assign t[59] = t[72] ^ x[19];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[20];
  assign t[61] = t[74] ^ x[22];
  assign t[62] = t[75] ^ x[23];
  assign t[63] = t[76] ^ x[25];
  assign t[64] = t[77] ^ x[26];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[3]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[15]);
  assign t[72] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[18]);
  assign t[74] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[21]);
  assign t[76] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[14] : t[33];
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(x[12]);
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[34] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[8]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[34] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[36] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[35] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[36]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[2]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[8]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[16]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(x[12]);
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[34] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[8]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[34] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[36] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[35] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[36]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[1]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[15]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(x[12]);
  assign t[13] = ~(t[15]);
  assign t[14] = ~(t[16] | t[17]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[34] & t[22]);
  assign t[18] = ~(t[23] | t[24]);
  assign t[19] = ~(t[8]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[34] | t[25]);
  assign t[24] = ~(t[26]);
  assign t[25] = ~(t[36] & t[27]);
  assign t[26] = ~(t[20] & t[28]);
  assign t[27] = ~(t[35] | t[29]);
  assign t[28] = t[30] & t[37];
  assign t[29] = ~(t[22]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[34] | t[36]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[14]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind156(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind161(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind166(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind171(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [46:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[22];
  assign t[101] = t[123] ^ x[24];
  assign t[102] = t[124] ^ x[25];
  assign t[103] = t[125] ^ x[27];
  assign t[104] = t[126] ^ x[28];
  assign t[105] = t[127] ^ x[30];
  assign t[106] = t[128] ^ x[31];
  assign t[107] = t[129] ^ x[32];
  assign t[108] = t[130] ^ x[33];
  assign t[109] = t[131] ^ x[35];
  assign t[10] = x[12] ? x[19] : t[53];
  assign t[110] = t[132] ^ x[36];
  assign t[111] = t[133] ^ x[38];
  assign t[112] = t[134] ^ x[39];
  assign t[113] = t[135] ^ x[44];
  assign t[114] = t[136] ^ x[45];
  assign t[115] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[116] = (x[0]);
  assign t[117] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[118] = (x[6]);
  assign t[119] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[11] = ~(t[3]);
  assign t[120] = (x[14]);
  assign t[121] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[20]);
  assign t[123] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[23]);
  assign t[125] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[26]);
  assign t[127] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[29]);
  assign t[129] = (x[1]);
  assign t[12] = ~(t[54] | t[16]);
  assign t[130] = (x[7]);
  assign t[131] = (x[2]);
  assign t[132] = (x[8]);
  assign t[133] = (x[3]);
  assign t[134] = (x[9]);
  assign t[135] = (x[40] & ~x[41] & ~x[42] & ~x[43]) | (~x[40] & x[41] & ~x[42] & ~x[43]) | (~x[40] & ~x[41] & x[42] & ~x[43]) | (~x[40] & ~x[41] & ~x[42] & x[43]) | (x[40] & x[41] & x[42] & ~x[43]) | (x[40] & x[41] & ~x[42] & x[43]) | (x[40] & ~x[41] & x[42] & x[43]) | (~x[40] & x[41] & x[42] & x[43]);
  assign t[136] = (x[41]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[55] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[56] | t[24]);
  assign t[21] = ~(t[56]);
  assign t[22] = t[25] & t[57];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[54] | t[55]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[54] & t[28]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[55]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[31] & t[32]);
  assign t[31] = t[3] ? t[34] : t[33];
  assign t[32] = ~(t[6] & t[58]);
  assign t[33] = ~(t[59]);
  assign t[34] = ~(t[9] & t[35]);
  assign t[35] = t[36] ? x[34] : t[59];
  assign t[36] = ~(t[37]);
  assign t[37] = ~(x[12]);
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = ~(t[6] & t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = ~(t[9] & t[43]);
  assign t[43] = t[44] ? x[37] : t[58];
  assign t[44] = ~(t[37]);
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[62]);
  assign t[48] = ~(t[63]);
  assign t[49] = ~(t[9] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[46] : t[64];
  assign t[51] = (t[65]);
  assign t[52] = (t[66]);
  assign t[53] = (t[67]);
  assign t[54] = (t[68]);
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = t[79] ^ x[5];
  assign t[66] = t[80] ^ x[11];
  assign t[67] = t[81] ^ x[18];
  assign t[68] = t[82] ^ x[22];
  assign t[69] = t[83] ^ x[25];
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = t[84] ^ x[28];
  assign t[71] = t[85] ^ x[31];
  assign t[72] = t[86] ^ x[32];
  assign t[73] = t[87] ^ x[33];
  assign t[74] = t[88] ^ x[35];
  assign t[75] = t[89] ^ x[36];
  assign t[76] = t[90] ^ x[38];
  assign t[77] = t[91] ^ x[39];
  assign t[78] = t[92] ^ x[45];
  assign t[79] = (~t[93] & t[94]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[93] & t[107]);
  assign t[87] = (~t[95] & t[108]);
  assign t[88] = (~t[93] & t[109]);
  assign t[89] = (~t[95] & t[110]);
  assign t[8] = ~(t[14]);
  assign t[90] = (~t[93] & t[111]);
  assign t[91] = (~t[95] & t[112]);
  assign t[92] = (~t[113] & t[114]);
  assign t[93] = t[115] ^ x[4];
  assign t[94] = t[116] ^ x[5];
  assign t[95] = t[117] ^ x[10];
  assign t[96] = t[118] ^ x[11];
  assign t[97] = t[119] ^ x[17];
  assign t[98] = t[120] ^ x[18];
  assign t[99] = t[121] ^ x[21];
  assign t[9] = ~(t[15]);
  assign y = (t[0] & ~t[30] & ~t[38] & ~t[45]) | (~t[0] & t[30] & ~t[38] & ~t[45]) | (~t[0] & ~t[30] & t[38] & ~t[45]) | (~t[0] & ~t[30] & ~t[38] & t[45]) | (t[0] & t[30] & t[38] & ~t[45]) | (t[0] & t[30] & ~t[38] & t[45]) | (t[0] & ~t[30] & t[38] & t[45]) | (~t[0] & t[30] & t[38] & t[45]);
endmodule

module R2ind176(x, y);
 input [31:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = x[12] ? x[19] : t[32];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[33] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[34] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35] | t[24]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[25] & t[36];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[33] | t[34]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[33] & t[28]);
  assign t[28] = ~(t[36]);
  assign t[29] = ~(t[34]);
  assign t[2] = ~(t[6] & t[30]);
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = t[44] ^ x[5];
  assign t[38] = t[45] ^ x[11];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[22];
  assign t[41] = t[48] ^ x[25];
  assign t[42] = t[49] ^ x[28];
  assign t[43] = t[50] ^ x[31];
  assign t[44] = (~t[51] & t[52]);
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[31]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = t[65] ^ x[4];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[25];
  assign t[61] = t[75] ^ x[27];
  assign t[62] = t[76] ^ x[28];
  assign t[63] = t[77] ^ x[30];
  assign t[64] = t[78] ^ x[31];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[3]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[9]);
  assign t[69] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[14]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[75] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[26]);
  assign t[77] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[29]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[13] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[20]);
  assign t[21] = ~(x[20]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[12];
  assign t[42] = t[49] ^ x[16];
  assign t[43] = t[50] ^ x[19];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[53] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[12];
  assign t[58] = t[71] ^ x[15];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[73] ^ x[18];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[2]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[8]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[1]);
  assign t[71] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[14]);
  assign t[73] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[17]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [25:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[12] : t[33];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[34] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[35] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(x[19]);
  assign t[22] = ~(t[36] | t[26]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[27] & t[37];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[34] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[37]);
  assign t[31] = ~(t[35]);
  assign t[32] = (t[38]);
  assign t[33] = (t[39]);
  assign t[34] = (t[40]);
  assign t[35] = (t[41]);
  assign t[36] = (t[42]);
  assign t[37] = (t[43]);
  assign t[38] = t[44] ^ x[5];
  assign t[39] = t[45] ^ x[11];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[46] ^ x[15];
  assign t[41] = t[47] ^ x[18];
  assign t[42] = t[48] ^ x[22];
  assign t[43] = t[49] ^ x[25];
  assign t[44] = (~t[50] & t[51]);
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[33]);
  assign t[50] = t[62] ^ x[4];
  assign t[51] = t[63] ^ x[5];
  assign t[52] = t[64] ^ x[10];
  assign t[53] = t[65] ^ x[11];
  assign t[54] = t[66] ^ x[14];
  assign t[55] = t[67] ^ x[15];
  assign t[56] = t[68] ^ x[17];
  assign t[57] = t[69] ^ x[18];
  assign t[58] = t[70] ^ x[21];
  assign t[59] = t[71] ^ x[22];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[72] ^ x[24];
  assign t[61] = t[73] ^ x[25];
  assign t[62] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[63] = (x[1]);
  assign t[64] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[65] = (x[7]);
  assign t[66] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[13]);
  assign t[68] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[20]);
  assign t[72] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[23]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [31:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = x[12] ? x[19] : t[32];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[33] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[34] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35] | t[24]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[25] & t[36];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[33] | t[34]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[33] & t[28]);
  assign t[28] = ~(t[36]);
  assign t[29] = ~(t[34]);
  assign t[2] = ~(t[6] & t[30]);
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = t[44] ^ x[5];
  assign t[38] = t[45] ^ x[11];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[22];
  assign t[41] = t[48] ^ x[25];
  assign t[42] = t[49] ^ x[28];
  assign t[43] = t[50] ^ x[31];
  assign t[44] = (~t[51] & t[52]);
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[31]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = t[65] ^ x[4];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[25];
  assign t[61] = t[75] ^ x[27];
  assign t[62] = t[76] ^ x[28];
  assign t[63] = t[77] ^ x[30];
  assign t[64] = t[78] ^ x[31];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[0]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[6]);
  assign t[69] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[14]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[75] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[26]);
  assign t[77] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[29]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [58:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[10];
  assign t[102] = t[128] ^ x[11];
  assign t[103] = t[129] ^ x[16];
  assign t[104] = t[130] ^ x[17];
  assign t[105] = t[131] ^ x[20];
  assign t[106] = t[132] ^ x[21];
  assign t[107] = t[133] ^ x[23];
  assign t[108] = t[134] ^ x[24];
  assign t[109] = t[135] ^ x[27];
  assign t[10] = t[16] ? x[18] : t[53];
  assign t[110] = t[136] ^ x[28];
  assign t[111] = t[137] ^ x[30];
  assign t[112] = t[138] ^ x[31];
  assign t[113] = t[139] ^ x[32];
  assign t[114] = t[140] ^ x[33];
  assign t[115] = t[141] ^ x[38];
  assign t[116] = t[142] ^ x[39];
  assign t[117] = t[143] ^ x[41];
  assign t[118] = t[144] ^ x[42];
  assign t[119] = t[145] ^ x[47];
  assign t[11] = ~(t[3]);
  assign t[120] = t[146] ^ x[48];
  assign t[121] = t[147] ^ x[50];
  assign t[122] = t[148] ^ x[51];
  assign t[123] = t[149] ^ x[56];
  assign t[124] = t[150] ^ x[57];
  assign t[125] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[126] = (x[0]);
  assign t[127] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[128] = (x[6]);
  assign t[129] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[12] = ~(t[54] | t[17]);
  assign t[130] = (x[13]);
  assign t[131] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[19]);
  assign t[133] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[22]);
  assign t[135] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[26]);
  assign t[137] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[29]);
  assign t[139] = (x[1]);
  assign t[13] = ~(t[18]);
  assign t[140] = (x[7]);
  assign t[141] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[142] = (x[35]);
  assign t[143] = (x[2]);
  assign t[144] = (x[8]);
  assign t[145] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[146] = (x[44]);
  assign t[147] = (x[3]);
  assign t[148] = (x[9]);
  assign t[149] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[150] = (x[53]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[55] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[56] | t[26]);
  assign t[23] = ~(t[56]);
  assign t[24] = t[27] & t[57];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[54] | t[55]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[54] & t[30]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = ~(t[57]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[58]);
  assign t[35] = ~(t[59]);
  assign t[36] = ~(t[9] & t[37]);
  assign t[37] = t[38] ? x[40] : t[60];
  assign t[38] = ~(t[21]);
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[9] & t[44]);
  assign t[44] = x[25] ? x[49] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[9] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[25] ? x[58] : t[66];
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = t[83] ^ x[5];
  assign t[68] = t[84] ^ x[11];
  assign t[69] = t[85] ^ x[17];
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = t[86] ^ x[21];
  assign t[71] = t[87] ^ x[24];
  assign t[72] = t[88] ^ x[28];
  assign t[73] = t[89] ^ x[31];
  assign t[74] = t[90] ^ x[32];
  assign t[75] = t[91] ^ x[33];
  assign t[76] = t[92] ^ x[39];
  assign t[77] = t[93] ^ x[41];
  assign t[78] = t[94] ^ x[42];
  assign t[79] = t[95] ^ x[48];
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = t[96] ^ x[50];
  assign t[81] = t[97] ^ x[51];
  assign t[82] = t[98] ^ x[57];
  assign t[83] = (~t[99] & t[100]);
  assign t[84] = (~t[101] & t[102]);
  assign t[85] = (~t[103] & t[104]);
  assign t[86] = (~t[105] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[109] & t[110]);
  assign t[89] = (~t[111] & t[112]);
  assign t[8] = ~(t[14]);
  assign t[90] = (~t[99] & t[113]);
  assign t[91] = (~t[101] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = (~t[99] & t[117]);
  assign t[94] = (~t[101] & t[118]);
  assign t[95] = (~t[119] & t[120]);
  assign t[96] = (~t[99] & t[121]);
  assign t[97] = (~t[101] & t[122]);
  assign t[98] = (~t[123] & t[124]);
  assign t[99] = t[125] ^ x[4];
  assign t[9] = ~(t[15]);
  assign y = (t[0] & ~t[32] & ~t[39] & ~t[45]) | (~t[0] & t[32] & ~t[39] & ~t[45]) | (~t[0] & ~t[32] & t[39] & ~t[45]) | (~t[0] & ~t[32] & ~t[39] & t[45]) | (t[0] & t[32] & t[39] & ~t[45]) | (t[0] & t[32] & ~t[39] & t[45]) | (t[0] & ~t[32] & t[39] & t[45]) | (~t[0] & t[32] & t[39] & t[45]);
endmodule

module R2ind181(x, y);
 input [31:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = x[12] ? x[19] : t[32];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[33] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[34] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35] | t[24]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[25] & t[36];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[33] | t[34]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[33] & t[28]);
  assign t[28] = ~(t[36]);
  assign t[29] = ~(t[34]);
  assign t[2] = ~(t[6] & t[30]);
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = t[44] ^ x[5];
  assign t[38] = t[45] ^ x[11];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[22];
  assign t[41] = t[48] ^ x[25];
  assign t[42] = t[49] ^ x[28];
  assign t[43] = t[50] ^ x[31];
  assign t[44] = (~t[51] & t[52]);
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[31]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = t[65] ^ x[4];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[25];
  assign t[61] = t[75] ^ x[27];
  assign t[62] = t[76] ^ x[28];
  assign t[63] = t[77] ^ x[30];
  assign t[64] = t[78] ^ x[31];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[3]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[9]);
  assign t[69] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[14]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[75] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[26]);
  assign t[77] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[29]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [31:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = x[12] ? x[19] : t[32];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[33] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[34] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[35] | t[24]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[25] & t[36];
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[33] | t[34]);
  assign t[26] = ~(t[21] & t[29]);
  assign t[27] = ~(t[33] & t[28]);
  assign t[28] = ~(t[36]);
  assign t[29] = ~(t[34]);
  assign t[2] = ~(t[6] & t[30]);
  assign t[30] = (t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = t[44] ^ x[5];
  assign t[38] = t[45] ^ x[11];
  assign t[39] = t[46] ^ x[18];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[22];
  assign t[41] = t[48] ^ x[25];
  assign t[42] = t[49] ^ x[28];
  assign t[43] = t[50] ^ x[31];
  assign t[44] = (~t[51] & t[52]);
  assign t[45] = (~t[53] & t[54]);
  assign t[46] = (~t[55] & t[56]);
  assign t[47] = (~t[57] & t[58]);
  assign t[48] = (~t[59] & t[60]);
  assign t[49] = (~t[61] & t[62]);
  assign t[4] = ~(t[31]);
  assign t[50] = (~t[63] & t[64]);
  assign t[51] = t[65] ^ x[4];
  assign t[52] = t[66] ^ x[5];
  assign t[53] = t[67] ^ x[10];
  assign t[54] = t[68] ^ x[11];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[18];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[25];
  assign t[61] = t[75] ^ x[27];
  assign t[62] = t[76] ^ x[28];
  assign t[63] = t[77] ^ x[30];
  assign t[64] = t[78] ^ x[31];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[2]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[8]);
  assign t[69] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[14]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[75] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[26]);
  assign t[77] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[29]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[7]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[13]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[16] ? x[18] : t[34];
  assign t[11] = ~(t[3]);
  assign t[12] = ~(t[35] | t[17]);
  assign t[13] = ~(t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[14]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[36] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[25]);
  assign t[21] = ~(x[25]);
  assign t[22] = ~(t[37] | t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[27] & t[38];
  assign t[25] = ~(t[28] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[23] & t[31]);
  assign t[29] = ~(t[35] & t[30]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[38]);
  assign t[31] = ~(t[36]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[21];
  assign t[43] = t[50] ^ x[24];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[16];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[20];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[23];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[9] | t[11]);
  assign t[70] = (x[6]);
  assign t[71] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[72] = (x[13]);
  assign t[73] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[19]);
  assign t[75] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[22]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[12] | t[13]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [58:0] x;
 output y;

 wire [152:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (~t[125] & t[126]);
  assign t[101] = t[127] ^ x[4];
  assign t[102] = t[128] ^ x[5];
  assign t[103] = t[129] ^ x[10];
  assign t[104] = t[130] ^ x[11];
  assign t[105] = t[131] ^ x[17];
  assign t[106] = t[132] ^ x[18];
  assign t[107] = t[133] ^ x[21];
  assign t[108] = t[134] ^ x[22];
  assign t[109] = t[135] ^ x[24];
  assign t[10] = ~(t[12] & t[13]);
  assign t[110] = t[136] ^ x[25];
  assign t[111] = t[137] ^ x[27];
  assign t[112] = t[138] ^ x[28];
  assign t[113] = t[139] ^ x[30];
  assign t[114] = t[140] ^ x[31];
  assign t[115] = t[141] ^ x[32];
  assign t[116] = t[142] ^ x[33];
  assign t[117] = t[143] ^ x[38];
  assign t[118] = t[144] ^ x[39];
  assign t[119] = t[145] ^ x[41];
  assign t[11] = ~(t[14]);
  assign t[120] = t[146] ^ x[42];
  assign t[121] = t[147] ^ x[47];
  assign t[122] = t[148] ^ x[48];
  assign t[123] = t[149] ^ x[50];
  assign t[124] = t[150] ^ x[51];
  assign t[125] = t[151] ^ x[56];
  assign t[126] = t[152] ^ x[57];
  assign t[127] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[128] = (x[0]);
  assign t[129] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (x[6]);
  assign t[131] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[132] = (x[13]);
  assign t[133] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[20]);
  assign t[135] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[23]);
  assign t[137] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[26]);
  assign t[139] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[13] = ~(t[14]);
  assign t[140] = (x[29]);
  assign t[141] = (x[1]);
  assign t[142] = (x[7]);
  assign t[143] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[144] = (x[34]);
  assign t[145] = (x[2]);
  assign t[146] = (x[8]);
  assign t[147] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[148] = (x[43]);
  assign t[149] = (x[3]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[150] = (x[9]);
  assign t[151] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[152] = (x[55]);
  assign t[15] = ~(t[56] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[57] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[58] | t[27]);
  assign t[23] = ~(t[58]);
  assign t[24] = t[28] & t[59];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[56] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[56] | t[57]);
  assign t[29] = ~(t[57]);
  assign t[2] = ~(t[6] & t[53]);
  assign t[30] = ~(t[59]);
  assign t[31] = ~(t[32] & t[33]);
  assign t[32] = t[3] ? t[35] : t[34];
  assign t[33] = ~(t[6] & t[60]);
  assign t[34] = ~(t[61]);
  assign t[35] = ~(t[8] & t[36]);
  assign t[36] = t[37] ? x[40] : t[62];
  assign t[37] = ~(t[38]);
  assign t[38] = ~(x[12]);
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[63]);
  assign t[42] = ~(t[64]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[45] ? x[49] : t[65];
  assign t[45] = ~(t[38]);
  assign t[46] = ~(t[47] & t[48]);
  assign t[47] = t[3] ? t[50] : t[49];
  assign t[48] = ~(t[6] & t[66]);
  assign t[49] = ~(t[67]);
  assign t[4] = ~(t[54]);
  assign t[50] = ~(t[8] & t[51]);
  assign t[51] = t[52] ? x[58] : t[68];
  assign t[52] = ~(t[38]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = (t[83]);
  assign t[68] = (t[84]);
  assign t[69] = t[85] ^ x[5];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[11];
  assign t[71] = t[87] ^ x[18];
  assign t[72] = t[88] ^ x[22];
  assign t[73] = t[89] ^ x[25];
  assign t[74] = t[90] ^ x[28];
  assign t[75] = t[91] ^ x[31];
  assign t[76] = t[92] ^ x[32];
  assign t[77] = t[93] ^ x[33];
  assign t[78] = t[94] ^ x[39];
  assign t[79] = t[95] ^ x[41];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[42];
  assign t[81] = t[97] ^ x[48];
  assign t[82] = t[98] ^ x[50];
  assign t[83] = t[99] ^ x[51];
  assign t[84] = t[100] ^ x[57];
  assign t[85] = (~t[101] & t[102]);
  assign t[86] = (~t[103] & t[104]);
  assign t[87] = (~t[105] & t[106]);
  assign t[88] = (~t[107] & t[108]);
  assign t[89] = (~t[109] & t[110]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[111] & t[112]);
  assign t[91] = (~t[113] & t[114]);
  assign t[92] = (~t[101] & t[115]);
  assign t[93] = (~t[103] & t[116]);
  assign t[94] = (~t[117] & t[118]);
  assign t[95] = (~t[101] & t[119]);
  assign t[96] = (~t[103] & t[120]);
  assign t[97] = (~t[121] & t[122]);
  assign t[98] = (~t[101] & t[123]);
  assign t[99] = (~t[103] & t[124]);
  assign t[9] = x[12] ? x[19] : t[55];
  assign y = (t[0] & ~t[31] & ~t[39] & ~t[46]) | (~t[0] & t[31] & ~t[39] & ~t[46]) | (~t[0] & ~t[31] & t[39] & ~t[46]) | (~t[0] & ~t[31] & ~t[39] & t[46]) | (t[0] & t[31] & t[39] & ~t[46]) | (t[0] & t[31] & ~t[39] & t[46]) | (t[0] & ~t[31] & t[39] & t[46]) | (~t[0] & t[31] & t[39] & t[46]);
endmodule

module R2ind186(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[12]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[12]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [58:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[11];
  assign t[101] = t[127] ^ x[17];
  assign t[102] = t[128] ^ x[18];
  assign t[103] = t[129] ^ x[21];
  assign t[104] = t[130] ^ x[22];
  assign t[105] = t[131] ^ x[24];
  assign t[106] = t[132] ^ x[25];
  assign t[107] = t[133] ^ x[27];
  assign t[108] = t[134] ^ x[28];
  assign t[109] = t[135] ^ x[30];
  assign t[10] = ~(t[12] & t[13]);
  assign t[110] = t[136] ^ x[31];
  assign t[111] = t[137] ^ x[32];
  assign t[112] = t[138] ^ x[33];
  assign t[113] = t[139] ^ x[38];
  assign t[114] = t[140] ^ x[39];
  assign t[115] = t[141] ^ x[41];
  assign t[116] = t[142] ^ x[42];
  assign t[117] = t[143] ^ x[47];
  assign t[118] = t[144] ^ x[48];
  assign t[119] = t[145] ^ x[50];
  assign t[11] = ~(t[14]);
  assign t[120] = t[146] ^ x[51];
  assign t[121] = t[147] ^ x[56];
  assign t[122] = t[148] ^ x[57];
  assign t[123] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[124] = (x[0]);
  assign t[125] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[126] = (x[6]);
  assign t[127] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[128] = (x[13]);
  assign t[129] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (x[20]);
  assign t[131] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[23]);
  assign t[133] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[26]);
  assign t[135] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[29]);
  assign t[137] = (x[1]);
  assign t[138] = (x[7]);
  assign t[139] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[13] = ~(t[14]);
  assign t[140] = (x[34]);
  assign t[141] = (x[2]);
  assign t[142] = (x[8]);
  assign t[143] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[144] = (x[43]);
  assign t[145] = (x[3]);
  assign t[146] = (x[9]);
  assign t[147] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[148] = (x[52]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[52] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[53] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[54] | t[27]);
  assign t[23] = ~(t[54]);
  assign t[24] = t[28] & t[55];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[52] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[52] | t[53]);
  assign t[29] = ~(t[53]);
  assign t[2] = ~(t[6] & t[49]);
  assign t[30] = ~(t[55]);
  assign t[31] = ~(t[32] & t[33]);
  assign t[32] = t[3] ? t[35] : t[34];
  assign t[33] = ~(t[6] & t[56]);
  assign t[34] = ~(t[57]);
  assign t[35] = ~(t[8] & t[36]);
  assign t[36] = x[12] ? x[40] : t[58];
  assign t[37] = ~(t[38] & t[39]);
  assign t[38] = t[3] ? t[41] : t[40];
  assign t[39] = ~(t[6] & t[59]);
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[8] & t[42]);
  assign t[42] = x[12] ? x[49] : t[61];
  assign t[43] = ~(t[44] & t[45]);
  assign t[44] = t[3] ? t[47] : t[46];
  assign t[45] = ~(t[6] & t[62]);
  assign t[46] = ~(t[63]);
  assign t[47] = ~(t[8] & t[48]);
  assign t[48] = x[12] ? x[58] : t[64];
  assign t[49] = (t[65]);
  assign t[4] = ~(t[50]);
  assign t[50] = (t[66]);
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = t[81] ^ x[5];
  assign t[66] = t[82] ^ x[11];
  assign t[67] = t[83] ^ x[18];
  assign t[68] = t[84] ^ x[22];
  assign t[69] = t[85] ^ x[25];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[28];
  assign t[71] = t[87] ^ x[31];
  assign t[72] = t[88] ^ x[32];
  assign t[73] = t[89] ^ x[33];
  assign t[74] = t[90] ^ x[39];
  assign t[75] = t[91] ^ x[41];
  assign t[76] = t[92] ^ x[42];
  assign t[77] = t[93] ^ x[48];
  assign t[78] = t[94] ^ x[50];
  assign t[79] = t[95] ^ x[51];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[57];
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[109] & t[110]);
  assign t[88] = (~t[97] & t[111]);
  assign t[89] = (~t[99] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[113] & t[114]);
  assign t[91] = (~t[97] & t[115]);
  assign t[92] = (~t[99] & t[116]);
  assign t[93] = (~t[117] & t[118]);
  assign t[94] = (~t[97] & t[119]);
  assign t[95] = (~t[99] & t[120]);
  assign t[96] = (~t[121] & t[122]);
  assign t[97] = t[123] ^ x[4];
  assign t[98] = t[124] ^ x[5];
  assign t[99] = t[125] ^ x[10];
  assign t[9] = x[12] ? x[19] : t[51];
  assign y = (t[0] & ~t[31] & ~t[37] & ~t[43]) | (~t[0] & t[31] & ~t[37] & ~t[43]) | (~t[0] & ~t[31] & t[37] & ~t[43]) | (~t[0] & ~t[31] & ~t[37] & t[43]) | (t[0] & t[31] & t[37] & ~t[43]) | (t[0] & t[31] & ~t[37] & t[43]) | (t[0] & ~t[31] & t[37] & t[43]) | (~t[0] & t[31] & t[37] & t[43]);
endmodule

module R2ind191(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[2]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[8]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[1]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [58:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[126] ^ x[11];
  assign t[101] = t[127] ^ x[17];
  assign t[102] = t[128] ^ x[18];
  assign t[103] = t[129] ^ x[21];
  assign t[104] = t[130] ^ x[22];
  assign t[105] = t[131] ^ x[24];
  assign t[106] = t[132] ^ x[25];
  assign t[107] = t[133] ^ x[27];
  assign t[108] = t[134] ^ x[28];
  assign t[109] = t[135] ^ x[30];
  assign t[10] = ~(t[12] & t[13]);
  assign t[110] = t[136] ^ x[31];
  assign t[111] = t[137] ^ x[32];
  assign t[112] = t[138] ^ x[33];
  assign t[113] = t[139] ^ x[38];
  assign t[114] = t[140] ^ x[39];
  assign t[115] = t[141] ^ x[41];
  assign t[116] = t[142] ^ x[42];
  assign t[117] = t[143] ^ x[47];
  assign t[118] = t[144] ^ x[48];
  assign t[119] = t[145] ^ x[50];
  assign t[11] = ~(t[14]);
  assign t[120] = t[146] ^ x[51];
  assign t[121] = t[147] ^ x[56];
  assign t[122] = t[148] ^ x[57];
  assign t[123] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[124] = (x[0]);
  assign t[125] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[126] = (x[6]);
  assign t[127] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[128] = (x[13]);
  assign t[129] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (x[20]);
  assign t[131] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[23]);
  assign t[133] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[26]);
  assign t[135] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[29]);
  assign t[137] = (x[1]);
  assign t[138] = (x[7]);
  assign t[139] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[13] = ~(t[14]);
  assign t[140] = (x[34]);
  assign t[141] = (x[2]);
  assign t[142] = (x[8]);
  assign t[143] = (x[43] & ~x[44] & ~x[45] & ~x[46]) | (~x[43] & x[44] & ~x[45] & ~x[46]) | (~x[43] & ~x[44] & x[45] & ~x[46]) | (~x[43] & ~x[44] & ~x[45] & x[46]) | (x[43] & x[44] & x[45] & ~x[46]) | (x[43] & x[44] & ~x[45] & x[46]) | (x[43] & ~x[44] & x[45] & x[46]) | (~x[43] & x[44] & x[45] & x[46]);
  assign t[144] = (x[43]);
  assign t[145] = (x[3]);
  assign t[146] = (x[9]);
  assign t[147] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[148] = (x[52]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[52] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[53] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[54] | t[27]);
  assign t[23] = ~(t[54]);
  assign t[24] = t[28] & t[55];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[52] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[52] | t[53]);
  assign t[29] = ~(t[53]);
  assign t[2] = ~(t[6] & t[49]);
  assign t[30] = ~(t[55]);
  assign t[31] = ~(t[32] & t[33]);
  assign t[32] = t[3] ? t[35] : t[34];
  assign t[33] = ~(t[6] & t[56]);
  assign t[34] = ~(t[57]);
  assign t[35] = ~(t[8] & t[36]);
  assign t[36] = x[12] ? x[40] : t[58];
  assign t[37] = ~(t[38] & t[39]);
  assign t[38] = t[3] ? t[41] : t[40];
  assign t[39] = ~(t[6] & t[59]);
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[8] & t[42]);
  assign t[42] = x[12] ? x[49] : t[61];
  assign t[43] = ~(t[44] & t[45]);
  assign t[44] = t[3] ? t[47] : t[46];
  assign t[45] = ~(t[6] & t[62]);
  assign t[46] = ~(t[63]);
  assign t[47] = ~(t[8] & t[48]);
  assign t[48] = x[12] ? x[58] : t[64];
  assign t[49] = (t[65]);
  assign t[4] = ~(t[50]);
  assign t[50] = (t[66]);
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = t[81] ^ x[5];
  assign t[66] = t[82] ^ x[11];
  assign t[67] = t[83] ^ x[18];
  assign t[68] = t[84] ^ x[22];
  assign t[69] = t[85] ^ x[25];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[28];
  assign t[71] = t[87] ^ x[31];
  assign t[72] = t[88] ^ x[32];
  assign t[73] = t[89] ^ x[33];
  assign t[74] = t[90] ^ x[39];
  assign t[75] = t[91] ^ x[41];
  assign t[76] = t[92] ^ x[42];
  assign t[77] = t[93] ^ x[48];
  assign t[78] = t[94] ^ x[50];
  assign t[79] = t[95] ^ x[51];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[57];
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[109] & t[110]);
  assign t[88] = (~t[97] & t[111]);
  assign t[89] = (~t[99] & t[112]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[113] & t[114]);
  assign t[91] = (~t[97] & t[115]);
  assign t[92] = (~t[99] & t[116]);
  assign t[93] = (~t[117] & t[118]);
  assign t[94] = (~t[97] & t[119]);
  assign t[95] = (~t[99] & t[120]);
  assign t[96] = (~t[121] & t[122]);
  assign t[97] = t[123] ^ x[4];
  assign t[98] = t[124] ^ x[5];
  assign t[99] = t[125] ^ x[10];
  assign t[9] = x[12] ? x[19] : t[51];
  assign y = (t[0] & ~t[31] & ~t[37] & ~t[43]) | (~t[0] & t[31] & ~t[37] & ~t[43]) | (~t[0] & ~t[31] & t[37] & ~t[43]) | (~t[0] & ~t[31] & ~t[37] & t[43]) | (t[0] & t[31] & t[37] & ~t[43]) | (t[0] & t[31] & ~t[37] & t[43]) | (t[0] & ~t[31] & t[37] & t[43]) | (~t[0] & t[31] & t[37] & t[43]);
endmodule

module R2ind196(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[2]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[8]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[1]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [31:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[18];
  assign t[41] = t[48] ^ x[22];
  assign t[42] = t[49] ^ x[25];
  assign t[43] = t[50] ^ x[28];
  assign t[44] = t[51] ^ x[31];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[56] & t[57]);
  assign t[48] = (~t[58] & t[59]);
  assign t[49] = (~t[60] & t[61]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[62] & t[63]);
  assign t[51] = (~t[64] & t[65]);
  assign t[52] = t[66] ^ x[4];
  assign t[53] = t[67] ^ x[5];
  assign t[54] = t[68] ^ x[10];
  assign t[55] = t[69] ^ x[11];
  assign t[56] = t[70] ^ x[17];
  assign t[57] = t[71] ^ x[18];
  assign t[58] = t[72] ^ x[21];
  assign t[59] = t[73] ^ x[22];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[24];
  assign t[61] = t[75] ^ x[25];
  assign t[62] = t[76] ^ x[27];
  assign t[63] = t[77] ^ x[28];
  assign t[64] = t[78] ^ x[30];
  assign t[65] = t[79] ^ x[31];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[71] = (x[13]);
  assign t[72] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[20]);
  assign t[74] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[23]);
  assign t[76] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[26]);
  assign t[78] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[29]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[33];
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [46:0] x;
 output y;

 wire [137:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[18];
  assign t[101] = t[123] ^ x[19];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[26];
  assign t[107] = t[129] ^ x[27];
  assign t[108] = t[130] ^ x[29];
  assign t[109] = t[131] ^ x[30];
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = t[132] ^ x[35];
  assign t[111] = t[133] ^ x[36];
  assign t[112] = t[134] ^ x[38];
  assign t[113] = t[135] ^ x[39];
  assign t[114] = t[136] ^ x[44];
  assign t[115] = t[137] ^ x[45];
  assign t[116] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[117] = (x[0]);
  assign t[118] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[119] = (x[6]);
  assign t[11] = ~(t[15]);
  assign t[120] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[14]);
  assign t[122] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[17]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[1]);
  assign t[129] = (x[7]);
  assign t[12] = ~(t[16]);
  assign t[130] = (x[2]);
  assign t[131] = (x[8]);
  assign t[132] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[133] = (x[31]);
  assign t[134] = (x[3]);
  assign t[135] = (x[9]);
  assign t[136] = (x[40] & ~x[41] & ~x[42] & ~x[43]) | (~x[40] & x[41] & ~x[42] & ~x[43]) | (~x[40] & ~x[41] & x[42] & ~x[43]) | (~x[40] & ~x[41] & ~x[42] & x[43]) | (x[40] & x[41] & x[42] & ~x[43]) | (x[40] & x[41] & ~x[42] & x[43]) | (x[40] & ~x[41] & x[42] & x[43]) | (~x[40] & x[41] & x[42] & x[43]);
  assign t[137] = (x[40]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[13]);
  assign t[17] = ~(t[54] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[13]);
  assign t[21] = ~(t[55] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[56] | t[29]);
  assign t[25] = ~(t[56]);
  assign t[26] = t[30] & t[57];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[54] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[52]);
  assign t[30] = ~(t[54] | t[55]);
  assign t[31] = ~(t[55]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[13] ? x[28] : t[52];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[60]);
  assign t[42] = ~(t[61]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = t[12] ? x[37] : t[62];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[63]);
  assign t[48] = ~(t[64]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[53]);
  assign t[50] = t[51] ? x[46] : t[65];
  assign t[51] = ~(t[16]);
  assign t[52] = (t[66]);
  assign t[53] = (t[67]);
  assign t[54] = (t[68]);
  assign t[55] = (t[69]);
  assign t[56] = (t[70]);
  assign t[57] = (t[71]);
  assign t[58] = (t[72]);
  assign t[59] = (t[73]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[74]);
  assign t[61] = (t[75]);
  assign t[62] = (t[76]);
  assign t[63] = (t[77]);
  assign t[64] = (t[78]);
  assign t[65] = (t[79]);
  assign t[66] = t[80] ^ x[5];
  assign t[67] = t[81] ^ x[11];
  assign t[68] = t[82] ^ x[16];
  assign t[69] = t[83] ^ x[19];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[84] ^ x[22];
  assign t[71] = t[85] ^ x[25];
  assign t[72] = t[86] ^ x[26];
  assign t[73] = t[87] ^ x[27];
  assign t[74] = t[88] ^ x[29];
  assign t[75] = t[89] ^ x[30];
  assign t[76] = t[90] ^ x[36];
  assign t[77] = t[91] ^ x[38];
  assign t[78] = t[92] ^ x[39];
  assign t[79] = t[93] ^ x[45];
  assign t[7] = ~(t[10]);
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[94] & t[106]);
  assign t[87] = (~t[96] & t[107]);
  assign t[88] = (~t[94] & t[108]);
  assign t[89] = (~t[96] & t[109]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[110] & t[111]);
  assign t[91] = (~t[94] & t[112]);
  assign t[92] = (~t[96] & t[113]);
  assign t[93] = (~t[114] & t[115]);
  assign t[94] = t[116] ^ x[4];
  assign t[95] = t[117] ^ x[5];
  assign t[96] = t[118] ^ x[10];
  assign t[97] = t[119] ^ x[11];
  assign t[98] = t[120] ^ x[15];
  assign t[99] = t[121] ^ x[16];
  assign t[9] = t[12] ? x[12] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind201(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[12]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[19]);
  assign t[17] = ~(t[36] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[19]);
  assign t[21] = ~(t[37] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[38] | t[29]);
  assign t[25] = ~(t[38]);
  assign t[26] = t[30] & t[39];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[36] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[37]);
  assign t[32] = ~(t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[16];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[12] & ~x[13] & ~x[14] & ~x[15]) | (~x[12] & x[13] & ~x[14] & ~x[15]) | (~x[12] & ~x[13] & x[14] & ~x[15]) | (~x[12] & ~x[13] & ~x[14] & x[15]) | (x[12] & x[13] & x[14] & ~x[15]) | (x[12] & x[13] & ~x[14] & x[15]) | (x[12] & ~x[13] & x[14] & x[15]) | (~x[12] & x[13] & x[14] & x[15]);
  assign t[73] = (x[12]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[18] : t[35];
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [26:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[14]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(x[12]);
  assign t[19] = ~(t[35] & t[22]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[36] | t[27]);
  assign t[23] = ~(t[36]);
  assign t[24] = t[28] & t[37];
  assign t[25] = ~(t[23] & t[29]);
  assign t[26] = ~(t[34] & t[30]);
  assign t[27] = ~(t[30]);
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[35]);
  assign t[2] = ~(t[6] & t[31]);
  assign t[30] = ~(t[37]);
  assign t[31] = (t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = t[45] ^ x[5];
  assign t[39] = t[46] ^ x[11];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[13];
  assign t[41] = t[48] ^ x[17];
  assign t[42] = t[49] ^ x[20];
  assign t[43] = t[50] ^ x[23];
  assign t[44] = t[51] ^ x[26];
  assign t[45] = (~t[52] & t[53]);
  assign t[46] = (~t[54] & t[55]);
  assign t[47] = (~t[52] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[32]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = t[65] ^ x[4];
  assign t[53] = t[66] ^ x[5];
  assign t[54] = t[67] ^ x[10];
  assign t[55] = t[68] ^ x[11];
  assign t[56] = t[69] ^ x[13];
  assign t[57] = t[70] ^ x[16];
  assign t[58] = t[71] ^ x[17];
  assign t[59] = t[72] ^ x[19];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[20];
  assign t[61] = t[74] ^ x[22];
  assign t[62] = t[75] ^ x[23];
  assign t[63] = t[76] ^ x[25];
  assign t[64] = t[77] ^ x[26];
  assign t[65] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[66] = (x[1]);
  assign t[67] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[68] = (x[7]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[15]);
  assign t[72] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[18]);
  assign t[74] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[21]);
  assign t[76] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[33];
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [25:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(x[13]);
  assign t[17] = ~(t[35] | t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(x[13]);
  assign t[21] = ~(t[36] & t[24]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[37] | t[29]);
  assign t[25] = ~(t[37]);
  assign t[26] = t[30] & t[38];
  assign t[27] = ~(t[25] & t[31]);
  assign t[28] = ~(t[35] & t[32]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = ~(t[35] | t[36]);
  assign t[31] = ~(t[36]);
  assign t[32] = ~(t[38]);
  assign t[33] = (t[39]);
  assign t[34] = (t[40]);
  assign t[35] = (t[41]);
  assign t[36] = (t[42]);
  assign t[37] = (t[43]);
  assign t[38] = (t[44]);
  assign t[39] = t[45] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[46] ^ x[11];
  assign t[41] = t[47] ^ x[16];
  assign t[42] = t[48] ^ x[19];
  assign t[43] = t[49] ^ x[22];
  assign t[44] = t[50] ^ x[25];
  assign t[45] = (~t[51] & t[52]);
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = t[63] ^ x[4];
  assign t[52] = t[64] ^ x[5];
  assign t[53] = t[65] ^ x[10];
  assign t[54] = t[66] ^ x[11];
  assign t[55] = t[67] ^ x[15];
  assign t[56] = t[68] ^ x[16];
  assign t[57] = t[69] ^ x[18];
  assign t[58] = t[70] ^ x[19];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[24];
  assign t[62] = t[74] ^ x[25];
  assign t[63] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[64] = (x[0]);
  assign t[65] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[66] = (x[6]);
  assign t[67] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[14]);
  assign t[69] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[17]);
  assign t[71] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[20]);
  assign t[73] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[23]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = t[12] ? x[12] : t[34];
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind206(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind211(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [42:0] x;
 output y;

 wire [138:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[18];
  assign t[101] = t[123] ^ x[21];
  assign t[102] = t[124] ^ x[22];
  assign t[103] = t[125] ^ x[24];
  assign t[104] = t[126] ^ x[25];
  assign t[105] = t[127] ^ x[27];
  assign t[106] = t[128] ^ x[28];
  assign t[107] = t[129] ^ x[30];
  assign t[108] = t[130] ^ x[31];
  assign t[109] = t[131] ^ x[32];
  assign t[10] = ~(t[3]);
  assign t[110] = t[132] ^ x[33];
  assign t[111] = t[133] ^ x[34];
  assign t[112] = t[134] ^ x[36];
  assign t[113] = t[135] ^ x[37];
  assign t[114] = t[136] ^ x[38];
  assign t[115] = t[137] ^ x[40];
  assign t[116] = t[138] ^ x[41];
  assign t[117] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[118] = (x[0]);
  assign t[119] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[120] = (x[6]);
  assign t[121] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[122] = (x[14]);
  assign t[123] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[20]);
  assign t[125] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[23]);
  assign t[127] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[26]);
  assign t[129] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15]);
  assign t[130] = (x[29]);
  assign t[131] = (x[1]);
  assign t[132] = (x[7]);
  assign t[133] = (x[15]);
  assign t[134] = (x[2]);
  assign t[135] = (x[8]);
  assign t[136] = (x[16]);
  assign t[137] = (x[3]);
  assign t[138] = (x[9]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[53] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[55] | t[28]);
  assign t[24] = ~(t[55]);
  assign t[25] = t[29] & t[56];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[53] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[53] | t[54]);
  assign t[2] = ~(t[6] & t[50]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[56]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[57]);
  assign t[35] = ~(t[58]);
  assign t[36] = ~(t[8] & t[37]);
  assign t[37] = x[12] ? x[35] : t[59];
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[6] & t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = ~(t[8] & t[43]);
  assign t[43] = x[12] ? x[39] : t[62];
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[63]);
  assign t[47] = ~(t[64]);
  assign t[48] = ~(t[8] & t[49]);
  assign t[49] = x[12] ? x[42] : t[51];
  assign t[4] = ~(t[51]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = t[80] ^ x[5];
  assign t[66] = t[81] ^ x[11];
  assign t[67] = t[82] ^ x[18];
  assign t[68] = t[83] ^ x[22];
  assign t[69] = t[84] ^ x[25];
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = t[85] ^ x[28];
  assign t[71] = t[86] ^ x[31];
  assign t[72] = t[87] ^ x[32];
  assign t[73] = t[88] ^ x[33];
  assign t[74] = t[89] ^ x[34];
  assign t[75] = t[90] ^ x[36];
  assign t[76] = t[91] ^ x[37];
  assign t[77] = t[92] ^ x[38];
  assign t[78] = t[93] ^ x[40];
  assign t[79] = t[94] ^ x[41];
  assign t[7] = ~(t[11]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[95] & t[109]);
  assign t[88] = (~t[97] & t[110]);
  assign t[89] = (~t[99] & t[111]);
  assign t[8] = ~(t[12]);
  assign t[90] = (~t[95] & t[112]);
  assign t[91] = (~t[97] & t[113]);
  assign t[92] = (~t[99] & t[114]);
  assign t[93] = (~t[95] & t[115]);
  assign t[94] = (~t[97] & t[116]);
  assign t[95] = t[117] ^ x[4];
  assign t[96] = t[118] ^ x[5];
  assign t[97] = t[119] ^ x[10];
  assign t[98] = t[120] ^ x[11];
  assign t[99] = t[121] ^ x[17];
  assign t[9] = x[12] ? x[19] : t[52];
  assign y = (t[0] & ~t[32] & ~t[38] & ~t[44]) | (~t[0] & t[32] & ~t[38] & ~t[44]) | (~t[0] & ~t[32] & t[38] & ~t[44]) | (~t[0] & ~t[32] & ~t[38] & t[44]) | (t[0] & t[32] & t[38] & ~t[44]) | (t[0] & t[32] & ~t[38] & t[44]) | (t[0] & ~t[32] & t[38] & t[44]) | (~t[0] & t[32] & t[38] & t[44]);
endmodule

module R2ind216(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[13];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[20];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[55] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[13];
  assign t[58] = t[71] ^ x[16];
  assign t[59] = t[72] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[19];
  assign t[61] = t[74] ^ x[20];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[15]);
  assign t[73] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[18]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[14] : t[34];
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[8]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[16]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[7]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[15]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[14]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [42:0] x;
 output y;

 wire [138:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[18];
  assign t[101] = t[123] ^ x[21];
  assign t[102] = t[124] ^ x[22];
  assign t[103] = t[125] ^ x[24];
  assign t[104] = t[126] ^ x[25];
  assign t[105] = t[127] ^ x[27];
  assign t[106] = t[128] ^ x[28];
  assign t[107] = t[129] ^ x[30];
  assign t[108] = t[130] ^ x[31];
  assign t[109] = t[131] ^ x[32];
  assign t[10] = ~(t[3]);
  assign t[110] = t[132] ^ x[33];
  assign t[111] = t[133] ^ x[34];
  assign t[112] = t[134] ^ x[36];
  assign t[113] = t[135] ^ x[37];
  assign t[114] = t[136] ^ x[38];
  assign t[115] = t[137] ^ x[40];
  assign t[116] = t[138] ^ x[41];
  assign t[117] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[118] = (x[0]);
  assign t[119] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[120] = (x[6]);
  assign t[121] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[122] = (x[14]);
  assign t[123] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[20]);
  assign t[125] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[23]);
  assign t[127] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[26]);
  assign t[129] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15]);
  assign t[130] = (x[29]);
  assign t[131] = (x[1]);
  assign t[132] = (x[7]);
  assign t[133] = (x[15]);
  assign t[134] = (x[2]);
  assign t[135] = (x[8]);
  assign t[136] = (x[16]);
  assign t[137] = (x[3]);
  assign t[138] = (x[9]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[53] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[55] | t[28]);
  assign t[24] = ~(t[55]);
  assign t[25] = t[29] & t[56];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[53] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[53] | t[54]);
  assign t[2] = ~(t[6] & t[50]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[56]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[57]);
  assign t[35] = ~(t[58]);
  assign t[36] = ~(t[8] & t[37]);
  assign t[37] = x[12] ? x[35] : t[59];
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[6] & t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = ~(t[8] & t[43]);
  assign t[43] = x[12] ? x[39] : t[62];
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[63]);
  assign t[47] = ~(t[64]);
  assign t[48] = ~(t[8] & t[49]);
  assign t[49] = x[12] ? x[42] : t[51];
  assign t[4] = ~(t[51]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = t[80] ^ x[5];
  assign t[66] = t[81] ^ x[11];
  assign t[67] = t[82] ^ x[18];
  assign t[68] = t[83] ^ x[22];
  assign t[69] = t[84] ^ x[25];
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = t[85] ^ x[28];
  assign t[71] = t[86] ^ x[31];
  assign t[72] = t[87] ^ x[32];
  assign t[73] = t[88] ^ x[33];
  assign t[74] = t[89] ^ x[34];
  assign t[75] = t[90] ^ x[36];
  assign t[76] = t[91] ^ x[37];
  assign t[77] = t[92] ^ x[38];
  assign t[78] = t[93] ^ x[40];
  assign t[79] = t[94] ^ x[41];
  assign t[7] = ~(t[11]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[95] & t[109]);
  assign t[88] = (~t[97] & t[110]);
  assign t[89] = (~t[99] & t[111]);
  assign t[8] = ~(t[12]);
  assign t[90] = (~t[95] & t[112]);
  assign t[91] = (~t[97] & t[113]);
  assign t[92] = (~t[99] & t[114]);
  assign t[93] = (~t[95] & t[115]);
  assign t[94] = (~t[97] & t[116]);
  assign t[95] = t[117] ^ x[4];
  assign t[96] = t[118] ^ x[5];
  assign t[97] = t[119] ^ x[10];
  assign t[98] = t[120] ^ x[11];
  assign t[99] = t[121] ^ x[17];
  assign t[9] = x[12] ? x[19] : t[52];
  assign y = (t[0] & ~t[32] & ~t[38] & ~t[44]) | (~t[0] & t[32] & ~t[38] & ~t[44]) | (~t[0] & ~t[32] & t[38] & ~t[44]) | (~t[0] & ~t[32] & ~t[38] & t[44]) | (t[0] & t[32] & t[38] & ~t[44]) | (t[0] & t[32] & ~t[38] & t[44]) | (t[0] & ~t[32] & t[38] & t[44]) | (~t[0] & t[32] & t[38] & t[44]);
endmodule

module R2ind221(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[13];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[20];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[55] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[13];
  assign t[58] = t[71] ^ x[16];
  assign t[59] = t[72] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[19];
  assign t[61] = t[74] ^ x[20];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[15]);
  assign t[73] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[18]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[14] : t[34];
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[8]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[16]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[7]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[15]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[14]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [42:0] x;
 output y;

 wire [138:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[18];
  assign t[101] = t[123] ^ x[21];
  assign t[102] = t[124] ^ x[22];
  assign t[103] = t[125] ^ x[24];
  assign t[104] = t[126] ^ x[25];
  assign t[105] = t[127] ^ x[27];
  assign t[106] = t[128] ^ x[28];
  assign t[107] = t[129] ^ x[30];
  assign t[108] = t[130] ^ x[31];
  assign t[109] = t[131] ^ x[32];
  assign t[10] = ~(t[3]);
  assign t[110] = t[132] ^ x[33];
  assign t[111] = t[133] ^ x[34];
  assign t[112] = t[134] ^ x[36];
  assign t[113] = t[135] ^ x[37];
  assign t[114] = t[136] ^ x[38];
  assign t[115] = t[137] ^ x[40];
  assign t[116] = t[138] ^ x[41];
  assign t[117] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[118] = (x[0]);
  assign t[119] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[120] = (x[6]);
  assign t[121] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[122] = (x[14]);
  assign t[123] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[20]);
  assign t[125] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[23]);
  assign t[127] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[26]);
  assign t[129] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[15]);
  assign t[130] = (x[29]);
  assign t[131] = (x[1]);
  assign t[132] = (x[7]);
  assign t[133] = (x[15]);
  assign t[134] = (x[2]);
  assign t[135] = (x[8]);
  assign t[136] = (x[16]);
  assign t[137] = (x[3]);
  assign t[138] = (x[9]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[53] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[55] | t[28]);
  assign t[24] = ~(t[55]);
  assign t[25] = t[29] & t[56];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[53] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[53] | t[54]);
  assign t[2] = ~(t[6] & t[50]);
  assign t[30] = ~(t[54]);
  assign t[31] = ~(t[56]);
  assign t[32] = ~(t[33] & t[34]);
  assign t[33] = t[3] ? t[36] : t[35];
  assign t[34] = ~(t[6] & t[57]);
  assign t[35] = ~(t[58]);
  assign t[36] = ~(t[8] & t[37]);
  assign t[37] = x[12] ? x[35] : t[59];
  assign t[38] = ~(t[39] & t[40]);
  assign t[39] = t[3] ? t[42] : t[41];
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[6] & t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = ~(t[8] & t[43]);
  assign t[43] = x[12] ? x[39] : t[62];
  assign t[44] = ~(t[45] & t[46]);
  assign t[45] = t[3] ? t[48] : t[47];
  assign t[46] = ~(t[6] & t[63]);
  assign t[47] = ~(t[64]);
  assign t[48] = ~(t[8] & t[49]);
  assign t[49] = x[12] ? x[42] : t[51];
  assign t[4] = ~(t[51]);
  assign t[50] = (t[65]);
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = t[80] ^ x[5];
  assign t[66] = t[81] ^ x[11];
  assign t[67] = t[82] ^ x[18];
  assign t[68] = t[83] ^ x[22];
  assign t[69] = t[84] ^ x[25];
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = t[85] ^ x[28];
  assign t[71] = t[86] ^ x[31];
  assign t[72] = t[87] ^ x[32];
  assign t[73] = t[88] ^ x[33];
  assign t[74] = t[89] ^ x[34];
  assign t[75] = t[90] ^ x[36];
  assign t[76] = t[91] ^ x[37];
  assign t[77] = t[92] ^ x[38];
  assign t[78] = t[93] ^ x[40];
  assign t[79] = t[94] ^ x[41];
  assign t[7] = ~(t[11]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = (~t[95] & t[109]);
  assign t[88] = (~t[97] & t[110]);
  assign t[89] = (~t[99] & t[111]);
  assign t[8] = ~(t[12]);
  assign t[90] = (~t[95] & t[112]);
  assign t[91] = (~t[97] & t[113]);
  assign t[92] = (~t[99] & t[114]);
  assign t[93] = (~t[95] & t[115]);
  assign t[94] = (~t[97] & t[116]);
  assign t[95] = t[117] ^ x[4];
  assign t[96] = t[118] ^ x[5];
  assign t[97] = t[119] ^ x[10];
  assign t[98] = t[120] ^ x[11];
  assign t[99] = t[121] ^ x[17];
  assign t[9] = x[12] ? x[19] : t[52];
  assign y = (t[0] & ~t[32] & ~t[38] & ~t[44]) | (~t[0] & t[32] & ~t[38] & ~t[44]) | (~t[0] & ~t[32] & t[38] & ~t[44]) | (~t[0] & ~t[32] & ~t[38] & t[44]) | (t[0] & t[32] & t[38] & ~t[44]) | (t[0] & t[32] & ~t[38] & t[44]) | (t[0] & ~t[32] & t[38] & t[44]) | (~t[0] & t[32] & t[38] & t[44]);
endmodule

module R2ind226(x, y);
 input [26:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[13];
  assign t[42] = t[49] ^ x[17];
  assign t[43] = t[50] ^ x[20];
  assign t[44] = t[51] ^ x[23];
  assign t[45] = t[52] ^ x[26];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[55] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = t[66] ^ x[4];
  assign t[54] = t[67] ^ x[5];
  assign t[55] = t[68] ^ x[10];
  assign t[56] = t[69] ^ x[11];
  assign t[57] = t[70] ^ x[13];
  assign t[58] = t[71] ^ x[16];
  assign t[59] = t[72] ^ x[17];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[19];
  assign t[61] = t[74] ^ x[20];
  assign t[62] = t[75] ^ x[22];
  assign t[63] = t[76] ^ x[23];
  assign t[64] = t[77] ^ x[25];
  assign t[65] = t[78] ^ x[26];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[15]);
  assign t[73] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[18]);
  assign t[75] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[21]);
  assign t[77] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[24]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[14] : t[34];
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[2]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[8]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[16]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[1]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[7]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[15]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [31:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[3]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[15]);
  assign t[15] = ~(t[18] & t[19]);
  assign t[16] = ~(t[35] | t[20]);
  assign t[17] = ~(t[21]);
  assign t[18] = ~(t[22]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] & t[23]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[37] | t[28]);
  assign t[24] = ~(t[37]);
  assign t[25] = t[29] & t[38];
  assign t[26] = ~(t[24] & t[30]);
  assign t[27] = ~(t[35] & t[31]);
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[6] & t[32]);
  assign t[30] = ~(t[36]);
  assign t[31] = ~(t[38]);
  assign t[32] = (t[39]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = t[46] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[11];
  assign t[41] = t[48] ^ x[18];
  assign t[42] = t[49] ^ x[22];
  assign t[43] = t[50] ^ x[25];
  assign t[44] = t[51] ^ x[28];
  assign t[45] = t[52] ^ x[31];
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = (~t[59] & t[60]);
  assign t[4] = ~(t[33]);
  assign t[50] = (~t[61] & t[62]);
  assign t[51] = (~t[63] & t[64]);
  assign t[52] = (~t[65] & t[66]);
  assign t[53] = t[67] ^ x[4];
  assign t[54] = t[68] ^ x[5];
  assign t[55] = t[69] ^ x[10];
  assign t[56] = t[70] ^ x[11];
  assign t[57] = t[71] ^ x[17];
  assign t[58] = t[72] ^ x[18];
  assign t[59] = t[73] ^ x[21];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[22];
  assign t[61] = t[75] ^ x[24];
  assign t[62] = t[76] ^ x[25];
  assign t[63] = t[77] ^ x[27];
  assign t[64] = t[78] ^ x[28];
  assign t[65] = t[79] ^ x[30];
  assign t[66] = t[80] ^ x[31];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[10]);
  assign t[70] = (x[6]);
  assign t[71] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[72] = (x[14]);
  assign t[73] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[20]);
  assign t[75] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[23]);
  assign t[77] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[26]);
  assign t[79] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[29]);
  assign t[8] = ~(t[12]);
  assign t[9] = x[12] ? x[19] : t[34];
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind231(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind236(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind241(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [42:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[122] ^ x[17];
  assign t[101] = t[123] ^ x[18];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[24];
  assign t[105] = t[127] ^ x[25];
  assign t[106] = t[128] ^ x[27];
  assign t[107] = t[129] ^ x[28];
  assign t[108] = t[130] ^ x[30];
  assign t[109] = t[131] ^ x[31];
  assign t[10] = ~(t[12]);
  assign t[110] = t[132] ^ x[32];
  assign t[111] = t[133] ^ x[33];
  assign t[112] = t[134] ^ x[34];
  assign t[113] = t[135] ^ x[36];
  assign t[114] = t[136] ^ x[37];
  assign t[115] = t[137] ^ x[38];
  assign t[116] = t[138] ^ x[40];
  assign t[117] = t[139] ^ x[41];
  assign t[118] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[119] = (x[0]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[121] = (x[6]);
  assign t[122] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[123] = (x[14]);
  assign t[124] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[20]);
  assign t[126] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[23]);
  assign t[128] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[26]);
  assign t[12] = ~(t[14]);
  assign t[130] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[29]);
  assign t[132] = (x[1]);
  assign t[133] = (x[7]);
  assign t[134] = (x[15]);
  assign t[135] = (x[2]);
  assign t[136] = (x[8]);
  assign t[137] = (x[16]);
  assign t[138] = (x[3]);
  assign t[139] = (x[9]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[54] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[54] & t[28]);
  assign t[24] = ~(t[55] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[55]);
  assign t[28] = ~(t[57]);
  assign t[29] = ~(t[56] | t[31]);
  assign t[2] = ~(t[6] & t[51]);
  assign t[30] = t[32] & t[57];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[54] | t[55]);
  assign t[33] = ~(t[34] & t[35]);
  assign t[34] = t[3] ? t[37] : t[36];
  assign t[35] = ~(t[6] & t[58]);
  assign t[36] = ~(t[59]);
  assign t[37] = ~(t[8] & t[38]);
  assign t[38] = x[12] ? x[35] : t[60];
  assign t[39] = ~(t[40] & t[41]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[3] ? t[43] : t[42];
  assign t[41] = ~(t[6] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[8] & t[44]);
  assign t[44] = x[12] ? x[39] : t[63];
  assign t[45] = ~(t[46] & t[47]);
  assign t[46] = t[3] ? t[49] : t[48];
  assign t[47] = ~(t[6] & t[64]);
  assign t[48] = ~(t[65]);
  assign t[49] = ~(t[8] & t[50]);
  assign t[4] = ~(t[52]);
  assign t[50] = x[12] ? x[42] : t[52];
  assign t[51] = (t[66]);
  assign t[52] = (t[67]);
  assign t[53] = (t[68]);
  assign t[54] = (t[69]);
  assign t[55] = (t[70]);
  assign t[56] = (t[71]);
  assign t[57] = (t[72]);
  assign t[58] = (t[73]);
  assign t[59] = (t[74]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[75]);
  assign t[61] = (t[76]);
  assign t[62] = (t[77]);
  assign t[63] = (t[78]);
  assign t[64] = (t[79]);
  assign t[65] = (t[80]);
  assign t[66] = t[81] ^ x[5];
  assign t[67] = t[82] ^ x[11];
  assign t[68] = t[83] ^ x[18];
  assign t[69] = t[84] ^ x[22];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[85] ^ x[25];
  assign t[71] = t[86] ^ x[28];
  assign t[72] = t[87] ^ x[31];
  assign t[73] = t[88] ^ x[32];
  assign t[74] = t[89] ^ x[33];
  assign t[75] = t[90] ^ x[34];
  assign t[76] = t[91] ^ x[36];
  assign t[77] = t[92] ^ x[37];
  assign t[78] = t[93] ^ x[38];
  assign t[79] = t[94] ^ x[40];
  assign t[7] = ~(t[10]);
  assign t[80] = t[95] ^ x[41];
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = (~t[96] & t[110]);
  assign t[89] = (~t[98] & t[111]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[100] & t[112]);
  assign t[91] = (~t[96] & t[113]);
  assign t[92] = (~t[98] & t[114]);
  assign t[93] = (~t[100] & t[115]);
  assign t[94] = (~t[96] & t[116]);
  assign t[95] = (~t[98] & t[117]);
  assign t[96] = t[118] ^ x[4];
  assign t[97] = t[119] ^ x[5];
  assign t[98] = t[120] ^ x[10];
  assign t[99] = t[121] ^ x[11];
  assign t[9] = x[12] ? x[19] : t[53];
  assign y = (t[0] & ~t[33] & ~t[39] & ~t[45]) | (~t[0] & t[33] & ~t[39] & ~t[45]) | (~t[0] & ~t[33] & t[39] & ~t[45]) | (~t[0] & ~t[33] & ~t[39] & t[45]) | (t[0] & t[33] & t[39] & ~t[45]) | (t[0] & t[33] & ~t[39] & t[45]) | (t[0] & ~t[33] & t[39] & t[45]) | (~t[0] & t[33] & t[39] & t[45]);
endmodule

module R2ind246(x, y);
 input [26:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[13];
  assign t[43] = t[50] ^ x[17];
  assign t[44] = t[51] ^ x[20];
  assign t[45] = t[52] ^ x[23];
  assign t[46] = t[53] ^ x[26];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[56] & t[58]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = (~t[61] & t[62]);
  assign t[52] = (~t[63] & t[64]);
  assign t[53] = (~t[65] & t[66]);
  assign t[54] = t[67] ^ x[4];
  assign t[55] = t[68] ^ x[5];
  assign t[56] = t[69] ^ x[10];
  assign t[57] = t[70] ^ x[11];
  assign t[58] = t[71] ^ x[13];
  assign t[59] = t[72] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[17];
  assign t[61] = t[74] ^ x[19];
  assign t[62] = t[75] ^ x[20];
  assign t[63] = t[76] ^ x[22];
  assign t[64] = t[77] ^ x[23];
  assign t[65] = t[78] ^ x[25];
  assign t[66] = t[79] ^ x[26];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[15]);
  assign t[74] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[18]);
  assign t[76] = (x[21] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[21] & 1'b0 & ~1'b0 & ~1'b0) | (~x[21] & ~1'b0 & 1'b0 & ~1'b0) | (~x[21] & ~1'b0 & ~1'b0 & 1'b0) | (x[21] & 1'b0 & 1'b0 & ~1'b0) | (x[21] & 1'b0 & ~1'b0 & 1'b0) | (x[21] & ~1'b0 & 1'b0 & 1'b0) | (~x[21] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[21]);
  assign t[78] = (x[24] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0 & ~1'b0) | (x[24] & 1'b0 & ~1'b0 & 1'b0) | (x[24] & ~1'b0 & 1'b0 & 1'b0) | (~x[24] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[24]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[14] : t[35];
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[2]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[8]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[16]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[1]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[7]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[15]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [31:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = ~(t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17] & t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(x[12]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[13]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[36] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[36] & t[28]);
  assign t[24] = ~(t[37] & t[29]);
  assign t[25] = ~(t[26] & t[30]);
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[37]);
  assign t[28] = ~(t[39]);
  assign t[29] = ~(t[38] | t[31]);
  assign t[2] = ~(t[6] & t[33]);
  assign t[30] = t[32] & t[39];
  assign t[31] = ~(t[28]);
  assign t[32] = ~(t[36] | t[37]);
  assign t[33] = (t[40]);
  assign t[34] = (t[41]);
  assign t[35] = (t[42]);
  assign t[36] = (t[43]);
  assign t[37] = (t[44]);
  assign t[38] = (t[45]);
  assign t[39] = (t[46]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[47] ^ x[5];
  assign t[41] = t[48] ^ x[11];
  assign t[42] = t[49] ^ x[18];
  assign t[43] = t[50] ^ x[22];
  assign t[44] = t[51] ^ x[25];
  assign t[45] = t[52] ^ x[28];
  assign t[46] = t[53] ^ x[31];
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[34]);
  assign t[50] = (~t[60] & t[61]);
  assign t[51] = (~t[62] & t[63]);
  assign t[52] = (~t[64] & t[65]);
  assign t[53] = (~t[66] & t[67]);
  assign t[54] = t[68] ^ x[4];
  assign t[55] = t[69] ^ x[5];
  assign t[56] = t[70] ^ x[10];
  assign t[57] = t[71] ^ x[11];
  assign t[58] = t[72] ^ x[17];
  assign t[59] = t[73] ^ x[18];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[74] ^ x[21];
  assign t[61] = t[75] ^ x[22];
  assign t[62] = t[76] ^ x[24];
  assign t[63] = t[77] ^ x[25];
  assign t[64] = t[78] ^ x[27];
  assign t[65] = t[79] ^ x[28];
  assign t[66] = t[80] ^ x[30];
  assign t[67] = t[81] ^ x[31];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[71] = (x[6]);
  assign t[72] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign t[73] = (x[14]);
  assign t[74] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[20]);
  assign t[76] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[23]);
  assign t[78] = (x[26] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[26] & 1'b0 & ~1'b0 & ~1'b0) | (~x[26] & ~1'b0 & 1'b0 & ~1'b0) | (~x[26] & ~1'b0 & ~1'b0 & 1'b0) | (x[26] & 1'b0 & 1'b0 & ~1'b0) | (x[26] & 1'b0 & ~1'b0 & 1'b0) | (x[26] & ~1'b0 & 1'b0 & 1'b0) | (~x[26] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[26]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[29]);
  assign t[8] = ~(t[11]);
  assign t[9] = x[12] ? x[19] : t[35];
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [51:0] x;
 output y;

 wire [194:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (t[119]);
  assign t[101] = (t[120]);
  assign t[102] = (t[121]);
  assign t[103] = t[122] ^ x[5];
  assign t[104] = t[123] ^ x[11];
  assign t[105] = t[124] ^ x[19];
  assign t[106] = t[125] ^ x[25];
  assign t[107] = t[126] ^ x[26];
  assign t[108] = t[127] ^ x[29];
  assign t[109] = t[128] ^ x[30];
  assign t[10] = ~(t[13]);
  assign t[110] = t[129] ^ x[31];
  assign t[111] = t[130] ^ x[32];
  assign t[112] = t[131] ^ x[33];
  assign t[113] = t[132] ^ x[34];
  assign t[114] = t[133] ^ x[37];
  assign t[115] = t[134] ^ x[40];
  assign t[116] = t[135] ^ x[43];
  assign t[117] = t[136] ^ x[44];
  assign t[118] = t[137] ^ x[45];
  assign t[119] = t[138] ^ x[46];
  assign t[11] = ~(t[14]);
  assign t[120] = t[139] ^ x[48];
  assign t[121] = t[140] ^ x[50];
  assign t[122] = (~t[141] & t[142]);
  assign t[123] = (~t[143] & t[144]);
  assign t[124] = (~t[145] & t[146]);
  assign t[125] = (~t[147] & t[148]);
  assign t[126] = (~t[145] & t[149]);
  assign t[127] = (~t[150] & t[151]);
  assign t[128] = (~t[143] & t[152]);
  assign t[129] = (~t[147] & t[153]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = (~t[145] & t[154]);
  assign t[131] = (~t[143] & t[155]);
  assign t[132] = (~t[147] & t[156]);
  assign t[133] = (~t[157] & t[158]);
  assign t[134] = (~t[159] & t[160]);
  assign t[135] = (~t[161] & t[162]);
  assign t[136] = (~t[143] & t[163]);
  assign t[137] = (~t[147] & t[164]);
  assign t[138] = (~t[141] & t[165]);
  assign t[139] = (~t[141] & t[166]);
  assign t[13] = ~(t[17]);
  assign t[140] = (~t[141] & t[167]);
  assign t[141] = t[168] ^ x[4];
  assign t[142] = t[169] ^ x[5];
  assign t[143] = t[170] ^ x[10];
  assign t[144] = t[171] ^ x[11];
  assign t[145] = t[172] ^ x[18];
  assign t[146] = t[173] ^ x[19];
  assign t[147] = t[174] ^ x[24];
  assign t[148] = t[175] ^ x[25];
  assign t[149] = t[176] ^ x[26];
  assign t[14] = ~(t[18] & t[19]);
  assign t[150] = t[177] ^ x[28];
  assign t[151] = t[178] ^ x[29];
  assign t[152] = t[179] ^ x[30];
  assign t[153] = t[180] ^ x[31];
  assign t[154] = t[181] ^ x[32];
  assign t[155] = t[182] ^ x[33];
  assign t[156] = t[183] ^ x[34];
  assign t[157] = t[184] ^ x[36];
  assign t[158] = t[185] ^ x[37];
  assign t[159] = t[186] ^ x[39];
  assign t[15] = t[20] ? t[22] : t[21];
  assign t[160] = t[187] ^ x[40];
  assign t[161] = t[188] ^ x[42];
  assign t[162] = t[189] ^ x[43];
  assign t[163] = t[190] ^ x[44];
  assign t[164] = t[191] ^ x[45];
  assign t[165] = t[192] ^ x[46];
  assign t[166] = t[193] ^ x[48];
  assign t[167] = t[194] ^ x[50];
  assign t[168] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[169] = (x[0]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[170] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[171] = (x[6]);
  assign t[172] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[173] = (x[15]);
  assign t[174] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[175] = (x[20]);
  assign t[176] = (x[17]);
  assign t[177] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[178] = (x[27]);
  assign t[179] = (x[8]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[22]);
  assign t[181] = (x[16]);
  assign t[182] = (x[9]);
  assign t[183] = (x[23]);
  assign t[184] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[185] = (x[35]);
  assign t[186] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[187] = (x[38]);
  assign t[188] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[189] = (x[41]);
  assign t[18] = ~(t[27]);
  assign t[190] = (x[7]);
  assign t[191] = (x[21]);
  assign t[192] = (x[1]);
  assign t[193] = (x[2]);
  assign t[194] = (x[3]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[27] ? t[86] : t[28];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = ~(t[20] | t[33]);
  assign t[24] = ~(t[29]);
  assign t[25] = ~(t[34] | t[35]);
  assign t[26] = ~(t[14]);
  assign t[27] = ~(t[36] | t[37]);
  assign t[28] = t[85] ^ t[87];
  assign t[29] = t[27] ? t[88] : t[38];
  assign t[2] = ~(t[6] & t[84]);
  assign t[30] = ~(t[39] & t[31]);
  assign t[31] = ~(t[40]);
  assign t[32] = ~(t[39] & t[24]);
  assign t[33] = t[27] ? t[85] : t[41];
  assign t[34] = ~(t[89] | t[42]);
  assign t[35] = ~(t[43]);
  assign t[36] = ~(t[44] & t[45]);
  assign t[37] = ~(t[89] & t[46]);
  assign t[38] = t[90] ^ t[91];
  assign t[39] = ~(t[33]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[27] ? t[92] : t[47];
  assign t[41] = t[93] ^ t[94];
  assign t[42] = ~(t[95] & t[48]);
  assign t[43] = ~(t[44] & t[49]);
  assign t[44] = ~(t[96]);
  assign t[45] = ~(t[95]);
  assign t[46] = ~(t[97]);
  assign t[47] = t[98] ^ t[99];
  assign t[48] = ~(t[96] | t[50]);
  assign t[49] = t[51] & t[97];
  assign t[4] = ~(t[85]);
  assign t[50] = ~(t[46]);
  assign t[51] = ~(t[89] | t[95]);
  assign t[52] = ~(t[53] & t[54]);
  assign t[53] = t[3] ? t[56] : t[55];
  assign t[54] = ~(t[6] & t[100]);
  assign t[55] = ~(t[98]);
  assign t[56] = ~(t[8] & t[57]);
  assign t[57] = x[12] ? x[47] : t[58];
  assign t[58] = ~(t[59] & t[60]);
  assign t[59] = ~(t[61] & t[21]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = ~(t[62] & t[63]);
  assign t[61] = ~(t[40] | t[64]);
  assign t[62] = ~(t[23] | t[31]);
  assign t[63] = t[20] ? t[21] : t[29];
  assign t[64] = ~(t[65] | t[32]);
  assign t[65] = ~(t[20]);
  assign t[66] = ~(t[67] & t[68]);
  assign t[67] = t[3] ? t[70] : t[69];
  assign t[68] = ~(t[6] & t[101]);
  assign t[69] = ~(t[90]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = ~(t[8] & t[71]);
  assign t[71] = x[12] ? x[49] : t[72];
  assign t[72] = ~(t[73] | t[74]);
  assign t[73] = ~(t[62] | t[63]);
  assign t[74] = ~(t[31] | t[75]);
  assign t[75] = ~(t[20] ^ t[33]);
  assign t[76] = ~(t[77] & t[78]);
  assign t[77] = t[3] ? t[80] : t[79];
  assign t[78] = ~(t[6] & t[102]);
  assign t[79] = ~(t[93]);
  assign t[7] = ~(t[10]);
  assign t[80] = ~(t[8] & t[81]);
  assign t[81] = x[12] ? x[51] : t[82];
  assign t[82] = ~(t[83] ^ t[75]);
  assign t[83] = ~(t[31] | t[29]);
  assign t[84] = (t[103]);
  assign t[85] = (t[104]);
  assign t[86] = (t[105]);
  assign t[87] = (t[106]);
  assign t[88] = (t[107]);
  assign t[89] = (t[108]);
  assign t[8] = ~(t[11]);
  assign t[90] = (t[109]);
  assign t[91] = (t[110]);
  assign t[92] = (t[111]);
  assign t[93] = (t[112]);
  assign t[94] = (t[113]);
  assign t[95] = (t[114]);
  assign t[96] = (t[115]);
  assign t[97] = (t[116]);
  assign t[98] = (t[117]);
  assign t[99] = (t[118]);
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0] & ~t[52] & ~t[66] & ~t[76]) | (~t[0] & t[52] & ~t[66] & ~t[76]) | (~t[0] & ~t[52] & t[66] & ~t[76]) | (~t[0] & ~t[52] & ~t[66] & t[76]) | (t[0] & t[52] & t[66] & ~t[76]) | (t[0] & t[52] & ~t[66] & t[76]) | (t[0] & ~t[52] & t[66] & t[76]) | (~t[0] & t[52] & t[66] & t[76]);
endmodule

module R2ind251(x, y);
 input [45:0] x;
 output y;

 wire [140:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[124] ^ x[21];
  assign t[101] = t[125] ^ x[22];
  assign t[102] = t[126] ^ x[23];
  assign t[103] = t[127] ^ x[28];
  assign t[104] = t[128] ^ x[29];
  assign t[105] = t[129] ^ x[30];
  assign t[106] = t[130] ^ x[31];
  assign t[107] = t[131] ^ x[33];
  assign t[108] = t[132] ^ x[34];
  assign t[109] = t[133] ^ x[35];
  assign t[10] = ~(t[13]);
  assign t[110] = t[134] ^ x[36];
  assign t[111] = t[135] ^ x[38];
  assign t[112] = t[136] ^ x[39];
  assign t[113] = t[137] ^ x[41];
  assign t[114] = t[138] ^ x[42];
  assign t[115] = t[139] ^ x[44];
  assign t[116] = t[140] ^ x[45];
  assign t[117] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[118] = (x[3]);
  assign t[119] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[11] = ~(t[14]);
  assign t[120] = (x[9]);
  assign t[121] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[122] = (x[17]);
  assign t[123] = (x[15]);
  assign t[124] = (x[6]);
  assign t[125] = (x[16]);
  assign t[126] = (x[8]);
  assign t[127] = (x[24] & ~x[25] & ~x[26] & ~x[27]) | (~x[24] & x[25] & ~x[26] & ~x[27]) | (~x[24] & ~x[25] & x[26] & ~x[27]) | (~x[24] & ~x[25] & ~x[26] & x[27]) | (x[24] & x[25] & x[26] & ~x[27]) | (x[24] & x[25] & ~x[26] & x[27]) | (x[24] & ~x[25] & x[26] & x[27]) | (~x[24] & x[25] & x[26] & x[27]);
  assign t[128] = (x[26]);
  assign t[129] = (x[24]);
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = (x[27]);
  assign t[131] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[32]);
  assign t[133] = (x[7]);
  assign t[134] = (x[25]);
  assign t[135] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[136] = (x[37]);
  assign t[137] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[138] = (x[40]);
  assign t[139] = (x[43] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0 & ~1'b0) | (x[43] & 1'b0 & ~1'b0 & 1'b0) | (x[43] & ~1'b0 & 1'b0 & 1'b0) | (~x[43] & 1'b0 & 1'b0 & 1'b0);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[43]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[22] ^ t[23]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[27]);
  assign t[21] = t[26] ? t[47] : t[28];
  assign t[22] = t[26] ? t[48] : t[29];
  assign t[23] = t[26] ? t[49] : t[30];
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[14]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[26] ? t[50] : t[35];
  assign t[28] = t[51] ^ t[52];
  assign t[29] = t[49] ^ t[53];
  assign t[2] = ~(t[6] & t[45]);
  assign t[30] = t[46] ^ t[54];
  assign t[31] = ~(t[55] | t[36]);
  assign t[32] = ~(t[37]);
  assign t[33] = ~(t[38] & t[39]);
  assign t[34] = ~(t[55] & t[40]);
  assign t[35] = t[56] ^ t[57];
  assign t[36] = ~(t[58] & t[41]);
  assign t[37] = ~(t[38] & t[42]);
  assign t[38] = ~(t[59]);
  assign t[39] = ~(t[58]);
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[59] | t[43]);
  assign t[42] = t[44] & t[60];
  assign t[43] = ~(t[40]);
  assign t[44] = ~(t[55] | t[58]);
  assign t[45] = (t[61]);
  assign t[46] = (t[62]);
  assign t[47] = (t[63]);
  assign t[48] = (t[64]);
  assign t[49] = (t[65]);
  assign t[4] = ~(t[46]);
  assign t[50] = (t[66]);
  assign t[51] = (t[67]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = t[77] ^ x[5];
  assign t[62] = t[78] ^ x[11];
  assign t[63] = t[79] ^ x[19];
  assign t[64] = t[80] ^ x[20];
  assign t[65] = t[81] ^ x[21];
  assign t[66] = t[82] ^ x[22];
  assign t[67] = t[83] ^ x[23];
  assign t[68] = t[84] ^ x[29];
  assign t[69] = t[85] ^ x[30];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[31];
  assign t[71] = t[87] ^ x[34];
  assign t[72] = t[88] ^ x[35];
  assign t[73] = t[89] ^ x[36];
  assign t[74] = t[90] ^ x[39];
  assign t[75] = t[91] ^ x[42];
  assign t[76] = t[92] ^ x[45];
  assign t[77] = (~t[93] & t[94]);
  assign t[78] = (~t[95] & t[96]);
  assign t[79] = (~t[97] & t[98]);
  assign t[7] = ~(t[10]);
  assign t[80] = (~t[97] & t[99]);
  assign t[81] = (~t[95] & t[100]);
  assign t[82] = (~t[97] & t[101]);
  assign t[83] = (~t[95] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[103] & t[105]);
  assign t[86] = (~t[103] & t[106]);
  assign t[87] = (~t[107] & t[108]);
  assign t[88] = (~t[95] & t[109]);
  assign t[89] = (~t[103] & t[110]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[111] & t[112]);
  assign t[91] = (~t[113] & t[114]);
  assign t[92] = (~t[115] & t[116]);
  assign t[93] = t[117] ^ x[4];
  assign t[94] = t[118] ^ x[5];
  assign t[95] = t[119] ^ x[10];
  assign t[96] = t[120] ^ x[11];
  assign t[97] = t[121] ^ x[18];
  assign t[98] = t[122] ^ x[19];
  assign t[99] = t[123] ^ x[20];
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [45:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[124] ^ x[4];
  assign t[101] = t[125] ^ x[5];
  assign t[102] = t[126] ^ x[10];
  assign t[103] = t[127] ^ x[11];
  assign t[104] = t[128] ^ x[18];
  assign t[105] = t[129] ^ x[19];
  assign t[106] = t[130] ^ x[20];
  assign t[107] = t[131] ^ x[21];
  assign t[108] = t[132] ^ x[22];
  assign t[109] = t[133] ^ x[24];
  assign t[10] = ~(t[13]);
  assign t[110] = t[134] ^ x[25];
  assign t[111] = t[135] ^ x[30];
  assign t[112] = t[136] ^ x[31];
  assign t[113] = t[137] ^ x[32];
  assign t[114] = t[138] ^ x[33];
  assign t[115] = t[139] ^ x[34];
  assign t[116] = t[140] ^ x[35];
  assign t[117] = t[141] ^ x[36];
  assign t[118] = t[142] ^ x[38];
  assign t[119] = t[143] ^ x[39];
  assign t[11] = ~(t[14]);
  assign t[120] = t[144] ^ x[41];
  assign t[121] = t[145] ^ x[42];
  assign t[122] = t[146] ^ x[44];
  assign t[123] = t[147] ^ x[45];
  assign t[124] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[125] = (x[2]);
  assign t[126] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[127] = (x[8]);
  assign t[128] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[129] = (x[15]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[130] = (x[17]);
  assign t[131] = (x[16]);
  assign t[132] = (x[6]);
  assign t[133] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[23]);
  assign t[135] = (x[26] & ~x[27] & ~x[28] & ~x[29]) | (~x[26] & x[27] & ~x[28] & ~x[29]) | (~x[26] & ~x[27] & x[28] & ~x[29]) | (~x[26] & ~x[27] & ~x[28] & x[29]) | (x[26] & x[27] & x[28] & ~x[29]) | (x[26] & x[27] & ~x[28] & x[29]) | (x[26] & ~x[27] & x[28] & x[29]) | (~x[26] & x[27] & x[28] & x[29]);
  assign t[136] = (x[26]);
  assign t[137] = (x[28]);
  assign t[138] = (x[7]);
  assign t[139] = (x[27]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[9]);
  assign t[141] = (x[29]);
  assign t[142] = (x[37] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[37] & 1'b0 & ~1'b0 & ~1'b0) | (~x[37] & ~1'b0 & 1'b0 & ~1'b0) | (~x[37] & ~1'b0 & ~1'b0 & 1'b0) | (x[37] & 1'b0 & 1'b0 & ~1'b0) | (x[37] & 1'b0 & ~1'b0 & 1'b0) | (x[37] & ~1'b0 & 1'b0 & 1'b0) | (~x[37] & 1'b0 & 1'b0 & 1'b0);
  assign t[143] = (x[37]);
  assign t[144] = (x[40] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0 & ~1'b0) | (x[40] & 1'b0 & ~1'b0 & 1'b0) | (x[40] & ~1'b0 & 1'b0 & 1'b0) | (~x[40] & 1'b0 & 1'b0 & 1'b0);
  assign t[145] = (x[40]);
  assign t[146] = (x[43] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[43] & 1'b0 & ~1'b0 & ~1'b0) | (~x[43] & ~1'b0 & 1'b0 & ~1'b0) | (~x[43] & ~1'b0 & ~1'b0 & 1'b0) | (x[43] & 1'b0 & 1'b0 & ~1'b0) | (x[43] & 1'b0 & ~1'b0 & 1'b0) | (x[43] & ~1'b0 & 1'b0 & 1'b0) | (~x[43] & 1'b0 & 1'b0 & 1'b0);
  assign t[147] = (x[43]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[22] | t[23]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[27] | t[22]);
  assign t[21] = t[28] ? t[30] : t[29];
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[28] ^ t[32]);
  assign t[24] = ~(t[33] | t[34]);
  assign t[25] = ~(t[14]);
  assign t[26] = ~(t[35] | t[36]);
  assign t[27] = ~(t[28] | t[32]);
  assign t[28] = t[26] ? t[54] : t[37];
  assign t[29] = t[26] ? t[55] : t[38];
  assign t[2] = ~(t[6] & t[52]);
  assign t[30] = ~(t[29] & t[39]);
  assign t[31] = t[26] ? t[56] : t[40];
  assign t[32] = t[26] ? t[57] : t[41];
  assign t[33] = ~(t[58] | t[42]);
  assign t[34] = ~(t[43]);
  assign t[35] = ~(t[44] & t[45]);
  assign t[36] = ~(t[58] & t[46]);
  assign t[37] = t[57] ^ t[59];
  assign t[38] = t[53] ^ t[60];
  assign t[39] = ~(t[47] & t[22]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] & t[48]);
  assign t[43] = ~(t[44] & t[49]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[65]);
  assign t[46] = ~(t[67]);
  assign t[47] = ~(t[32]);
  assign t[48] = ~(t[66] | t[50]);
  assign t[49] = t[51] & t[67];
  assign t[4] = ~(t[53]);
  assign t[50] = ~(t[46]);
  assign t[51] = ~(t[58] | t[65]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = (t[83]);
  assign t[68] = t[84] ^ x[5];
  assign t[69] = t[85] ^ x[11];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[19];
  assign t[71] = t[87] ^ x[20];
  assign t[72] = t[88] ^ x[21];
  assign t[73] = t[89] ^ x[22];
  assign t[74] = t[90] ^ x[25];
  assign t[75] = t[91] ^ x[31];
  assign t[76] = t[92] ^ x[32];
  assign t[77] = t[93] ^ x[33];
  assign t[78] = t[94] ^ x[34];
  assign t[79] = t[95] ^ x[35];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[36];
  assign t[81] = t[97] ^ x[39];
  assign t[82] = t[98] ^ x[42];
  assign t[83] = t[99] ^ x[45];
  assign t[84] = (~t[100] & t[101]);
  assign t[85] = (~t[102] & t[103]);
  assign t[86] = (~t[104] & t[105]);
  assign t[87] = (~t[104] & t[106]);
  assign t[88] = (~t[104] & t[107]);
  assign t[89] = (~t[102] & t[108]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[109] & t[110]);
  assign t[91] = (~t[111] & t[112]);
  assign t[92] = (~t[111] & t[113]);
  assign t[93] = (~t[102] & t[114]);
  assign t[94] = (~t[111] & t[115]);
  assign t[95] = (~t[102] & t[116]);
  assign t[96] = (~t[111] & t[117]);
  assign t[97] = (~t[118] & t[119]);
  assign t[98] = (~t[120] & t[121]);
  assign t[99] = (~t[122] & t[123]);
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [45:0] x;
 output y;

 wire [151:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (~t[122] & t[123]);
  assign t[101] = (~t[124] & t[125]);
  assign t[102] = (~t[106] & t[126]);
  assign t[103] = (~t[114] & t[127]);
  assign t[104] = t[128] ^ x[4];
  assign t[105] = t[129] ^ x[5];
  assign t[106] = t[130] ^ x[10];
  assign t[107] = t[131] ^ x[11];
  assign t[108] = t[132] ^ x[18];
  assign t[109] = t[133] ^ x[19];
  assign t[10] = ~(t[13]);
  assign t[110] = t[134] ^ x[20];
  assign t[111] = t[135] ^ x[21];
  assign t[112] = t[136] ^ x[23];
  assign t[113] = t[137] ^ x[24];
  assign t[114] = t[138] ^ x[29];
  assign t[115] = t[139] ^ x[30];
  assign t[116] = t[140] ^ x[31];
  assign t[117] = t[141] ^ x[32];
  assign t[118] = t[142] ^ x[33];
  assign t[119] = t[143] ^ x[34];
  assign t[11] = ~(t[14]);
  assign t[120] = t[144] ^ x[36];
  assign t[121] = t[145] ^ x[37];
  assign t[122] = t[146] ^ x[39];
  assign t[123] = t[147] ^ x[40];
  assign t[124] = t[148] ^ x[42];
  assign t[125] = t[149] ^ x[43];
  assign t[126] = t[150] ^ x[44];
  assign t[127] = t[151] ^ x[45];
  assign t[128] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[129] = (x[1]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[131] = (x[7]);
  assign t[132] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[133] = (x[16]);
  assign t[134] = (x[17]);
  assign t[135] = (x[15]);
  assign t[136] = (x[22] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[22] & 1'b0 & ~1'b0 & ~1'b0) | (~x[22] & ~1'b0 & 1'b0 & ~1'b0) | (~x[22] & ~1'b0 & ~1'b0 & 1'b0) | (x[22] & 1'b0 & 1'b0 & ~1'b0) | (x[22] & 1'b0 & ~1'b0 & 1'b0) | (x[22] & ~1'b0 & 1'b0 & 1'b0) | (~x[22] & 1'b0 & 1'b0 & 1'b0);
  assign t[137] = (x[22]);
  assign t[138] = (x[25] & ~x[26] & ~x[27] & ~x[28]) | (~x[25] & x[26] & ~x[27] & ~x[28]) | (~x[25] & ~x[26] & x[27] & ~x[28]) | (~x[25] & ~x[26] & ~x[27] & x[28]) | (x[25] & x[26] & x[27] & ~x[28]) | (x[25] & x[26] & ~x[27] & x[28]) | (x[25] & ~x[26] & x[27] & x[28]) | (~x[25] & x[26] & x[27] & x[28]);
  assign t[139] = (x[26]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[8]);
  assign t[141] = (x[27]);
  assign t[142] = (x[6]);
  assign t[143] = (x[25]);
  assign t[144] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[145] = (x[35]);
  assign t[146] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[147] = (x[38]);
  assign t[148] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[149] = (x[41]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[150] = (x[9]);
  assign t[151] = (x[28]);
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = t[33] ? t[21] : t[29];
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[14]);
  assign t[26] = ~(t[36] | t[37]);
  assign t[27] = t[26] ? t[58] : t[38];
  assign t[28] = ~(t[39] | t[40]);
  assign t[29] = t[26] ? t[59] : t[41];
  assign t[2] = ~(t[6] & t[56]);
  assign t[30] = ~(t[42] & t[32]);
  assign t[31] = ~(t[33] | t[43]);
  assign t[32] = ~(t[27]);
  assign t[33] = t[26] ? t[60] : t[44];
  assign t[34] = ~(t[61] | t[45]);
  assign t[35] = ~(t[46]);
  assign t[36] = ~(t[47] & t[48]);
  assign t[37] = ~(t[61] & t[49]);
  assign t[38] = t[57] ^ t[62];
  assign t[39] = ~(t[33]);
  assign t[3] = ~(t[7]);
  assign t[40] = ~(t[42] & t[50]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[43]);
  assign t[43] = t[26] ? t[65] : t[51];
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[67] & t[52]);
  assign t[46] = ~(t[47] & t[53]);
  assign t[47] = ~(t[68]);
  assign t[48] = ~(t[67]);
  assign t[49] = ~(t[69]);
  assign t[4] = ~(t[57]);
  assign t[50] = ~(t[29]);
  assign t[51] = t[70] ^ t[71];
  assign t[52] = ~(t[68] | t[54]);
  assign t[53] = t[55] & t[69];
  assign t[54] = ~(t[49]);
  assign t[55] = ~(t[61] | t[67]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = (t[83]);
  assign t[68] = (t[84]);
  assign t[69] = (t[85]);
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = (t[86]);
  assign t[71] = (t[87]);
  assign t[72] = t[88] ^ x[5];
  assign t[73] = t[89] ^ x[11];
  assign t[74] = t[90] ^ x[19];
  assign t[75] = t[91] ^ x[20];
  assign t[76] = t[92] ^ x[21];
  assign t[77] = t[93] ^ x[24];
  assign t[78] = t[94] ^ x[30];
  assign t[79] = t[95] ^ x[31];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[32];
  assign t[81] = t[97] ^ x[33];
  assign t[82] = t[98] ^ x[34];
  assign t[83] = t[99] ^ x[37];
  assign t[84] = t[100] ^ x[40];
  assign t[85] = t[101] ^ x[43];
  assign t[86] = t[102] ^ x[44];
  assign t[87] = t[103] ^ x[45];
  assign t[88] = (~t[104] & t[105]);
  assign t[89] = (~t[106] & t[107]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[108] & t[109]);
  assign t[91] = (~t[108] & t[110]);
  assign t[92] = (~t[108] & t[111]);
  assign t[93] = (~t[112] & t[113]);
  assign t[94] = (~t[114] & t[115]);
  assign t[95] = (~t[106] & t[116]);
  assign t[96] = (~t[114] & t[117]);
  assign t[97] = (~t[106] & t[118]);
  assign t[98] = (~t[114] & t[119]);
  assign t[99] = (~t[120] & t[121]);
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [45:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[124] ^ x[4];
  assign t[101] = t[125] ^ x[5];
  assign t[102] = t[126] ^ x[10];
  assign t[103] = t[127] ^ x[11];
  assign t[104] = t[128] ^ x[18];
  assign t[105] = t[129] ^ x[19];
  assign t[106] = t[130] ^ x[24];
  assign t[107] = t[131] ^ x[25];
  assign t[108] = t[132] ^ x[26];
  assign t[109] = t[133] ^ x[28];
  assign t[10] = ~(t[13]);
  assign t[110] = t[134] ^ x[29];
  assign t[111] = t[135] ^ x[30];
  assign t[112] = t[136] ^ x[31];
  assign t[113] = t[137] ^ x[32];
  assign t[114] = t[138] ^ x[33];
  assign t[115] = t[139] ^ x[34];
  assign t[116] = t[140] ^ x[36];
  assign t[117] = t[141] ^ x[37];
  assign t[118] = t[142] ^ x[39];
  assign t[119] = t[143] ^ x[40];
  assign t[11] = ~(t[14]);
  assign t[120] = t[144] ^ x[42];
  assign t[121] = t[145] ^ x[43];
  assign t[122] = t[146] ^ x[44];
  assign t[123] = t[147] ^ x[45];
  assign t[124] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[125] = (x[0]);
  assign t[126] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[127] = (x[6]);
  assign t[128] = (x[14] & ~x[15] & ~x[16] & ~x[17]) | (~x[14] & x[15] & ~x[16] & ~x[17]) | (~x[14] & ~x[15] & x[16] & ~x[17]) | (~x[14] & ~x[15] & ~x[16] & x[17]) | (x[14] & x[15] & x[16] & ~x[17]) | (x[14] & x[15] & ~x[16] & x[17]) | (x[14] & ~x[15] & x[16] & x[17]) | (~x[14] & x[15] & x[16] & x[17]);
  assign t[129] = (x[15]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[130] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[131] = (x[20]);
  assign t[132] = (x[17]);
  assign t[133] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[134] = (x[27]);
  assign t[135] = (x[8]);
  assign t[136] = (x[22]);
  assign t[137] = (x[16]);
  assign t[138] = (x[9]);
  assign t[139] = (x[23]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[141] = (x[35]);
  assign t[142] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[143] = (x[38]);
  assign t[144] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[145] = (x[41]);
  assign t[146] = (x[7]);
  assign t[147] = (x[21]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ? t[22] : t[21];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27]);
  assign t[19] = ~(x[12]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[27] ? t[54] : t[28];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = ~(t[20] | t[33]);
  assign t[24] = ~(t[29]);
  assign t[25] = ~(t[34] | t[35]);
  assign t[26] = ~(t[14]);
  assign t[27] = ~(t[36] | t[37]);
  assign t[28] = t[53] ^ t[55];
  assign t[29] = t[27] ? t[56] : t[38];
  assign t[2] = ~(t[6] & t[52]);
  assign t[30] = ~(t[39] & t[31]);
  assign t[31] = ~(t[40]);
  assign t[32] = ~(t[39] & t[24]);
  assign t[33] = t[27] ? t[53] : t[41];
  assign t[34] = ~(t[57] | t[42]);
  assign t[35] = ~(t[43]);
  assign t[36] = ~(t[44] & t[45]);
  assign t[37] = ~(t[57] & t[46]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = ~(t[33]);
  assign t[3] = ~(t[7]);
  assign t[40] = t[27] ? t[60] : t[47];
  assign t[41] = t[61] ^ t[62];
  assign t[42] = ~(t[63] & t[48]);
  assign t[43] = ~(t[44] & t[49]);
  assign t[44] = ~(t[64]);
  assign t[45] = ~(t[63]);
  assign t[46] = ~(t[65]);
  assign t[47] = t[66] ^ t[67];
  assign t[48] = ~(t[64] | t[50]);
  assign t[49] = t[51] & t[65];
  assign t[4] = ~(t[53]);
  assign t[50] = ~(t[46]);
  assign t[51] = ~(t[57] | t[63]);
  assign t[52] = (t[68]);
  assign t[53] = (t[69]);
  assign t[54] = (t[70]);
  assign t[55] = (t[71]);
  assign t[56] = (t[72]);
  assign t[57] = (t[73]);
  assign t[58] = (t[74]);
  assign t[59] = (t[75]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (t[76]);
  assign t[61] = (t[77]);
  assign t[62] = (t[78]);
  assign t[63] = (t[79]);
  assign t[64] = (t[80]);
  assign t[65] = (t[81]);
  assign t[66] = (t[82]);
  assign t[67] = (t[83]);
  assign t[68] = t[84] ^ x[5];
  assign t[69] = t[85] ^ x[11];
  assign t[6] = ~(t[8] | t[7]);
  assign t[70] = t[86] ^ x[19];
  assign t[71] = t[87] ^ x[25];
  assign t[72] = t[88] ^ x[26];
  assign t[73] = t[89] ^ x[29];
  assign t[74] = t[90] ^ x[30];
  assign t[75] = t[91] ^ x[31];
  assign t[76] = t[92] ^ x[32];
  assign t[77] = t[93] ^ x[33];
  assign t[78] = t[94] ^ x[34];
  assign t[79] = t[95] ^ x[37];
  assign t[7] = ~(t[10]);
  assign t[80] = t[96] ^ x[40];
  assign t[81] = t[97] ^ x[43];
  assign t[82] = t[98] ^ x[44];
  assign t[83] = t[99] ^ x[45];
  assign t[84] = (~t[100] & t[101]);
  assign t[85] = (~t[102] & t[103]);
  assign t[86] = (~t[104] & t[105]);
  assign t[87] = (~t[106] & t[107]);
  assign t[88] = (~t[104] & t[108]);
  assign t[89] = (~t[109] & t[110]);
  assign t[8] = ~(t[11]);
  assign t[90] = (~t[102] & t[111]);
  assign t[91] = (~t[106] & t[112]);
  assign t[92] = (~t[104] & t[113]);
  assign t[93] = (~t[102] & t[114]);
  assign t[94] = (~t[106] & t[115]);
  assign t[95] = (~t[116] & t[117]);
  assign t[96] = (~t[118] & t[119]);
  assign t[97] = (~t[120] & t[121]);
  assign t[98] = (~t[102] & t[122]);
  assign t[99] = (~t[106] & t[123]);
  assign t[9] = x[12] ? x[13] : t[12];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [513:0] x;
 output [254:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[30]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[30]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[14], x[13], x[12], x[30]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[14], x[13], x[12], x[30]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[36], x[35], x[34], x[30], x[42], x[41], x[40]}), .y(y[30]));
  R2ind31 R2ind31_inst(.y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[36], x[35], x[34], x[30], x[42], x[41], x[40]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[30], x[33], x[32], x[31], x[39], x[38], x[37]}), .y(y[35]));
  R2ind36 R2ind36_inst(.y(y[36]));
  R2ind37 R2ind37_inst(.y(y[37]));
  R2ind38 R2ind38_inst(.y(y[38]));
  R2ind39 R2ind39_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[30], x[33], x[32], x[31], x[39], x[38], x[37]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43], x[33], x[32], x[31]}), .y(y[40]));
  R2ind41 R2ind41_inst(.y(y[41]));
  R2ind42 R2ind42_inst(.y(y[42]));
  R2ind43 R2ind43_inst(.y(y[43]));
  R2ind44 R2ind44_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43], x[33], x[32], x[31]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43]}), .y(y[45]));
  R2ind46 R2ind46_inst(.y(y[46]));
  R2ind47 R2ind47_inst(.y(y[47]));
  R2ind48 R2ind48_inst(.y(y[48]));
  R2ind49 R2ind49_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[30], x[36], x[35], x[34]}), .y(y[50]));
  R2ind51 R2ind51_inst(.y(y[51]));
  R2ind52 R2ind52_inst(.y(y[52]));
  R2ind53 R2ind53_inst(.y(y[53]));
  R2ind54 R2ind54_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[30], x[36], x[35], x[34]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[26], x[25], x[24], x[30], x[29], x[28], x[27], x[20], x[19], x[18]}), .y(y[55]));
  R2ind56 R2ind56_inst(.y(y[56]));
  R2ind57 R2ind57_inst(.y(y[57]));
  R2ind58 R2ind58_inst(.y(y[58]));
  R2ind59 R2ind59_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[26], x[25], x[24], x[30], x[29], x[28], x[27], x[20], x[19], x[18]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[26], x[25], x[24], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[23], x[22], x[21]}), .y(y[60]));
  R2ind61 R2ind61_inst(.y(y[61]));
  R2ind62 R2ind62_inst(.y(y[62]));
  R2ind63 R2ind63_inst(.y(y[63]));
  R2ind64 R2ind64_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[26], x[25], x[24], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[23], x[22], x[21]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[26], x[25], x[24], x[29], x[28], x[27]}), .y(y[65]));
  R2ind66 R2ind66_inst(.y(y[66]));
  R2ind67 R2ind67_inst(.y(y[67]));
  R2ind68 R2ind68_inst(.y(y[68]));
  R2ind69 R2ind69_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[26], x[25], x[24], x[29], x[28], x[27]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[26], x[25], x[24]}), .y(y[70]));
  R2ind71 R2ind71_inst(.y(y[71]));
  R2ind72 R2ind72_inst(.y(y[72]));
  R2ind73 R2ind73_inst(.y(y[73]));
  R2ind74 R2ind74_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[26], x[25], x[24]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[14], x[13], x[12], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[17], x[16], x[15], x[11], x[10], x[9], x[30], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[8], x[7], x[6], x[52], x[51], x[50], x[49], x[48], x[47], x[46]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[78], x[77], x[64], x[58], x[73], x[75], x[74], x[70], x[14], x[13], x[12], x[71], x[69], x[68], x[67], x[66], x[65], x[17], x[16], x[15], x[11], x[10], x[9], x[30], x[76], x[63], x[62], x[61], x[60], x[59], x[72], x[57], x[56], x[55], x[54], x[53], x[8], x[7], x[6], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[50], x[49], x[48], x[47], x[46]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[64], x[58], x[76], x[72], x[75], x[74], x[71], x[70], x[73], x[69], x[68], x[67], x[66], x[65], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[30], x[78], x[63], x[62], x[61], x[60], x[59], x[77], x[57], x[56], x[55], x[54], x[53], x[8], x[7], x[6], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[50], x[49], x[48], x[47], x[46]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[64], x[58], x[78], x[77], x[76], x[72], x[73], x[70], x[71], x[69], x[68], x[67], x[66], x[65], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[30], x[75], x[63], x[62], x[61], x[60], x[59], x[74], x[57], x[56], x[55], x[54], x[53], x[8], x[7], x[6], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[50], x[49], x[48], x[47], x[46]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[78], x[77], x[76], x[75], x[74], x[73], x[14], x[13], x[12], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[17], x[16], x[15], x[11], x[10], x[9], x[30], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[8], x[7], x[6], x[52], x[51], x[50], x[49], x[48], x[47], x[46]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[85], x[51], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[79], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[87], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[84], x[83], x[82], x[81], x[80], x[95], x[50], x[49], x[48], x[47], x[46]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[85], x[84], x[83], x[82], x[81], x[80], x[51], x[50], x[49], x[48], x[47], x[46]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[84], x[83], x[82], x[81], x[80], x[79], x[50], x[49], x[48], x[47], x[46]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[84], x[83], x[82], x[81], x[80], x[87], x[50], x[49], x[48], x[47], x[46]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[84], x[83], x[82], x[81], x[80], x[95], x[50], x[49], x[48], x[47], x[46]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[93], x[85], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[119], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[111], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[92], x[91], x[90], x[89], x[88], x[103], x[84], x[83], x[82], x[81], x[80]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[93], x[92], x[91], x[90], x[89], x[88], x[85], x[84], x[83], x[82], x[81], x[80]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[92], x[91], x[90], x[89], x[88], x[119], x[84], x[83], x[82], x[81], x[80]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[92], x[91], x[90], x[89], x[88], x[111], x[84], x[83], x[82], x[81], x[80]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[92], x[91], x[90], x[89], x[88], x[103], x[84], x[83], x[82], x[81], x[80]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[101], x[93], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[150], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[142], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[166], x[64], x[63], x[62], x[61], x[60], x[59], x[165], x[100], x[99], x[98], x[97], x[96], x[134], x[92], x[91], x[90], x[89], x[88]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[101], x[100], x[99], x[98], x[97], x[96], x[93], x[92], x[91], x[90], x[89], x[88]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[100], x[99], x[98], x[97], x[96], x[150], x[92], x[91], x[90], x[89], x[88]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[100], x[99], x[98], x[97], x[96], x[142], x[92], x[91], x[90], x[89], x[88]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[166], x[64], x[63], x[62], x[61], x[60], x[59], x[165], x[100], x[99], x[98], x[97], x[96], x[134], x[92], x[91], x[90], x[89], x[88]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[196], x[79], x[50], x[49], x[48], x[47], x[46], x[132], x[101], x[195], x[119], x[84], x[83], x[82], x[81], x[80], x[194], x[193], x[150], x[92], x[91], x[90], x[89], x[88], x[192], x[167], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[191], x[175], x[190], x[131], x[130], x[129], x[128], x[127], x[165], x[100], x[99], x[98], x[97], x[96]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[196], x[79], x[50], x[49], x[48], x[47], x[46], x[132], x[131], x[130], x[129], x[128], x[127], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[195], x[119], x[84], x[83], x[82], x[81], x[80], x[194], x[131], x[130], x[129], x[128], x[127], x[175], x[100], x[99], x[98], x[97], x[96]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[193], x[150], x[92], x[91], x[90], x[89], x[88], x[192], x[131], x[130], x[129], x[128], x[127], x[167], x[100], x[99], x[98], x[97], x[96]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[191], x[175], x[190], x[131], x[130], x[129], x[128], x[127], x[165], x[100], x[99], x[98], x[97], x[96]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[205], x[125], x[132], x[204], x[203], x[194], x[202], x[201], x[116], x[115], x[114], x[113], x[112], x[200], x[192], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[199], x[198], x[108], x[107], x[106], x[105], x[104], x[197], x[124], x[123], x[122], x[121], x[120], x[190], x[131], x[130], x[129], x[128], x[127]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[205], x[194], x[125], x[124], x[123], x[122], x[121], x[120], x[132], x[131], x[130], x[129], x[128], x[127]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[204], x[203], x[124], x[123], x[122], x[121], x[120], x[194], x[131], x[130], x[129], x[128], x[127]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[202], x[201], x[116], x[115], x[114], x[113], x[112], x[200], x[124], x[123], x[122], x[121], x[120], x[192], x[131], x[130], x[129], x[128], x[127]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[199], x[198], x[108], x[107], x[106], x[105], x[104], x[197], x[124], x[123], x[122], x[121], x[120], x[190], x[131], x[130], x[129], x[128], x[127]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[215], x[214], x[162], x[161], x[160], x[159], x[158], x[117], x[125], x[213], x[212], x[155], x[154], x[153], x[152], x[151], x[201], x[203], x[211], x[210], x[147], x[146], x[145], x[144], x[143], x[209], x[200], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[208], x[207], x[139], x[138], x[137], x[136], x[135], x[206], x[116], x[115], x[114], x[113], x[112], x[197], x[124], x[123], x[122], x[121], x[120]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[215], x[214], x[162], x[161], x[160], x[159], x[158], x[117], x[116], x[115], x[114], x[113], x[112], x[125], x[124], x[123], x[122], x[121], x[120]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[213], x[212], x[155], x[154], x[153], x[152], x[151], x[201], x[116], x[115], x[114], x[113], x[112], x[203], x[124], x[123], x[122], x[121], x[120]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[211], x[210], x[147], x[146], x[145], x[144], x[143], x[209], x[116], x[115], x[114], x[113], x[112], x[200], x[124], x[123], x[122], x[121], x[120]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[208], x[207], x[139], x[138], x[137], x[136], x[135], x[206], x[116], x[115], x[114], x[113], x[112], x[197], x[124], x[123], x[122], x[121], x[120]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[224], x[223], x[187], x[186], x[185], x[184], x[183], x[109], x[117], x[222], x[221], x[180], x[179], x[178], x[177], x[176], x[198], x[201], x[220], x[219], x[172], x[171], x[170], x[169], x[168], x[218], x[209], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[217], x[75], x[63], x[62], x[61], x[60], x[59], x[216], x[108], x[107], x[106], x[105], x[104], x[206], x[116], x[115], x[114], x[113], x[112]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[224], x[223], x[187], x[186], x[185], x[184], x[183], x[109], x[108], x[107], x[106], x[105], x[104], x[117], x[116], x[115], x[114], x[113], x[112]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[222], x[221], x[180], x[179], x[178], x[177], x[176], x[198], x[108], x[107], x[106], x[105], x[104], x[201], x[116], x[115], x[114], x[113], x[112]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[220], x[219], x[172], x[171], x[170], x[169], x[168], x[218], x[108], x[107], x[106], x[105], x[104], x[209], x[116], x[115], x[114], x[113], x[112]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[217], x[75], x[63], x[62], x[61], x[60], x[59], x[216], x[108], x[107], x[106], x[105], x[104], x[206], x[116], x[115], x[114], x[113], x[112]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[230], x[87], x[50], x[49], x[48], x[47], x[46], x[163], x[109], x[229], x[111], x[84], x[83], x[82], x[81], x[80], x[214], x[198], x[228], x[142], x[92], x[91], x[90], x[89], x[88], x[227], x[218], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[226], x[167], x[100], x[99], x[98], x[97], x[96], x[225], x[162], x[161], x[160], x[159], x[158], x[216], x[108], x[107], x[106], x[105], x[104]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[230], x[87], x[50], x[49], x[48], x[47], x[46], x[163], x[162], x[161], x[160], x[159], x[158], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[229], x[111], x[84], x[83], x[82], x[81], x[80], x[214], x[162], x[161], x[160], x[159], x[158], x[198], x[108], x[107], x[106], x[105], x[104]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[228], x[142], x[92], x[91], x[90], x[89], x[88], x[227], x[162], x[161], x[160], x[159], x[158], x[218], x[108], x[107], x[106], x[105], x[104]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[226], x[167], x[100], x[99], x[98], x[97], x[96], x[225], x[162], x[161], x[160], x[159], x[158], x[216], x[108], x[107], x[106], x[105], x[104]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[236], x[192], x[131], x[130], x[129], x[128], x[127], x[156], x[163], x[235], x[200], x[124], x[123], x[122], x[121], x[120], x[212], x[214], x[234], x[209], x[116], x[115], x[114], x[113], x[112], x[233], x[227], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[232], x[218], x[108], x[107], x[106], x[105], x[104], x[30], x[231], x[155], x[154], x[153], x[152], x[151], x[225], x[162], x[161], x[160], x[159], x[158]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[236], x[192], x[131], x[130], x[129], x[128], x[127], x[156], x[155], x[154], x[153], x[152], x[151], x[163], x[162], x[161], x[160], x[159], x[158]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[235], x[200], x[124], x[123], x[122], x[121], x[120], x[212], x[155], x[154], x[153], x[152], x[151], x[214], x[162], x[161], x[160], x[159], x[158]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[234], x[209], x[116], x[115], x[114], x[113], x[112], x[233], x[155], x[154], x[153], x[152], x[151], x[227], x[162], x[161], x[160], x[159], x[158]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[232], x[218], x[108], x[107], x[106], x[105], x[104], x[30], x[231], x[155], x[154], x[153], x[152], x[151], x[225], x[162], x[161], x[160], x[159], x[158]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[249], x[70], x[58], x[248], x[247], x[73], x[74], x[246], x[245], x[71], x[77], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[30], x[237], x[69], x[68], x[67], x[66], x[65], x[72], x[57], x[56], x[55], x[54], x[53]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[249], x[237], x[30], x[70], x[69], x[68], x[67], x[66], x[65], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[248], x[247], x[242], x[241], x[240], x[239], x[238], x[30], x[73], x[69], x[68], x[67], x[66], x[65], x[74], x[57], x[56], x[55], x[54], x[53]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[246], x[245], x[242], x[241], x[240], x[239], x[238], x[30], x[71], x[69], x[68], x[67], x[66], x[65], x[77], x[57], x[56], x[55], x[54], x[53]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[30], x[237], x[69], x[68], x[67], x[66], x[65], x[72], x[57], x[56], x[55], x[54], x[53]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[262], x[247], x[70], x[261], x[260], x[245], x[73], x[259], x[258], x[243], x[71], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[30], x[250], x[242], x[241], x[240], x[239], x[238], x[237], x[69], x[68], x[67], x[66], x[65]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[262], x[250], x[30], x[247], x[242], x[241], x[240], x[239], x[238], x[70], x[69], x[68], x[67], x[66], x[65]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[261], x[260], x[255], x[254], x[253], x[252], x[251], x[30], x[245], x[242], x[241], x[240], x[239], x[238], x[73], x[69], x[68], x[67], x[66], x[65]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[259], x[258], x[255], x[254], x[253], x[252], x[251], x[30], x[243], x[242], x[241], x[240], x[239], x[238], x[71], x[69], x[68], x[67], x[66], x[65]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[30], x[250], x[242], x[241], x[240], x[239], x[238], x[237], x[69], x[68], x[67], x[66], x[65]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[275], x[260], x[247], x[274], x[273], x[258], x[245], x[272], x[271], x[256], x[243], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[30], x[263], x[255], x[254], x[253], x[252], x[251], x[250], x[242], x[241], x[240], x[239], x[238]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[275], x[263], x[30], x[260], x[255], x[254], x[253], x[252], x[251], x[247], x[242], x[241], x[240], x[239], x[238]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[274], x[273], x[268], x[267], x[266], x[265], x[264], x[30], x[258], x[255], x[254], x[253], x[252], x[251], x[245], x[242], x[241], x[240], x[239], x[238]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[272], x[271], x[268], x[267], x[266], x[265], x[264], x[30], x[256], x[255], x[254], x[253], x[252], x[251], x[243], x[242], x[241], x[240], x[239], x[238]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[30], x[263], x[255], x[254], x[253], x[252], x[251], x[250], x[242], x[241], x[240], x[239], x[238]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[288], x[273], x[260], x[287], x[286], x[271], x[258], x[285], x[284], x[269], x[256], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[283], x[282], x[281], x[280], x[279], x[278], x[45], x[44], x[43], x[277], x[30], x[276], x[268], x[267], x[266], x[265], x[264], x[263], x[255], x[254], x[253], x[252], x[251]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[288], x[276], x[30], x[273], x[268], x[267], x[266], x[265], x[264], x[260], x[255], x[254], x[253], x[252], x[251]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[287], x[286], x[282], x[281], x[280], x[279], x[278], x[30], x[271], x[268], x[267], x[266], x[265], x[264], x[258], x[255], x[254], x[253], x[252], x[251]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[285], x[284], x[282], x[281], x[280], x[279], x[278], x[30], x[269], x[268], x[267], x[266], x[265], x[264], x[256], x[255], x[254], x[253], x[252], x[251]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[283], x[282], x[281], x[280], x[279], x[278], x[45], x[44], x[43], x[277], x[30], x[276], x[268], x[267], x[266], x[265], x[264], x[263], x[255], x[254], x[253], x[252], x[251]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[33], x[32], x[31], x[301], x[286], x[273], x[300], x[39], x[38], x[37], x[299], x[284], x[271], x[298], x[36], x[35], x[34], x[297], x[283], x[269], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[296], x[295], x[294], x[293], x[292], x[291], x[42], x[41], x[40], x[290], x[30], x[289], x[282], x[281], x[280], x[279], x[278], x[276], x[268], x[267], x[266], x[265], x[264]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[289], x[33], x[32], x[31], x[301], x[30], x[286], x[282], x[281], x[280], x[279], x[278], x[273], x[268], x[267], x[266], x[265], x[264]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[300], x[295], x[294], x[293], x[292], x[291], x[39], x[38], x[37], x[299], x[30], x[284], x[282], x[281], x[280], x[279], x[278], x[271], x[268], x[267], x[266], x[265], x[264]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[298], x[295], x[294], x[293], x[292], x[291], x[36], x[35], x[34], x[297], x[30], x[283], x[282], x[281], x[280], x[279], x[278], x[269], x[268], x[267], x[266], x[265], x[264]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[296], x[295], x[294], x[293], x[292], x[291], x[42], x[41], x[40], x[290], x[30], x[289], x[282], x[281], x[280], x[279], x[278], x[276], x[268], x[267], x[266], x[265], x[264]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[314], x[300], x[286], x[313], x[312], x[298], x[284], x[311], x[310], x[296], x[283], x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[30], x[302], x[295], x[294], x[293], x[292], x[291], x[289], x[282], x[281], x[280], x[279], x[278]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[314], x[302], x[30], x[300], x[295], x[294], x[293], x[292], x[291], x[286], x[282], x[281], x[280], x[279], x[278]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[313], x[312], x[307], x[306], x[305], x[304], x[303], x[30], x[298], x[295], x[294], x[293], x[292], x[291], x[284], x[282], x[281], x[280], x[279], x[278]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[311], x[310], x[307], x[306], x[305], x[304], x[303], x[30], x[296], x[295], x[294], x[293], x[292], x[291], x[283], x[282], x[281], x[280], x[279], x[278]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[30], x[302], x[295], x[294], x[293], x[292], x[291], x[289], x[282], x[281], x[280], x[279], x[278]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[327], x[312], x[300], x[326], x[325], x[310], x[298], x[324], x[323], x[308], x[296], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[30], x[315], x[307], x[306], x[305], x[304], x[303], x[302], x[295], x[294], x[293], x[292], x[291]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[327], x[315], x[30], x[312], x[307], x[306], x[305], x[304], x[303], x[300], x[295], x[294], x[293], x[292], x[291]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[326], x[325], x[320], x[319], x[318], x[317], x[316], x[30], x[310], x[307], x[306], x[305], x[304], x[303], x[298], x[295], x[294], x[293], x[292], x[291]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[324], x[323], x[320], x[319], x[318], x[317], x[316], x[30], x[308], x[307], x[306], x[305], x[304], x[303], x[296], x[295], x[294], x[293], x[292], x[291]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[30], x[315], x[307], x[306], x[305], x[304], x[303], x[302], x[295], x[294], x[293], x[292], x[291]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[340], x[325], x[312], x[339], x[338], x[323], x[310], x[337], x[336], x[321], x[308], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[30], x[328], x[320], x[319], x[318], x[317], x[316], x[315], x[307], x[306], x[305], x[304], x[303]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[340], x[328], x[30], x[325], x[320], x[319], x[318], x[317], x[316], x[312], x[307], x[306], x[305], x[304], x[303]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[339], x[338], x[333], x[332], x[331], x[330], x[329], x[30], x[323], x[320], x[319], x[318], x[317], x[316], x[310], x[307], x[306], x[305], x[304], x[303]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[337], x[336], x[333], x[332], x[331], x[330], x[329], x[30], x[321], x[320], x[319], x[318], x[317], x[316], x[308], x[307], x[306], x[305], x[304], x[303]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[30], x[328], x[320], x[319], x[318], x[317], x[316], x[315], x[307], x[306], x[305], x[304], x[303]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[353], x[338], x[325], x[352], x[351], x[336], x[323], x[350], x[349], x[334], x[321], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[30], x[341], x[333], x[332], x[331], x[330], x[329], x[328], x[320], x[319], x[318], x[317], x[316]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[353], x[341], x[30], x[338], x[333], x[332], x[331], x[330], x[329], x[325], x[320], x[319], x[318], x[317], x[316]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[352], x[351], x[346], x[345], x[344], x[343], x[342], x[30], x[336], x[333], x[332], x[331], x[330], x[329], x[323], x[320], x[319], x[318], x[317], x[316]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[350], x[349], x[346], x[345], x[344], x[343], x[342], x[30], x[334], x[333], x[332], x[331], x[330], x[329], x[321], x[320], x[319], x[318], x[317], x[316]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[348], x[347], x[346], x[345], x[344], x[343], x[342], x[30], x[341], x[333], x[332], x[331], x[330], x[329], x[328], x[320], x[319], x[318], x[317], x[316]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[366], x[351], x[338], x[365], x[364], x[349], x[336], x[363], x[362], x[347], x[334], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[30], x[354], x[346], x[345], x[344], x[343], x[342], x[341], x[333], x[332], x[331], x[330], x[329]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[366], x[354], x[30], x[351], x[346], x[345], x[344], x[343], x[342], x[338], x[333], x[332], x[331], x[330], x[329]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[365], x[364], x[359], x[358], x[357], x[356], x[355], x[30], x[349], x[346], x[345], x[344], x[343], x[342], x[336], x[333], x[332], x[331], x[330], x[329]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[363], x[362], x[359], x[358], x[357], x[356], x[355], x[30], x[347], x[346], x[345], x[344], x[343], x[342], x[334], x[333], x[332], x[331], x[330], x[329]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[30], x[354], x[346], x[345], x[344], x[343], x[342], x[341], x[333], x[332], x[331], x[330], x[329]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[373], x[227], x[162], x[161], x[160], x[159], x[158], x[148], x[156], x[372], x[210], x[212], x[371], x[370], x[233], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[369], x[368], x[139], x[138], x[137], x[136], x[135], x[30], x[367], x[147], x[146], x[145], x[144], x[143], x[231], x[155], x[154], x[153], x[152], x[151]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[373], x[227], x[162], x[161], x[160], x[159], x[158], x[30], x[148], x[147], x[146], x[145], x[144], x[143], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[372], x[233], x[210], x[147], x[146], x[145], x[144], x[143], x[212], x[155], x[154], x[153], x[152], x[151]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[371], x[370], x[147], x[146], x[145], x[144], x[143], x[233], x[155], x[154], x[153], x[152], x[151]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[369], x[368], x[139], x[138], x[137], x[136], x[135], x[30], x[367], x[147], x[146], x[145], x[144], x[143], x[231], x[155], x[154], x[153], x[152], x[151]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[381], x[380], x[187], x[186], x[185], x[184], x[183], x[140], x[148], x[379], x[378], x[180], x[179], x[178], x[177], x[176], x[207], x[210], x[377], x[376], x[172], x[171], x[170], x[169], x[168], x[368], x[370], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[375], x[78], x[63], x[62], x[61], x[60], x[59], x[374], x[139], x[138], x[137], x[136], x[135], x[367], x[147], x[146], x[145], x[144], x[143]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[381], x[380], x[187], x[186], x[185], x[184], x[183], x[30], x[140], x[139], x[138], x[137], x[136], x[135], x[148], x[147], x[146], x[145], x[144], x[143]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[379], x[378], x[180], x[179], x[178], x[177], x[176], x[30], x[207], x[139], x[138], x[137], x[136], x[135], x[210], x[147], x[146], x[145], x[144], x[143]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[377], x[376], x[172], x[171], x[170], x[169], x[168], x[368], x[139], x[138], x[137], x[136], x[135], x[370], x[147], x[146], x[145], x[144], x[143]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[11], x[10], x[9], x[8], x[7], x[6], x[375], x[78], x[63], x[62], x[61], x[60], x[59], x[374], x[139], x[138], x[137], x[136], x[135], x[367], x[147], x[146], x[145], x[144], x[143]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[386], x[95], x[50], x[49], x[48], x[47], x[46], x[188], x[140], x[385], x[103], x[84], x[83], x[82], x[81], x[80], x[223], x[207], x[384], x[134], x[92], x[91], x[90], x[89], x[88], x[380], x[368], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[383], x[165], x[100], x[99], x[98], x[97], x[96], x[30], x[382], x[187], x[186], x[185], x[184], x[183], x[374], x[139], x[138], x[137], x[136], x[135]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[386], x[95], x[50], x[49], x[48], x[47], x[46], x[188], x[187], x[186], x[185], x[184], x[183], x[140], x[139], x[138], x[137], x[136], x[135]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[385], x[103], x[84], x[83], x[82], x[81], x[80], x[223], x[187], x[186], x[185], x[184], x[183], x[207], x[139], x[138], x[137], x[136], x[135]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[384], x[134], x[92], x[91], x[90], x[89], x[88], x[380], x[187], x[186], x[185], x[184], x[183], x[368], x[139], x[138], x[137], x[136], x[135]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[383], x[165], x[100], x[99], x[98], x[97], x[96], x[30], x[382], x[187], x[186], x[185], x[184], x[183], x[374], x[139], x[138], x[137], x[136], x[135]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[391], x[190], x[131], x[130], x[129], x[128], x[127], x[181], x[188], x[390], x[197], x[124], x[123], x[122], x[121], x[120], x[221], x[223], x[389], x[206], x[116], x[115], x[114], x[113], x[112], x[378], x[380], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[388], x[216], x[108], x[107], x[106], x[105], x[104], x[30], x[387], x[180], x[179], x[178], x[177], x[176], x[382], x[187], x[186], x[185], x[184], x[183]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[391], x[190], x[131], x[130], x[129], x[128], x[127], x[30], x[181], x[180], x[179], x[178], x[177], x[176], x[188], x[187], x[186], x[185], x[184], x[183]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[390], x[197], x[124], x[123], x[122], x[121], x[120], x[30], x[221], x[180], x[179], x[178], x[177], x[176], x[223], x[187], x[186], x[185], x[184], x[183]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[389], x[206], x[116], x[115], x[114], x[113], x[112], x[30], x[378], x[180], x[179], x[178], x[177], x[176], x[380], x[187], x[186], x[185], x[184], x[183]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[388], x[216], x[108], x[107], x[106], x[105], x[104], x[30], x[387], x[180], x[179], x[178], x[177], x[176], x[382], x[187], x[186], x[185], x[184], x[183]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[396], x[225], x[162], x[161], x[160], x[159], x[158], x[173], x[181], x[395], x[231], x[155], x[154], x[153], x[152], x[151], x[219], x[221], x[394], x[367], x[147], x[146], x[145], x[144], x[143], x[376], x[378], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[393], x[374], x[139], x[138], x[137], x[136], x[135], x[30], x[392], x[172], x[171], x[170], x[169], x[168], x[387], x[180], x[179], x[178], x[177], x[176]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[396], x[225], x[162], x[161], x[160], x[159], x[158], x[30], x[173], x[172], x[171], x[170], x[169], x[168], x[181], x[180], x[179], x[178], x[177], x[176]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[395], x[231], x[155], x[154], x[153], x[152], x[151], x[30], x[219], x[172], x[171], x[170], x[169], x[168], x[221], x[180], x[179], x[178], x[177], x[176]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[394], x[367], x[147], x[146], x[145], x[144], x[143], x[30], x[376], x[172], x[171], x[170], x[169], x[168], x[378], x[180], x[179], x[178], x[177], x[176]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[393], x[374], x[139], x[138], x[137], x[136], x[135], x[30], x[392], x[172], x[171], x[170], x[169], x[168], x[387], x[180], x[179], x[178], x[177], x[176]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[400], x[382], x[187], x[186], x[185], x[184], x[183], x[64], x[173], x[399], x[387], x[180], x[179], x[178], x[177], x[176], x[75], x[219], x[398], x[78], x[376], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[397], x[76], x[63], x[62], x[61], x[60], x[59], x[392], x[172], x[171], x[170], x[169], x[168]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[400], x[382], x[187], x[186], x[185], x[184], x[183], x[64], x[63], x[62], x[61], x[60], x[59], x[173], x[172], x[171], x[170], x[169], x[168]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[399], x[387], x[180], x[179], x[178], x[177], x[176], x[75], x[63], x[62], x[61], x[60], x[59], x[219], x[172], x[171], x[170], x[169], x[168]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[398], x[392], x[30], x[78], x[63], x[62], x[61], x[60], x[59], x[376], x[172], x[171], x[170], x[169], x[168]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[30], x[397], x[76], x[63], x[62], x[61], x[60], x[59], x[392], x[172], x[171], x[170], x[169], x[168]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[413], x[364], x[351], x[412], x[411], x[362], x[349], x[410], x[409], x[360], x[347], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[30], x[401], x[359], x[358], x[357], x[356], x[355], x[354], x[346], x[345], x[344], x[343], x[342]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[413], x[401], x[30], x[364], x[359], x[358], x[357], x[356], x[355], x[351], x[346], x[345], x[344], x[343], x[342]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[412], x[411], x[406], x[405], x[404], x[403], x[402], x[30], x[362], x[359], x[358], x[357], x[356], x[355], x[349], x[346], x[345], x[344], x[343], x[342]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[410], x[409], x[406], x[405], x[404], x[403], x[402], x[30], x[360], x[359], x[358], x[357], x[356], x[355], x[347], x[346], x[345], x[344], x[343], x[342]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[30], x[401], x[359], x[358], x[357], x[356], x[355], x[354], x[346], x[345], x[344], x[343], x[342]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[426], x[411], x[364], x[425], x[424], x[409], x[362], x[423], x[422], x[407], x[360], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[30], x[414], x[406], x[405], x[404], x[403], x[402], x[401], x[359], x[358], x[357], x[356], x[355]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[426], x[414], x[30], x[411], x[406], x[405], x[404], x[403], x[402], x[364], x[359], x[358], x[357], x[356], x[355]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[425], x[424], x[419], x[418], x[417], x[416], x[415], x[30], x[409], x[406], x[405], x[404], x[403], x[402], x[362], x[359], x[358], x[357], x[356], x[355]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[423], x[422], x[419], x[418], x[417], x[416], x[415], x[30], x[407], x[406], x[405], x[404], x[403], x[402], x[360], x[359], x[358], x[357], x[356], x[355]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[30], x[414], x[406], x[405], x[404], x[403], x[402], x[401], x[359], x[358], x[357], x[356], x[355]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[439], x[424], x[411], x[438], x[437], x[422], x[409], x[436], x[435], x[420], x[407], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[30], x[427], x[419], x[418], x[417], x[416], x[415], x[414], x[406], x[405], x[404], x[403], x[402]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[439], x[427], x[30], x[424], x[419], x[418], x[417], x[416], x[415], x[411], x[406], x[405], x[404], x[403], x[402]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[438], x[437], x[432], x[431], x[430], x[429], x[428], x[30], x[422], x[419], x[418], x[417], x[416], x[415], x[409], x[406], x[405], x[404], x[403], x[402]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[436], x[435], x[432], x[431], x[430], x[429], x[428], x[30], x[420], x[419], x[418], x[417], x[416], x[415], x[407], x[406], x[405], x[404], x[403], x[402]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[30], x[427], x[419], x[418], x[417], x[416], x[415], x[414], x[406], x[405], x[404], x[403], x[402]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[452], x[437], x[424], x[451], x[450], x[435], x[422], x[449], x[448], x[433], x[420], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[30], x[440], x[432], x[431], x[430], x[429], x[428], x[427], x[419], x[418], x[417], x[416], x[415]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[452], x[440], x[30], x[437], x[432], x[431], x[430], x[429], x[428], x[424], x[419], x[418], x[417], x[416], x[415]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[451], x[450], x[445], x[444], x[443], x[442], x[441], x[30], x[435], x[432], x[431], x[430], x[429], x[428], x[422], x[419], x[418], x[417], x[416], x[415]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[449], x[448], x[445], x[444], x[443], x[442], x[441], x[30], x[433], x[432], x[431], x[430], x[429], x[428], x[420], x[419], x[418], x[417], x[416], x[415]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[30], x[440], x[432], x[431], x[430], x[429], x[428], x[427], x[419], x[418], x[417], x[416], x[415]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[465], x[450], x[437], x[464], x[463], x[448], x[435], x[462], x[461], x[446], x[433], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[460], x[459], x[458], x[457], x[456], x[455], x[454], x[30], x[453], x[445], x[444], x[443], x[442], x[441], x[440], x[432], x[431], x[430], x[429], x[428]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[465], x[453], x[30], x[450], x[445], x[444], x[443], x[442], x[441], x[437], x[432], x[431], x[430], x[429], x[428]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[464], x[463], x[458], x[457], x[456], x[455], x[454], x[30], x[448], x[445], x[444], x[443], x[442], x[441], x[435], x[432], x[431], x[430], x[429], x[428]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[462], x[461], x[458], x[457], x[456], x[455], x[454], x[30], x[446], x[445], x[444], x[443], x[442], x[441], x[433], x[432], x[431], x[430], x[429], x[428]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[460], x[459], x[458], x[457], x[456], x[455], x[454], x[30], x[453], x[445], x[444], x[443], x[442], x[441], x[440], x[432], x[431], x[430], x[429], x[428]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[478], x[463], x[450], x[477], x[476], x[461], x[448], x[475], x[474], x[459], x[446], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[473], x[472], x[471], x[470], x[469], x[468], x[467], x[30], x[466], x[458], x[457], x[456], x[455], x[454], x[453], x[445], x[444], x[443], x[442], x[441]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[478], x[466], x[30], x[463], x[458], x[457], x[456], x[455], x[454], x[450], x[445], x[444], x[443], x[442], x[441]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[477], x[476], x[471], x[470], x[469], x[468], x[467], x[30], x[461], x[458], x[457], x[456], x[455], x[454], x[448], x[445], x[444], x[443], x[442], x[441]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[475], x[474], x[471], x[470], x[469], x[468], x[467], x[30], x[459], x[458], x[457], x[456], x[455], x[454], x[446], x[445], x[444], x[443], x[442], x[441]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[473], x[472], x[471], x[470], x[469], x[468], x[467], x[30], x[466], x[458], x[457], x[456], x[455], x[454], x[453], x[445], x[444], x[443], x[442], x[441]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[491], x[476], x[463], x[490], x[489], x[474], x[461], x[488], x[487], x[472], x[459], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[30], x[479], x[471], x[470], x[469], x[468], x[467], x[466], x[458], x[457], x[456], x[455], x[454]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[491], x[479], x[30], x[476], x[471], x[470], x[469], x[468], x[467], x[463], x[458], x[457], x[456], x[455], x[454]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[490], x[489], x[484], x[483], x[482], x[481], x[480], x[30], x[474], x[471], x[470], x[469], x[468], x[467], x[461], x[458], x[457], x[456], x[455], x[454]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[488], x[487], x[484], x[483], x[482], x[481], x[480], x[30], x[472], x[471], x[470], x[469], x[468], x[467], x[459], x[458], x[457], x[456], x[455], x[454]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[30], x[479], x[471], x[470], x[469], x[468], x[467], x[466], x[458], x[457], x[456], x[455], x[454]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[504], x[489], x[476], x[503], x[502], x[487], x[474], x[501], x[500], x[485], x[472], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[30], x[492], x[484], x[483], x[482], x[481], x[480], x[479], x[471], x[470], x[469], x[468], x[467]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[504], x[492], x[30], x[489], x[484], x[483], x[482], x[481], x[480], x[476], x[471], x[470], x[469], x[468], x[467]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[503], x[502], x[497], x[496], x[495], x[494], x[493], x[30], x[487], x[484], x[483], x[482], x[481], x[480], x[474], x[471], x[470], x[469], x[468], x[467]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[501], x[500], x[497], x[496], x[495], x[494], x[493], x[30], x[485], x[484], x[483], x[482], x[481], x[480], x[472], x[471], x[470], x[469], x[468], x[467]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[30], x[492], x[484], x[483], x[482], x[481], x[480], x[479], x[471], x[470], x[469], x[468], x[467]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[509], x[502], x[489], x[508], x[58], x[500], x[487], x[507], x[74], x[498], x[485], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[506], x[77], x[57], x[56], x[55], x[54], x[53], x[30], x[505], x[497], x[496], x[495], x[494], x[493], x[492], x[484], x[483], x[482], x[481], x[480]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[509], x[505], x[30], x[502], x[497], x[496], x[495], x[494], x[493], x[489], x[484], x[483], x[482], x[481], x[480]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[508], x[58], x[57], x[56], x[55], x[54], x[53], x[30], x[500], x[497], x[496], x[495], x[494], x[493], x[487], x[484], x[483], x[482], x[481], x[480]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[507], x[74], x[57], x[56], x[55], x[54], x[53], x[30], x[498], x[497], x[496], x[495], x[494], x[493], x[485], x[484], x[483], x[482], x[481], x[480]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[506], x[77], x[57], x[56], x[55], x[54], x[53], x[30], x[505], x[497], x[496], x[495], x[494], x[493], x[492], x[484], x[483], x[482], x[481], x[480]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[513], x[502], x[512], x[500], x[511], x[498], x[78], x[77], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[64], x[58], x[73], x[75], x[74], x[8], x[7], x[6], x[70], x[76], x[63], x[62], x[61], x[60], x[59], x[71], x[69], x[68], x[67], x[66], x[65], x[510], x[30], x[72], x[57], x[56], x[55], x[54], x[53], x[505], x[497], x[496], x[495], x[494], x[493]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[78], x[77], x[8], x[7], x[6], x[64], x[76], x[75], x[63], x[62], x[61], x[60], x[59], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[513], x[30], x[58], x[57], x[56], x[55], x[54], x[53], x[502], x[497], x[496], x[495], x[494], x[493]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[64], x[58], x[78], x[77], x[75], x[76], x[63], x[62], x[61], x[60], x[59], x[8], x[7], x[6], x[72], x[73], x[70], x[71], x[69], x[68], x[67], x[66], x[65], x[512], x[30], x[74], x[57], x[56], x[55], x[54], x[53], x[500], x[497], x[496], x[495], x[494], x[493]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[64], x[58], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[76], x[72], x[75], x[74], x[78], x[63], x[62], x[61], x[60], x[59], x[8], x[7], x[6], x[71], x[70], x[73], x[69], x[68], x[67], x[66], x[65], x[511], x[30], x[77], x[57], x[56], x[55], x[54], x[53], x[498], x[497], x[496], x[495], x[494], x[493]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[78], x[77], x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[64], x[58], x[73], x[75], x[74], x[8], x[7], x[6], x[70], x[76], x[63], x[62], x[61], x[60], x[59], x[71], x[69], x[68], x[67], x[66], x[65], x[510], x[30], x[72], x[57], x[56], x[55], x[54], x[53], x[505], x[497], x[496], x[495], x[494], x[493]}), .y(y[254]));
endmodule

