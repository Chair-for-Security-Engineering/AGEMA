/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 12 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 13 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d4 (SI_s0, clk, SI_s1, SI_s2, SI_s3, SI_s4, Fresh, SO_s0, SO_s1, SO_s2, SO_s3, SO_s4);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [3:0] SI_s3 ;
    input [3:0] SI_s4 ;
    input [169:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    output [3:0] SO_s3 ;
    output [3:0] SO_s4 ;
    wire signal_15 ;
    wire signal_16 ;
    wire signal_17 ;
    wire signal_18 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_57 ;
    wire signal_58 ;
    wire signal_59 ;
    wire signal_60 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_69 ;
    wire signal_70 ;
    wire signal_71 ;
    wire signal_72 ;
    wire signal_77 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_85 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_113 ;
    wire signal_114 ;
    wire signal_115 ;
    wire signal_116 ;
    wire signal_117 ;
    wire signal_118 ;
    wire signal_119 ;
    wire signal_120 ;
    wire signal_121 ;
    wire signal_122 ;
    wire signal_123 ;
    wire signal_124 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_141 ;
    wire signal_142 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(1)) cell_23 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_72, signal_71, signal_70, signal_69, signal_34}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_24 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({signal_80, signal_79, signal_78, signal_77, signal_35}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_25 ( .a ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({signal_88, signal_87, signal_86, signal_85, signal_36}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_26 ( .a ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({signal_96, signal_95, signal_94, signal_93, signal_37}) ) ;

    /* cells in depth 1 */
    buf_clk cell_58 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_407 ) ) ;
    buf_clk cell_60 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_409 ) ) ;
    buf_clk cell_62 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( signal_411 ) ) ;
    buf_clk cell_64 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( signal_413 ) ) ;
    buf_clk cell_66 ( .C ( clk ), .D ( SI_s4[3] ), .Q ( signal_415 ) ) ;
    buf_clk cell_68 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_417 ) ) ;
    buf_clk cell_70 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_419 ) ) ;
    buf_clk cell_72 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( signal_421 ) ) ;
    buf_clk cell_74 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( signal_423 ) ) ;
    buf_clk cell_76 ( .C ( clk ), .D ( SI_s4[0] ), .Q ( signal_425 ) ) ;
    buf_clk cell_78 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_427 ) ) ;
    buf_clk cell_80 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_429 ) ) ;
    buf_clk cell_82 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( signal_431 ) ) ;
    buf_clk cell_84 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( signal_433 ) ) ;
    buf_clk cell_86 ( .C ( clk ), .D ( SI_s4[2] ), .Q ( signal_435 ) ) ;
    buf_clk cell_88 ( .C ( clk ), .D ( signal_34 ), .Q ( signal_437 ) ) ;
    buf_clk cell_90 ( .C ( clk ), .D ( signal_69 ), .Q ( signal_439 ) ) ;
    buf_clk cell_92 ( .C ( clk ), .D ( signal_70 ), .Q ( signal_441 ) ) ;
    buf_clk cell_94 ( .C ( clk ), .D ( signal_71 ), .Q ( signal_443 ) ) ;
    buf_clk cell_96 ( .C ( clk ), .D ( signal_72 ), .Q ( signal_445 ) ) ;
    buf_clk cell_98 ( .C ( clk ), .D ( signal_36 ), .Q ( signal_447 ) ) ;
    buf_clk cell_100 ( .C ( clk ), .D ( signal_85 ), .Q ( signal_449 ) ) ;
    buf_clk cell_102 ( .C ( clk ), .D ( signal_86 ), .Q ( signal_451 ) ) ;
    buf_clk cell_104 ( .C ( clk ), .D ( signal_87 ), .Q ( signal_453 ) ) ;
    buf_clk cell_106 ( .C ( clk ), .D ( signal_88 ), .Q ( signal_455 ) ) ;
    buf_clk cell_138 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_487 ) ) ;
    buf_clk cell_144 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_493 ) ) ;
    buf_clk cell_150 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( signal_499 ) ) ;
    buf_clk cell_156 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( signal_505 ) ) ;
    buf_clk cell_162 ( .C ( clk ), .D ( SI_s4[1] ), .Q ( signal_511 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_27 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_100, signal_99, signal_98, signal_97, signal_38}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_28 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({signal_104, signal_103, signal_102, signal_101, signal_39}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_29 ( .a ({signal_100, signal_99, signal_98, signal_97, signal_38}), .b ({signal_108, signal_107, signal_106, signal_105, signal_40}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_30 ( .a ({signal_104, signal_103, signal_102, signal_101, signal_39}), .b ({signal_112, signal_111, signal_110, signal_109, signal_41}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_31 ( .a ({signal_80, signal_79, signal_78, signal_77, signal_35}), .b ({signal_88, signal_87, signal_86, signal_85, signal_36}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({signal_116, signal_115, signal_114, signal_113, signal_42}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_32 ( .a ({signal_72, signal_71, signal_70, signal_69, signal_34}), .b ({signal_96, signal_95, signal_94, signal_93, signal_37}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_120, signal_119, signal_118, signal_117, signal_43}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_33 ( .a ({signal_80, signal_79, signal_78, signal_77, signal_35}), .b ({signal_96, signal_95, signal_94, signal_93, signal_37}), .clk ( clk ), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({signal_124, signal_123, signal_122, signal_121, signal_44}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_34 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({signal_80, signal_79, signal_78, signal_77, signal_35}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({signal_128, signal_127, signal_126, signal_125, signal_45}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_35 ( .a ({signal_72, signal_71, signal_70, signal_69, signal_34}), .b ({signal_80, signal_79, signal_78, signal_77, signal_35}), .clk ( clk ), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_132, signal_131, signal_130, signal_129, signal_46}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_36 ( .a ({signal_124, signal_123, signal_122, signal_121, signal_44}), .b ({signal_136, signal_135, signal_134, signal_133, signal_47}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_39 ( .a ({signal_416, signal_414, signal_412, signal_410, signal_408}), .b ({signal_116, signal_115, signal_114, signal_113, signal_42}), .c ({signal_148, signal_147, signal_146, signal_145, signal_16}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_40 ( .a ({signal_426, signal_424, signal_422, signal_420, signal_418}), .b ({signal_128, signal_127, signal_126, signal_125, signal_45}), .c ({signal_152, signal_151, signal_150, signal_149, signal_50}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) cell_41 ( .a ({signal_426, signal_424, signal_422, signal_420, signal_418}), .b ({signal_132, signal_131, signal_130, signal_129, signal_46}), .c ({signal_156, signal_155, signal_154, signal_153, signal_15}) ) ;
    buf_clk cell_59 ( .C ( clk ), .D ( signal_407 ), .Q ( signal_408 ) ) ;
    buf_clk cell_61 ( .C ( clk ), .D ( signal_409 ), .Q ( signal_410 ) ) ;
    buf_clk cell_63 ( .C ( clk ), .D ( signal_411 ), .Q ( signal_412 ) ) ;
    buf_clk cell_65 ( .C ( clk ), .D ( signal_413 ), .Q ( signal_414 ) ) ;
    buf_clk cell_67 ( .C ( clk ), .D ( signal_415 ), .Q ( signal_416 ) ) ;
    buf_clk cell_69 ( .C ( clk ), .D ( signal_417 ), .Q ( signal_418 ) ) ;
    buf_clk cell_71 ( .C ( clk ), .D ( signal_419 ), .Q ( signal_420 ) ) ;
    buf_clk cell_73 ( .C ( clk ), .D ( signal_421 ), .Q ( signal_422 ) ) ;
    buf_clk cell_75 ( .C ( clk ), .D ( signal_423 ), .Q ( signal_424 ) ) ;
    buf_clk cell_77 ( .C ( clk ), .D ( signal_425 ), .Q ( signal_426 ) ) ;
    buf_clk cell_79 ( .C ( clk ), .D ( signal_427 ), .Q ( signal_428 ) ) ;
    buf_clk cell_81 ( .C ( clk ), .D ( signal_429 ), .Q ( signal_430 ) ) ;
    buf_clk cell_83 ( .C ( clk ), .D ( signal_431 ), .Q ( signal_432 ) ) ;
    buf_clk cell_85 ( .C ( clk ), .D ( signal_433 ), .Q ( signal_434 ) ) ;
    buf_clk cell_87 ( .C ( clk ), .D ( signal_435 ), .Q ( signal_436 ) ) ;
    buf_clk cell_89 ( .C ( clk ), .D ( signal_437 ), .Q ( signal_438 ) ) ;
    buf_clk cell_91 ( .C ( clk ), .D ( signal_439 ), .Q ( signal_440 ) ) ;
    buf_clk cell_93 ( .C ( clk ), .D ( signal_441 ), .Q ( signal_442 ) ) ;
    buf_clk cell_95 ( .C ( clk ), .D ( signal_443 ), .Q ( signal_444 ) ) ;
    buf_clk cell_97 ( .C ( clk ), .D ( signal_445 ), .Q ( signal_446 ) ) ;
    buf_clk cell_99 ( .C ( clk ), .D ( signal_447 ), .Q ( signal_448 ) ) ;
    buf_clk cell_101 ( .C ( clk ), .D ( signal_449 ), .Q ( signal_450 ) ) ;
    buf_clk cell_103 ( .C ( clk ), .D ( signal_451 ), .Q ( signal_452 ) ) ;
    buf_clk cell_105 ( .C ( clk ), .D ( signal_453 ), .Q ( signal_454 ) ) ;
    buf_clk cell_107 ( .C ( clk ), .D ( signal_455 ), .Q ( signal_456 ) ) ;
    buf_clk cell_139 ( .C ( clk ), .D ( signal_487 ), .Q ( signal_488 ) ) ;
    buf_clk cell_145 ( .C ( clk ), .D ( signal_493 ), .Q ( signal_494 ) ) ;
    buf_clk cell_151 ( .C ( clk ), .D ( signal_499 ), .Q ( signal_500 ) ) ;
    buf_clk cell_157 ( .C ( clk ), .D ( signal_505 ), .Q ( signal_506 ) ) ;
    buf_clk cell_163 ( .C ( clk ), .D ( signal_511 ), .Q ( signal_512 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_108 ( .C ( clk ), .D ( signal_40 ), .Q ( signal_457 ) ) ;
    buf_clk cell_110 ( .C ( clk ), .D ( signal_105 ), .Q ( signal_459 ) ) ;
    buf_clk cell_112 ( .C ( clk ), .D ( signal_106 ), .Q ( signal_461 ) ) ;
    buf_clk cell_114 ( .C ( clk ), .D ( signal_107 ), .Q ( signal_463 ) ) ;
    buf_clk cell_116 ( .C ( clk ), .D ( signal_108 ), .Q ( signal_465 ) ) ;
    buf_clk cell_118 ( .C ( clk ), .D ( signal_448 ), .Q ( signal_467 ) ) ;
    buf_clk cell_120 ( .C ( clk ), .D ( signal_450 ), .Q ( signal_469 ) ) ;
    buf_clk cell_122 ( .C ( clk ), .D ( signal_452 ), .Q ( signal_471 ) ) ;
    buf_clk cell_124 ( .C ( clk ), .D ( signal_454 ), .Q ( signal_473 ) ) ;
    buf_clk cell_126 ( .C ( clk ), .D ( signal_456 ), .Q ( signal_475 ) ) ;
    buf_clk cell_128 ( .C ( clk ), .D ( signal_41 ), .Q ( signal_477 ) ) ;
    buf_clk cell_130 ( .C ( clk ), .D ( signal_109 ), .Q ( signal_479 ) ) ;
    buf_clk cell_132 ( .C ( clk ), .D ( signal_110 ), .Q ( signal_481 ) ) ;
    buf_clk cell_134 ( .C ( clk ), .D ( signal_111 ), .Q ( signal_483 ) ) ;
    buf_clk cell_136 ( .C ( clk ), .D ( signal_112 ), .Q ( signal_485 ) ) ;
    buf_clk cell_140 ( .C ( clk ), .D ( signal_488 ), .Q ( signal_489 ) ) ;
    buf_clk cell_146 ( .C ( clk ), .D ( signal_494 ), .Q ( signal_495 ) ) ;
    buf_clk cell_152 ( .C ( clk ), .D ( signal_500 ), .Q ( signal_501 ) ) ;
    buf_clk cell_158 ( .C ( clk ), .D ( signal_506 ), .Q ( signal_507 ) ) ;
    buf_clk cell_164 ( .C ( clk ), .D ( signal_512 ), .Q ( signal_513 ) ) ;
    buf_clk cell_208 ( .C ( clk ), .D ( signal_15 ), .Q ( signal_557 ) ) ;
    buf_clk cell_218 ( .C ( clk ), .D ( signal_153 ), .Q ( signal_567 ) ) ;
    buf_clk cell_228 ( .C ( clk ), .D ( signal_154 ), .Q ( signal_577 ) ) ;
    buf_clk cell_238 ( .C ( clk ), .D ( signal_155 ), .Q ( signal_587 ) ) ;
    buf_clk cell_248 ( .C ( clk ), .D ( signal_156 ), .Q ( signal_597 ) ) ;
    buf_clk cell_258 ( .C ( clk ), .D ( signal_16 ), .Q ( signal_607 ) ) ;
    buf_clk cell_268 ( .C ( clk ), .D ( signal_145 ), .Q ( signal_617 ) ) ;
    buf_clk cell_278 ( .C ( clk ), .D ( signal_146 ), .Q ( signal_627 ) ) ;
    buf_clk cell_288 ( .C ( clk ), .D ( signal_147 ), .Q ( signal_637 ) ) ;
    buf_clk cell_298 ( .C ( clk ), .D ( signal_148 ), .Q ( signal_647 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_37 ( .a ({signal_436, signal_434, signal_432, signal_430, signal_428}), .b ({signal_120, signal_119, signal_118, signal_117, signal_43}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({signal_140, signal_139, signal_138, signal_137, signal_48}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_38 ( .a ({signal_416, signal_414, signal_412, signal_410, signal_408}), .b ({signal_124, signal_123, signal_122, signal_121, signal_44}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({signal_144, signal_143, signal_142, signal_141, signal_49}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_42 ( .a ({signal_140, signal_139, signal_138, signal_137, signal_48}), .b ({signal_160, signal_159, signal_158, signal_157, signal_51}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_43 ( .a ({signal_144, signal_143, signal_142, signal_141, signal_49}), .b ({signal_164, signal_163, signal_162, signal_161, signal_52}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_44 ( .a ({signal_446, signal_444, signal_442, signal_440, signal_438}), .b ({signal_136, signal_135, signal_134, signal_133, signal_47}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_168, signal_167, signal_166, signal_165, signal_53}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_45 ( .a ({signal_456, signal_454, signal_452, signal_450, signal_448}), .b ({signal_152, signal_151, signal_150, signal_149, signal_50}), .clk ( clk ), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({signal_172, signal_171, signal_170, signal_169, signal_54}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_46 ( .a ({signal_172, signal_171, signal_170, signal_169, signal_54}), .b ({signal_176, signal_175, signal_174, signal_173, signal_55}) ) ;
    buf_clk cell_109 ( .C ( clk ), .D ( signal_457 ), .Q ( signal_458 ) ) ;
    buf_clk cell_111 ( .C ( clk ), .D ( signal_459 ), .Q ( signal_460 ) ) ;
    buf_clk cell_113 ( .C ( clk ), .D ( signal_461 ), .Q ( signal_462 ) ) ;
    buf_clk cell_115 ( .C ( clk ), .D ( signal_463 ), .Q ( signal_464 ) ) ;
    buf_clk cell_117 ( .C ( clk ), .D ( signal_465 ), .Q ( signal_466 ) ) ;
    buf_clk cell_119 ( .C ( clk ), .D ( signal_467 ), .Q ( signal_468 ) ) ;
    buf_clk cell_121 ( .C ( clk ), .D ( signal_469 ), .Q ( signal_470 ) ) ;
    buf_clk cell_123 ( .C ( clk ), .D ( signal_471 ), .Q ( signal_472 ) ) ;
    buf_clk cell_125 ( .C ( clk ), .D ( signal_473 ), .Q ( signal_474 ) ) ;
    buf_clk cell_127 ( .C ( clk ), .D ( signal_475 ), .Q ( signal_476 ) ) ;
    buf_clk cell_129 ( .C ( clk ), .D ( signal_477 ), .Q ( signal_478 ) ) ;
    buf_clk cell_131 ( .C ( clk ), .D ( signal_479 ), .Q ( signal_480 ) ) ;
    buf_clk cell_133 ( .C ( clk ), .D ( signal_481 ), .Q ( signal_482 ) ) ;
    buf_clk cell_135 ( .C ( clk ), .D ( signal_483 ), .Q ( signal_484 ) ) ;
    buf_clk cell_137 ( .C ( clk ), .D ( signal_485 ), .Q ( signal_486 ) ) ;
    buf_clk cell_141 ( .C ( clk ), .D ( signal_489 ), .Q ( signal_490 ) ) ;
    buf_clk cell_147 ( .C ( clk ), .D ( signal_495 ), .Q ( signal_496 ) ) ;
    buf_clk cell_153 ( .C ( clk ), .D ( signal_501 ), .Q ( signal_502 ) ) ;
    buf_clk cell_159 ( .C ( clk ), .D ( signal_507 ), .Q ( signal_508 ) ) ;
    buf_clk cell_165 ( .C ( clk ), .D ( signal_513 ), .Q ( signal_514 ) ) ;
    buf_clk cell_209 ( .C ( clk ), .D ( signal_557 ), .Q ( signal_558 ) ) ;
    buf_clk cell_219 ( .C ( clk ), .D ( signal_567 ), .Q ( signal_568 ) ) ;
    buf_clk cell_229 ( .C ( clk ), .D ( signal_577 ), .Q ( signal_578 ) ) ;
    buf_clk cell_239 ( .C ( clk ), .D ( signal_587 ), .Q ( signal_588 ) ) ;
    buf_clk cell_249 ( .C ( clk ), .D ( signal_597 ), .Q ( signal_598 ) ) ;
    buf_clk cell_259 ( .C ( clk ), .D ( signal_607 ), .Q ( signal_608 ) ) ;
    buf_clk cell_269 ( .C ( clk ), .D ( signal_617 ), .Q ( signal_618 ) ) ;
    buf_clk cell_279 ( .C ( clk ), .D ( signal_627 ), .Q ( signal_628 ) ) ;
    buf_clk cell_289 ( .C ( clk ), .D ( signal_637 ), .Q ( signal_638 ) ) ;
    buf_clk cell_299 ( .C ( clk ), .D ( signal_647 ), .Q ( signal_648 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_142 ( .C ( clk ), .D ( signal_490 ), .Q ( signal_491 ) ) ;
    buf_clk cell_148 ( .C ( clk ), .D ( signal_496 ), .Q ( signal_497 ) ) ;
    buf_clk cell_154 ( .C ( clk ), .D ( signal_502 ), .Q ( signal_503 ) ) ;
    buf_clk cell_160 ( .C ( clk ), .D ( signal_508 ), .Q ( signal_509 ) ) ;
    buf_clk cell_166 ( .C ( clk ), .D ( signal_514 ), .Q ( signal_515 ) ) ;
    buf_clk cell_178 ( .C ( clk ), .D ( signal_52 ), .Q ( signal_527 ) ) ;
    buf_clk cell_184 ( .C ( clk ), .D ( signal_161 ), .Q ( signal_533 ) ) ;
    buf_clk cell_190 ( .C ( clk ), .D ( signal_162 ), .Q ( signal_539 ) ) ;
    buf_clk cell_196 ( .C ( clk ), .D ( signal_163 ), .Q ( signal_545 ) ) ;
    buf_clk cell_202 ( .C ( clk ), .D ( signal_164 ), .Q ( signal_551 ) ) ;
    buf_clk cell_210 ( .C ( clk ), .D ( signal_558 ), .Q ( signal_559 ) ) ;
    buf_clk cell_220 ( .C ( clk ), .D ( signal_568 ), .Q ( signal_569 ) ) ;
    buf_clk cell_230 ( .C ( clk ), .D ( signal_578 ), .Q ( signal_579 ) ) ;
    buf_clk cell_240 ( .C ( clk ), .D ( signal_588 ), .Q ( signal_589 ) ) ;
    buf_clk cell_250 ( .C ( clk ), .D ( signal_598 ), .Q ( signal_599 ) ) ;
    buf_clk cell_260 ( .C ( clk ), .D ( signal_608 ), .Q ( signal_609 ) ) ;
    buf_clk cell_270 ( .C ( clk ), .D ( signal_618 ), .Q ( signal_619 ) ) ;
    buf_clk cell_280 ( .C ( clk ), .D ( signal_628 ), .Q ( signal_629 ) ) ;
    buf_clk cell_290 ( .C ( clk ), .D ( signal_638 ), .Q ( signal_639 ) ) ;
    buf_clk cell_300 ( .C ( clk ), .D ( signal_648 ), .Q ( signal_649 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_47 ( .a ({signal_466, signal_464, signal_462, signal_460, signal_458}), .b ({signal_168, signal_167, signal_166, signal_165, signal_53}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({signal_180, signal_179, signal_178, signal_177, signal_56}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_48 ( .a ({signal_476, signal_474, signal_472, signal_470, signal_468}), .b ({signal_160, signal_159, signal_158, signal_157, signal_51}), .clk ( clk ), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_184, signal_183, signal_182, signal_181, signal_57}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_49 ( .a ({signal_184, signal_183, signal_182, signal_181, signal_57}), .b ({signal_188, signal_187, signal_186, signal_185, signal_58}) ) ;
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_50 ( .a ({signal_176, signal_175, signal_174, signal_173, signal_55}), .b ({signal_486, signal_484, signal_482, signal_480, signal_478}), .clk ( clk ), .r ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .c ({signal_192, signal_191, signal_190, signal_189, signal_59}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_52 ( .a ({signal_192, signal_191, signal_190, signal_189, signal_59}), .b ({signal_200, signal_199, signal_198, signal_197, signal_17}) ) ;
    buf_clk cell_143 ( .C ( clk ), .D ( signal_491 ), .Q ( signal_492 ) ) ;
    buf_clk cell_149 ( .C ( clk ), .D ( signal_497 ), .Q ( signal_498 ) ) ;
    buf_clk cell_155 ( .C ( clk ), .D ( signal_503 ), .Q ( signal_504 ) ) ;
    buf_clk cell_161 ( .C ( clk ), .D ( signal_509 ), .Q ( signal_510 ) ) ;
    buf_clk cell_167 ( .C ( clk ), .D ( signal_515 ), .Q ( signal_516 ) ) ;
    buf_clk cell_179 ( .C ( clk ), .D ( signal_527 ), .Q ( signal_528 ) ) ;
    buf_clk cell_185 ( .C ( clk ), .D ( signal_533 ), .Q ( signal_534 ) ) ;
    buf_clk cell_191 ( .C ( clk ), .D ( signal_539 ), .Q ( signal_540 ) ) ;
    buf_clk cell_197 ( .C ( clk ), .D ( signal_545 ), .Q ( signal_546 ) ) ;
    buf_clk cell_203 ( .C ( clk ), .D ( signal_551 ), .Q ( signal_552 ) ) ;
    buf_clk cell_211 ( .C ( clk ), .D ( signal_559 ), .Q ( signal_560 ) ) ;
    buf_clk cell_221 ( .C ( clk ), .D ( signal_569 ), .Q ( signal_570 ) ) ;
    buf_clk cell_231 ( .C ( clk ), .D ( signal_579 ), .Q ( signal_580 ) ) ;
    buf_clk cell_241 ( .C ( clk ), .D ( signal_589 ), .Q ( signal_590 ) ) ;
    buf_clk cell_251 ( .C ( clk ), .D ( signal_599 ), .Q ( signal_600 ) ) ;
    buf_clk cell_261 ( .C ( clk ), .D ( signal_609 ), .Q ( signal_610 ) ) ;
    buf_clk cell_271 ( .C ( clk ), .D ( signal_619 ), .Q ( signal_620 ) ) ;
    buf_clk cell_281 ( .C ( clk ), .D ( signal_629 ), .Q ( signal_630 ) ) ;
    buf_clk cell_291 ( .C ( clk ), .D ( signal_639 ), .Q ( signal_640 ) ) ;
    buf_clk cell_301 ( .C ( clk ), .D ( signal_649 ), .Q ( signal_650 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_168 ( .C ( clk ), .D ( signal_58 ), .Q ( signal_517 ) ) ;
    buf_clk cell_170 ( .C ( clk ), .D ( signal_185 ), .Q ( signal_519 ) ) ;
    buf_clk cell_172 ( .C ( clk ), .D ( signal_186 ), .Q ( signal_521 ) ) ;
    buf_clk cell_174 ( .C ( clk ), .D ( signal_187 ), .Q ( signal_523 ) ) ;
    buf_clk cell_176 ( .C ( clk ), .D ( signal_188 ), .Q ( signal_525 ) ) ;
    buf_clk cell_180 ( .C ( clk ), .D ( signal_528 ), .Q ( signal_529 ) ) ;
    buf_clk cell_186 ( .C ( clk ), .D ( signal_534 ), .Q ( signal_535 ) ) ;
    buf_clk cell_192 ( .C ( clk ), .D ( signal_540 ), .Q ( signal_541 ) ) ;
    buf_clk cell_198 ( .C ( clk ), .D ( signal_546 ), .Q ( signal_547 ) ) ;
    buf_clk cell_204 ( .C ( clk ), .D ( signal_552 ), .Q ( signal_553 ) ) ;
    buf_clk cell_212 ( .C ( clk ), .D ( signal_560 ), .Q ( signal_561 ) ) ;
    buf_clk cell_222 ( .C ( clk ), .D ( signal_570 ), .Q ( signal_571 ) ) ;
    buf_clk cell_232 ( .C ( clk ), .D ( signal_580 ), .Q ( signal_581 ) ) ;
    buf_clk cell_242 ( .C ( clk ), .D ( signal_590 ), .Q ( signal_591 ) ) ;
    buf_clk cell_252 ( .C ( clk ), .D ( signal_600 ), .Q ( signal_601 ) ) ;
    buf_clk cell_262 ( .C ( clk ), .D ( signal_610 ), .Q ( signal_611 ) ) ;
    buf_clk cell_272 ( .C ( clk ), .D ( signal_620 ), .Q ( signal_621 ) ) ;
    buf_clk cell_282 ( .C ( clk ), .D ( signal_630 ), .Q ( signal_631 ) ) ;
    buf_clk cell_292 ( .C ( clk ), .D ( signal_640 ), .Q ( signal_641 ) ) ;
    buf_clk cell_302 ( .C ( clk ), .D ( signal_650 ), .Q ( signal_651 ) ) ;
    buf_clk cell_308 ( .C ( clk ), .D ( signal_17 ), .Q ( signal_657 ) ) ;
    buf_clk cell_314 ( .C ( clk ), .D ( signal_197 ), .Q ( signal_663 ) ) ;
    buf_clk cell_320 ( .C ( clk ), .D ( signal_198 ), .Q ( signal_669 ) ) ;
    buf_clk cell_326 ( .C ( clk ), .D ( signal_199 ), .Q ( signal_675 ) ) ;
    buf_clk cell_332 ( .C ( clk ), .D ( signal_200 ), .Q ( signal_681 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_51 ( .a ({signal_516, signal_510, signal_504, signal_498, signal_492}), .b ({signal_180, signal_179, signal_178, signal_177, signal_56}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .c ({signal_196, signal_195, signal_194, signal_193, signal_60}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_53 ( .a ({signal_196, signal_195, signal_194, signal_193, signal_60}), .b ({signal_204, signal_203, signal_202, signal_201, signal_61}) ) ;
    buf_clk cell_169 ( .C ( clk ), .D ( signal_517 ), .Q ( signal_518 ) ) ;
    buf_clk cell_171 ( .C ( clk ), .D ( signal_519 ), .Q ( signal_520 ) ) ;
    buf_clk cell_173 ( .C ( clk ), .D ( signal_521 ), .Q ( signal_522 ) ) ;
    buf_clk cell_175 ( .C ( clk ), .D ( signal_523 ), .Q ( signal_524 ) ) ;
    buf_clk cell_177 ( .C ( clk ), .D ( signal_525 ), .Q ( signal_526 ) ) ;
    buf_clk cell_181 ( .C ( clk ), .D ( signal_529 ), .Q ( signal_530 ) ) ;
    buf_clk cell_187 ( .C ( clk ), .D ( signal_535 ), .Q ( signal_536 ) ) ;
    buf_clk cell_193 ( .C ( clk ), .D ( signal_541 ), .Q ( signal_542 ) ) ;
    buf_clk cell_199 ( .C ( clk ), .D ( signal_547 ), .Q ( signal_548 ) ) ;
    buf_clk cell_205 ( .C ( clk ), .D ( signal_553 ), .Q ( signal_554 ) ) ;
    buf_clk cell_213 ( .C ( clk ), .D ( signal_561 ), .Q ( signal_562 ) ) ;
    buf_clk cell_223 ( .C ( clk ), .D ( signal_571 ), .Q ( signal_572 ) ) ;
    buf_clk cell_233 ( .C ( clk ), .D ( signal_581 ), .Q ( signal_582 ) ) ;
    buf_clk cell_243 ( .C ( clk ), .D ( signal_591 ), .Q ( signal_592 ) ) ;
    buf_clk cell_253 ( .C ( clk ), .D ( signal_601 ), .Q ( signal_602 ) ) ;
    buf_clk cell_263 ( .C ( clk ), .D ( signal_611 ), .Q ( signal_612 ) ) ;
    buf_clk cell_273 ( .C ( clk ), .D ( signal_621 ), .Q ( signal_622 ) ) ;
    buf_clk cell_283 ( .C ( clk ), .D ( signal_631 ), .Q ( signal_632 ) ) ;
    buf_clk cell_293 ( .C ( clk ), .D ( signal_641 ), .Q ( signal_642 ) ) ;
    buf_clk cell_303 ( .C ( clk ), .D ( signal_651 ), .Q ( signal_652 ) ) ;
    buf_clk cell_309 ( .C ( clk ), .D ( signal_657 ), .Q ( signal_658 ) ) ;
    buf_clk cell_315 ( .C ( clk ), .D ( signal_663 ), .Q ( signal_664 ) ) ;
    buf_clk cell_321 ( .C ( clk ), .D ( signal_669 ), .Q ( signal_670 ) ) ;
    buf_clk cell_327 ( .C ( clk ), .D ( signal_675 ), .Q ( signal_676 ) ) ;
    buf_clk cell_333 ( .C ( clk ), .D ( signal_681 ), .Q ( signal_682 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_182 ( .C ( clk ), .D ( signal_530 ), .Q ( signal_531 ) ) ;
    buf_clk cell_188 ( .C ( clk ), .D ( signal_536 ), .Q ( signal_537 ) ) ;
    buf_clk cell_194 ( .C ( clk ), .D ( signal_542 ), .Q ( signal_543 ) ) ;
    buf_clk cell_200 ( .C ( clk ), .D ( signal_548 ), .Q ( signal_549 ) ) ;
    buf_clk cell_206 ( .C ( clk ), .D ( signal_554 ), .Q ( signal_555 ) ) ;
    buf_clk cell_214 ( .C ( clk ), .D ( signal_562 ), .Q ( signal_563 ) ) ;
    buf_clk cell_224 ( .C ( clk ), .D ( signal_572 ), .Q ( signal_573 ) ) ;
    buf_clk cell_234 ( .C ( clk ), .D ( signal_582 ), .Q ( signal_583 ) ) ;
    buf_clk cell_244 ( .C ( clk ), .D ( signal_592 ), .Q ( signal_593 ) ) ;
    buf_clk cell_254 ( .C ( clk ), .D ( signal_602 ), .Q ( signal_603 ) ) ;
    buf_clk cell_264 ( .C ( clk ), .D ( signal_612 ), .Q ( signal_613 ) ) ;
    buf_clk cell_274 ( .C ( clk ), .D ( signal_622 ), .Q ( signal_623 ) ) ;
    buf_clk cell_284 ( .C ( clk ), .D ( signal_632 ), .Q ( signal_633 ) ) ;
    buf_clk cell_294 ( .C ( clk ), .D ( signal_642 ), .Q ( signal_643 ) ) ;
    buf_clk cell_304 ( .C ( clk ), .D ( signal_652 ), .Q ( signal_653 ) ) ;
    buf_clk cell_310 ( .C ( clk ), .D ( signal_658 ), .Q ( signal_659 ) ) ;
    buf_clk cell_316 ( .C ( clk ), .D ( signal_664 ), .Q ( signal_665 ) ) ;
    buf_clk cell_322 ( .C ( clk ), .D ( signal_670 ), .Q ( signal_671 ) ) ;
    buf_clk cell_328 ( .C ( clk ), .D ( signal_676 ), .Q ( signal_677 ) ) ;
    buf_clk cell_334 ( .C ( clk ), .D ( signal_682 ), .Q ( signal_683 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_54 ( .a ({signal_526, signal_524, signal_522, signal_520, signal_518}), .b ({signal_204, signal_203, signal_202, signal_201, signal_61}), .clk ( clk ), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_208, signal_207, signal_206, signal_205, signal_62}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_55 ( .a ({signal_208, signal_207, signal_206, signal_205, signal_62}), .b ({signal_212, signal_211, signal_210, signal_209, signal_63}) ) ;
    buf_clk cell_183 ( .C ( clk ), .D ( signal_531 ), .Q ( signal_532 ) ) ;
    buf_clk cell_189 ( .C ( clk ), .D ( signal_537 ), .Q ( signal_538 ) ) ;
    buf_clk cell_195 ( .C ( clk ), .D ( signal_543 ), .Q ( signal_544 ) ) ;
    buf_clk cell_201 ( .C ( clk ), .D ( signal_549 ), .Q ( signal_550 ) ) ;
    buf_clk cell_207 ( .C ( clk ), .D ( signal_555 ), .Q ( signal_556 ) ) ;
    buf_clk cell_215 ( .C ( clk ), .D ( signal_563 ), .Q ( signal_564 ) ) ;
    buf_clk cell_225 ( .C ( clk ), .D ( signal_573 ), .Q ( signal_574 ) ) ;
    buf_clk cell_235 ( .C ( clk ), .D ( signal_583 ), .Q ( signal_584 ) ) ;
    buf_clk cell_245 ( .C ( clk ), .D ( signal_593 ), .Q ( signal_594 ) ) ;
    buf_clk cell_255 ( .C ( clk ), .D ( signal_603 ), .Q ( signal_604 ) ) ;
    buf_clk cell_265 ( .C ( clk ), .D ( signal_613 ), .Q ( signal_614 ) ) ;
    buf_clk cell_275 ( .C ( clk ), .D ( signal_623 ), .Q ( signal_624 ) ) ;
    buf_clk cell_285 ( .C ( clk ), .D ( signal_633 ), .Q ( signal_634 ) ) ;
    buf_clk cell_295 ( .C ( clk ), .D ( signal_643 ), .Q ( signal_644 ) ) ;
    buf_clk cell_305 ( .C ( clk ), .D ( signal_653 ), .Q ( signal_654 ) ) ;
    buf_clk cell_311 ( .C ( clk ), .D ( signal_659 ), .Q ( signal_660 ) ) ;
    buf_clk cell_317 ( .C ( clk ), .D ( signal_665 ), .Q ( signal_666 ) ) ;
    buf_clk cell_323 ( .C ( clk ), .D ( signal_671 ), .Q ( signal_672 ) ) ;
    buf_clk cell_329 ( .C ( clk ), .D ( signal_677 ), .Q ( signal_678 ) ) ;
    buf_clk cell_335 ( .C ( clk ), .D ( signal_683 ), .Q ( signal_684 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_216 ( .C ( clk ), .D ( signal_564 ), .Q ( signal_565 ) ) ;
    buf_clk cell_226 ( .C ( clk ), .D ( signal_574 ), .Q ( signal_575 ) ) ;
    buf_clk cell_236 ( .C ( clk ), .D ( signal_584 ), .Q ( signal_585 ) ) ;
    buf_clk cell_246 ( .C ( clk ), .D ( signal_594 ), .Q ( signal_595 ) ) ;
    buf_clk cell_256 ( .C ( clk ), .D ( signal_604 ), .Q ( signal_605 ) ) ;
    buf_clk cell_266 ( .C ( clk ), .D ( signal_614 ), .Q ( signal_615 ) ) ;
    buf_clk cell_276 ( .C ( clk ), .D ( signal_624 ), .Q ( signal_625 ) ) ;
    buf_clk cell_286 ( .C ( clk ), .D ( signal_634 ), .Q ( signal_635 ) ) ;
    buf_clk cell_296 ( .C ( clk ), .D ( signal_644 ), .Q ( signal_645 ) ) ;
    buf_clk cell_306 ( .C ( clk ), .D ( signal_654 ), .Q ( signal_655 ) ) ;
    buf_clk cell_312 ( .C ( clk ), .D ( signal_660 ), .Q ( signal_661 ) ) ;
    buf_clk cell_318 ( .C ( clk ), .D ( signal_666 ), .Q ( signal_667 ) ) ;
    buf_clk cell_324 ( .C ( clk ), .D ( signal_672 ), .Q ( signal_673 ) ) ;
    buf_clk cell_330 ( .C ( clk ), .D ( signal_678 ), .Q ( signal_679 ) ) ;
    buf_clk cell_336 ( .C ( clk ), .D ( signal_684 ), .Q ( signal_685 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(4), .pipeline(1)) cell_56 ( .a ({signal_556, signal_550, signal_544, signal_538, signal_532}), .b ({signal_212, signal_211, signal_210, signal_209, signal_63}), .clk ( clk ), .r ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .c ({signal_216, signal_215, signal_214, signal_213, signal_64}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) cell_57 ( .a ({signal_216, signal_215, signal_214, signal_213, signal_64}), .b ({signal_220, signal_219, signal_218, signal_217, signal_18}) ) ;
    buf_clk cell_217 ( .C ( clk ), .D ( signal_565 ), .Q ( signal_566 ) ) ;
    buf_clk cell_227 ( .C ( clk ), .D ( signal_575 ), .Q ( signal_576 ) ) ;
    buf_clk cell_237 ( .C ( clk ), .D ( signal_585 ), .Q ( signal_586 ) ) ;
    buf_clk cell_247 ( .C ( clk ), .D ( signal_595 ), .Q ( signal_596 ) ) ;
    buf_clk cell_257 ( .C ( clk ), .D ( signal_605 ), .Q ( signal_606 ) ) ;
    buf_clk cell_267 ( .C ( clk ), .D ( signal_615 ), .Q ( signal_616 ) ) ;
    buf_clk cell_277 ( .C ( clk ), .D ( signal_625 ), .Q ( signal_626 ) ) ;
    buf_clk cell_287 ( .C ( clk ), .D ( signal_635 ), .Q ( signal_636 ) ) ;
    buf_clk cell_297 ( .C ( clk ), .D ( signal_645 ), .Q ( signal_646 ) ) ;
    buf_clk cell_307 ( .C ( clk ), .D ( signal_655 ), .Q ( signal_656 ) ) ;
    buf_clk cell_313 ( .C ( clk ), .D ( signal_661 ), .Q ( signal_662 ) ) ;
    buf_clk cell_319 ( .C ( clk ), .D ( signal_667 ), .Q ( signal_668 ) ) ;
    buf_clk cell_325 ( .C ( clk ), .D ( signal_673 ), .Q ( signal_674 ) ) ;
    buf_clk cell_331 ( .C ( clk ), .D ( signal_679 ), .Q ( signal_680 ) ) ;
    buf_clk cell_337 ( .C ( clk ), .D ( signal_685 ), .Q ( signal_686 ) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_606, signal_596, signal_586, signal_576, signal_566}), .Q ({SO_s4[3], SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_656, signal_646, signal_636, signal_626, signal_616}), .Q ({SO_s4[2], SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_686, signal_680, signal_674, signal_668, signal_662}), .Q ({SO_s4[1], SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_220, signal_219, signal_218, signal_217, signal_18}), .Q ({SO_s4[0], SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
