/* modified netlist. Source: module CRAFT in file ../CaseStudies/09_CRAFT_round_based_encryption/FPGA_based/CRAFT_synthesis.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module CRAFT_GHPC_ClockGating_d1 (clk, rst, Input_s0, Key_s0, Key_s1, Input_s1, Fresh, done, Output_s0, Output_s1, Synch);
    input clk ;
    input rst ;
    input [63:0] Input_s0 ;
    input [127:0] Key_s0 ;
    input [127:0] Key_s1 ;
    input [63:0] Input_s1 ;
    input [63:0] Fresh ;
    output done ;
    output [63:0] Output_s0 ;
    output [63:0] Output_s1 ;
    output Synch ;
    wire [6:1] \FSM ;
    wire [6:2] \FSMUpdate ;
    wire done_internal ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N10 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N30 ;
    wire N32 ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N50 ;
    wire N52 ;
    wire N54 ;
    wire N55 ;
    wire N57 ;
    wire N58 ;
    wire N60 ;
    wire N61 ;
    wire N63 ;
    wire N64 ;
    wire N66 ;
    wire N67 ;
    wire N69 ;
    wire N70 ;
    wire N72 ;
    wire N73 ;
    wire N75 ;
    wire N77 ;
    wire N79 ;
    wire N81 ;
    wire N83 ;
    wire N85 ;
    wire N87 ;
    wire N89 ;
    wire N91 ;
    wire N93 ;
    wire N95 ;
    wire N97 ;
    wire N99 ;
    wire N101 ;
    wire N103 ;
    wire N105 ;
    wire N107 ;
    wire [6:0] \FSMRegInst/s_current_state ;
    wire [0:0] \selectsRegInst/s_current_state ;
    wire [0:0] selectsNext ;
    wire [63:0] Feedback ;
    wire [63:0] AddRoundKeyOutput ;
    wire new_AGEMA_signal_731 ;
    wire new_AGEMA_signal_732 ;
    wire new_AGEMA_signal_733 ;
    wire new_AGEMA_signal_734 ;
    wire new_AGEMA_signal_739 ;
    wire new_AGEMA_signal_740 ;
    wire new_AGEMA_signal_741 ;
    wire new_AGEMA_signal_742 ;
    wire new_AGEMA_signal_747 ;
    wire new_AGEMA_signal_748 ;
    wire new_AGEMA_signal_749 ;
    wire new_AGEMA_signal_750 ;
    wire new_AGEMA_signal_755 ;
    wire new_AGEMA_signal_756 ;
    wire new_AGEMA_signal_757 ;
    wire new_AGEMA_signal_758 ;
    wire new_AGEMA_signal_763 ;
    wire new_AGEMA_signal_764 ;
    wire new_AGEMA_signal_765 ;
    wire new_AGEMA_signal_766 ;
    wire new_AGEMA_signal_771 ;
    wire new_AGEMA_signal_772 ;
    wire new_AGEMA_signal_773 ;
    wire new_AGEMA_signal_774 ;
    wire new_AGEMA_signal_779 ;
    wire new_AGEMA_signal_780 ;
    wire new_AGEMA_signal_781 ;
    wire new_AGEMA_signal_782 ;
    wire new_AGEMA_signal_787 ;
    wire new_AGEMA_signal_788 ;
    wire new_AGEMA_signal_789 ;
    wire new_AGEMA_signal_790 ;
    wire new_AGEMA_signal_795 ;
    wire new_AGEMA_signal_796 ;
    wire new_AGEMA_signal_797 ;
    wire new_AGEMA_signal_798 ;
    wire new_AGEMA_signal_803 ;
    wire new_AGEMA_signal_804 ;
    wire new_AGEMA_signal_805 ;
    wire new_AGEMA_signal_806 ;
    wire new_AGEMA_signal_811 ;
    wire new_AGEMA_signal_812 ;
    wire new_AGEMA_signal_813 ;
    wire new_AGEMA_signal_814 ;
    wire new_AGEMA_signal_819 ;
    wire new_AGEMA_signal_820 ;
    wire new_AGEMA_signal_821 ;
    wire new_AGEMA_signal_822 ;
    wire new_AGEMA_signal_827 ;
    wire new_AGEMA_signal_828 ;
    wire new_AGEMA_signal_829 ;
    wire new_AGEMA_signal_830 ;
    wire new_AGEMA_signal_835 ;
    wire new_AGEMA_signal_836 ;
    wire new_AGEMA_signal_837 ;
    wire new_AGEMA_signal_838 ;
    wire new_AGEMA_signal_843 ;
    wire new_AGEMA_signal_844 ;
    wire new_AGEMA_signal_845 ;
    wire new_AGEMA_signal_846 ;
    wire new_AGEMA_signal_851 ;
    wire new_AGEMA_signal_852 ;
    wire new_AGEMA_signal_853 ;
    wire new_AGEMA_signal_854 ;
    wire new_AGEMA_signal_857 ;
    wire new_AGEMA_signal_860 ;
    wire new_AGEMA_signal_863 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_872 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_878 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_887 ;
    wire new_AGEMA_signal_890 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_896 ;
    wire new_AGEMA_signal_899 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_908 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[1].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [1]), .O (\FSM [1]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[2].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [2]), .O (\FSM [2]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[4].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [4]), .O (\FSM [4]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[5].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [5]), .O (\FSM [5]) ) ;
    LUT2 #( .INIT ( 4'h4 ) ) \FSMMUX/GEN[6].MUXInst/Mmux_Q11 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [6]), .O (\FSM [6]) ) ;
    LUT3 #( .INIT ( 8'h54 ) ) \FSMSignalsInst/done<6>_SW0 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [5]), .I2 (\FSMRegInst/s_current_state [4]), .O (N2) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[0].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[32], Key_s0[32]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[96], Key_s0[96]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_857, N4}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[1].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[33], Key_s0[33]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[97], Key_s0[97]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_860, N6}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[2].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[34], Key_s0[34]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[98], Key_s0[98]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_863, N8}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[3].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[35], Key_s0[35]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[99], Key_s0[99]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_866, N10}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[4].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[36], Key_s0[36]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[100], Key_s0[100]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_869, N12}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[5].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[37], Key_s0[37]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[101], Key_s0[101]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_872, N14}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[6].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[38], Key_s0[38]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[102], Key_s0[102]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_875, N16}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[7].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[39], Key_s0[39]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[103], Key_s0[103]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_878, N18}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[11].XOR_r1_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[43], Key_s0[43]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[107], Key_s0[107]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_881, N20}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[0].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[48], Key_s0[48]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[112], Key_s0[112]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_884, N22}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[1].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[49], Key_s0[49]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[113], Key_s0[113]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_887, N24}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[2].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[50], Key_s0[50]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[114], Key_s0[114]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_890, N26}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[3].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[51], Key_s0[51]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[115], Key_s0[115]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_893, N28}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[4].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[52], Key_s0[52]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[116], Key_s0[116]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_896, N30}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[5].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[53], Key_s0[53]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[117], Key_s0[117]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_899, N32}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[6].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[54], Key_s0[54]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[118], Key_s0[118]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_902, N34}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[7].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[55], Key_s0[55]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[119], Key_s0[119]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_905, N36}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[8].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[56], Key_s0[56]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[120], Key_s0[120]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_908, N38}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[9].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[57], Key_s0[57]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[121], Key_s0[121]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_911, N40}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[10].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[58], Key_s0[58]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[122], Key_s0[122]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_914, N42}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[11].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[59], Key_s0[59]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[123], Key_s0[123]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_917, N44}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[12].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[60], Key_s0[60]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[124], Key_s0[124]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_920, N46}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[13].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[61], Key_s0[61]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[125], Key_s0[125]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_923, N48}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[14].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[62], Key_s0[62]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[126], Key_s0[126]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_926, N50}) ) ;
    LUT4_masked #(.low_latency(0), .pipeline(0),  .INIT ( 16'h1D0F ) , .MASK ( 4'b1010 ), .INIT2 ( 16'hE2F0 ) ) \MCInst/GEN[15].XOR_r0_Inst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[63], Key_s0[63]}), .I1 ({1'b0, rst}), .I2 ({Key_s1[127], Key_s0[127]}), .I3 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_929, N52}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[46], Key_s0[46]}), .I1 ({Key_s1[110], Key_s0[110]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_932, N54}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[110], Key_s0[110]}), .I1 ({Input_s1[46], Input_s0[46]}), .I2 ({Input_s1[14], Input_s0[14]}), .O ({new_AGEMA_signal_935, N55}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[45], Key_s0[45]}), .I1 ({Key_s1[109], Key_s0[109]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_938, N57}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[109], Key_s0[109]}), .I1 ({Input_s1[45], Input_s0[45]}), .I2 ({Input_s1[13], Input_s0[13]}), .O ({new_AGEMA_signal_941, N58}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[47], Key_s0[47]}), .I1 ({Key_s1[111], Key_s0[111]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_944, N60}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[111], Key_s0[111]}), .I1 ({Input_s1[47], Input_s0[47]}), .I2 ({Input_s1[15], Input_s0[15]}), .O ({new_AGEMA_signal_947, N61}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[44], Key_s0[44]}), .I1 ({Key_s1[108], Key_s0[108]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_950, N63}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[108], Key_s0[108]}), .I1 ({Input_s1[44], Input_s0[44]}), .I2 ({Input_s1[12], Input_s0[12]}), .O ({new_AGEMA_signal_953, N64}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[42], Key_s0[42]}), .I1 ({Key_s1[106], Key_s0[106]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_956, N66}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[106], Key_s0[106]}), .I1 ({Input_s1[42], Input_s0[42]}), .I2 ({Input_s1[10], Input_s0[10]}), .O ({new_AGEMA_signal_959, N67}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[41], Key_s0[41]}), .I1 ({Key_s1[105], Key_s0[105]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_962, N69}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[105], Key_s0[105]}), .I1 ({Input_s1[9], Input_s0[9]}), .I2 ({Input_s1[41], Input_s0[41]}), .O ({new_AGEMA_signal_965, N70}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'hAC ) , .MASK ( 3'b100 ), .INIT2 ( 8'hAC ) ) \AddKeyConstXOR/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Key_s1[40], Key_s0[40]}), .I1 ({Key_s1[104], Key_s0[104]}), .I2 ({1'b0, \selectsRegInst/s_current_state [0]}), .O ({new_AGEMA_signal_968, N72}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyConstXOR/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW1 ( .I0 ({Key_s1[104], Key_s0[104]}), .I1 ({Input_s1[8], Input_s0[8]}), .I2 ({Input_s1[40], Input_s0[40]}), .O ({new_AGEMA_signal_971, N73}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[48], Input_s0[48]}), .I1 ({Input_s1[16], Input_s0[16]}), .I2 ({Input_s1[0], Input_s0[0]}), .O ({new_AGEMA_signal_975, N75}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[49], Input_s0[49]}), .I1 ({Input_s1[1], Input_s0[1]}), .I2 ({Input_s1[17], Input_s0[17]}), .O ({new_AGEMA_signal_979, N77}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[50], Input_s0[50]}), .I1 ({Input_s1[2], Input_s0[2]}), .I2 ({Input_s1[18], Input_s0[18]}), .O ({new_AGEMA_signal_983, N79}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[51], Input_s0[51]}), .I1 ({Input_s1[3], Input_s0[3]}), .I2 ({Input_s1[19], Input_s0[19]}), .O ({new_AGEMA_signal_987, N81}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[52], Input_s0[52]}), .I1 ({Input_s1[4], Input_s0[4]}), .I2 ({Input_s1[20], Input_s0[20]}), .O ({new_AGEMA_signal_991, N83}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[5], Input_s0[5]}), .I1 ({Input_s1[53], Input_s0[53]}), .I2 ({Input_s1[21], Input_s0[21]}), .O ({new_AGEMA_signal_995, N85}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[6], Input_s0[6]}), .I1 ({Input_s1[54], Input_s0[54]}), .I2 ({Input_s1[22], Input_s0[22]}), .O ({new_AGEMA_signal_999, N87}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[7], Input_s0[7]}), .I1 ({Input_s1[55], Input_s0[55]}), .I2 ({Input_s1[23], Input_s0[23]}), .O ({new_AGEMA_signal_1003, N89}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[8], Input_s0[8]}), .I1 ({Input_s1[56], Input_s0[56]}), .I2 ({Input_s1[24], Input_s0[24]}), .O ({new_AGEMA_signal_1006, N91}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[9], Input_s0[9]}), .I1 ({Input_s1[57], Input_s0[57]}), .I2 ({Input_s1[25], Input_s0[25]}), .O ({new_AGEMA_signal_1009, N93}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[58], Input_s0[58]}), .I1 ({Input_s1[26], Input_s0[26]}), .I2 ({Input_s1[10], Input_s0[10]}), .O ({new_AGEMA_signal_1012, N95}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[2].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[59], Input_s0[59]}), .I1 ({Input_s1[27], Input_s0[27]}), .I2 ({Input_s1[11], Input_s0[11]}), .O ({new_AGEMA_signal_1016, N97}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[0].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[60], Input_s0[60]}), .I1 ({Input_s1[28], Input_s0[28]}), .I2 ({Input_s1[12], Input_s0[12]}), .O ({new_AGEMA_signal_1019, N99}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[1].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[61], Input_s0[61]}), .I1 ({Input_s1[29], Input_s0[29]}), .I2 ({Input_s1[13], Input_s0[13]}), .O ({new_AGEMA_signal_1022, N101}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[2].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[62], Input_s0[62]}), .I1 ({Input_s1[30], Input_s0[30]}), .I2 ({Input_s1[14], Input_s0[14]}), .O ({new_AGEMA_signal_1025, N103}) ) ;
    LUT3_masked #(.low_latency(0), .pipeline(0),  .INIT ( 8'h96 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \AddKeyXOR1/GEN1[3].GEN2[3].XORInst/Mxor_Q_xo<0>1_SW0 ( .I0 ({Input_s1[63], Input_s0[63]}), .I1 ({Input_s1[31], Input_s0[31]}), .I2 ({Input_s1[15], Input_s0[15]}), .O ({new_AGEMA_signal_1028, N105}) ) ;
    LUT2 #( .INIT ( 4'hD ) ) \selectsUpdateInst/selectsNext<0>1 ( .I0 (\selectsRegInst/s_current_state [0]), .I1 (rst), .O (selectsNext[0]) ) ;
    LUT3 #( .INIT ( 8'hBE ) ) \FSMUpdateInst/Mxor_FSMUpdate<2>_xo<0>1 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [1]), .I2 (\FSMRegInst/s_current_state [0]), .O (\FSMUpdate [2]) ) ;
    LUT3 #( .INIT ( 8'hBE ) ) \FSMUpdateInst/Mxor_FSMUpdate<6>_xo<0>1 ( .I0 (rst), .I1 (\FSMRegInst/s_current_state [4]), .I2 (\FSMRegInst/s_current_state [3]), .O (\FSMUpdate [6]) ) ;
    MUXF7 \FSMSignalsInst/done<6> ( .S (N2), .I0 (N107), .I1 (1'b0), .O (done_internal) ) ;
    LUT6 #( .INIT ( 64'h0000000000000080 ) ) \FSMSignalsInst/done<6>_F ( .I0 (\FSMRegInst/s_current_state [0]), .I1 (\FSMRegInst/s_current_state [6]), .I2 (\FSMRegInst/s_current_state [2]), .I3 (rst), .I4 (\FSMRegInst/s_current_state [1]), .I5 (\FSMRegInst/s_current_state [3]), .O (N107) ) ;
    ClockGatingController #(3) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[0].SboxInst/y_0 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r (Fresh[0]), .O ({new_AGEMA_signal_731, Feedback[0]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[0].SboxInst/y_1 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r (Fresh[1]), .O ({new_AGEMA_signal_732, Feedback[1]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[0].SboxInst/y_2 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r (Fresh[2]), .O ({new_AGEMA_signal_733, Feedback[2]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[0].SboxInst/y_3 ( .I0 ({Output_s1[60], Output_s0[60]}), .I1 ({Output_s1[61], Output_s0[61]}), .I2 ({Output_s1[62], Output_s0[62]}), .I3 ({Output_s1[63], Output_s0[63]}), .clk (clk), .r (Fresh[3]), .O ({new_AGEMA_signal_734, Feedback[3]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[1].SboxInst/y_0 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r (Fresh[4]), .O ({new_AGEMA_signal_739, Feedback[4]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[1].SboxInst/y_1 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r (Fresh[5]), .O ({new_AGEMA_signal_740, Feedback[5]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[1].SboxInst/y_2 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r (Fresh[6]), .O ({new_AGEMA_signal_741, Feedback[6]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[1].SboxInst/y_3 ( .I0 ({Output_s1[48], Output_s0[48]}), .I1 ({Output_s1[49], Output_s0[49]}), .I2 ({Output_s1[50], Output_s0[50]}), .I3 ({Output_s1[51], Output_s0[51]}), .clk (clk), .r (Fresh[7]), .O ({new_AGEMA_signal_742, Feedback[7]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[2].SboxInst/y_0 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r (Fresh[8]), .O ({new_AGEMA_signal_747, Feedback[8]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[2].SboxInst/y_1 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r (Fresh[9]), .O ({new_AGEMA_signal_748, Feedback[9]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[2].SboxInst/y_2 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r (Fresh[10]), .O ({new_AGEMA_signal_749, Feedback[10]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[2].SboxInst/y_3 ( .I0 ({Output_s1[52], Output_s0[52]}), .I1 ({Output_s1[53], Output_s0[53]}), .I2 ({Output_s1[54], Output_s0[54]}), .I3 ({Output_s1[55], Output_s0[55]}), .clk (clk), .r (Fresh[11]), .O ({new_AGEMA_signal_750, Feedback[11]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[3].SboxInst/y_0 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r (Fresh[12]), .O ({new_AGEMA_signal_755, Feedback[12]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[3].SboxInst/y_1 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r (Fresh[13]), .O ({new_AGEMA_signal_756, Feedback[13]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[3].SboxInst/y_2 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r (Fresh[14]), .O ({new_AGEMA_signal_757, Feedback[14]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[3].SboxInst/y_3 ( .I0 ({Output_s1[56], Output_s0[56]}), .I1 ({Output_s1[57], Output_s0[57]}), .I2 ({Output_s1[58], Output_s0[58]}), .I3 ({Output_s1[59], Output_s0[59]}), .clk (clk), .r (Fresh[15]), .O ({new_AGEMA_signal_758, Feedback[15]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[4].SboxInst/y_0 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r (Fresh[16]), .O ({new_AGEMA_signal_763, Feedback[16]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[4].SboxInst/y_1 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r (Fresh[17]), .O ({new_AGEMA_signal_764, Feedback[17]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[4].SboxInst/y_2 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r (Fresh[18]), .O ({new_AGEMA_signal_765, Feedback[18]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[4].SboxInst/y_3 ( .I0 ({Output_s1[32], Output_s0[32]}), .I1 ({Output_s1[33], Output_s0[33]}), .I2 ({Output_s1[34], Output_s0[34]}), .I3 ({Output_s1[35], Output_s0[35]}), .clk (clk), .r (Fresh[19]), .O ({new_AGEMA_signal_766, Feedback[19]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[5].SboxInst/y_0 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r (Fresh[20]), .O ({new_AGEMA_signal_771, Feedback[20]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[5].SboxInst/y_1 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r (Fresh[21]), .O ({new_AGEMA_signal_772, Feedback[21]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[5].SboxInst/y_2 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r (Fresh[22]), .O ({new_AGEMA_signal_773, Feedback[22]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[5].SboxInst/y_3 ( .I0 ({Output_s1[44], Output_s0[44]}), .I1 ({Output_s1[45], Output_s0[45]}), .I2 ({Output_s1[46], Output_s0[46]}), .I3 ({Output_s1[47], Output_s0[47]}), .clk (clk), .r (Fresh[23]), .O ({new_AGEMA_signal_774, Feedback[23]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[6].SboxInst/y_0 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r (Fresh[24]), .O ({new_AGEMA_signal_779, Feedback[24]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[6].SboxInst/y_1 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r (Fresh[25]), .O ({new_AGEMA_signal_780, Feedback[25]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[6].SboxInst/y_2 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r (Fresh[26]), .O ({new_AGEMA_signal_781, Feedback[26]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[6].SboxInst/y_3 ( .I0 ({Output_s1[40], Output_s0[40]}), .I1 ({Output_s1[41], Output_s0[41]}), .I2 ({Output_s1[42], Output_s0[42]}), .I3 ({Output_s1[43], Output_s0[43]}), .clk (clk), .r (Fresh[27]), .O ({new_AGEMA_signal_782, Feedback[27]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[7].SboxInst/y_0 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r (Fresh[28]), .O ({new_AGEMA_signal_787, Feedback[28]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[7].SboxInst/y_1 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r (Fresh[29]), .O ({new_AGEMA_signal_788, Feedback[29]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[7].SboxInst/y_2 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r (Fresh[30]), .O ({new_AGEMA_signal_789, Feedback[30]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[7].SboxInst/y_3 ( .I0 ({Output_s1[36], Output_s0[36]}), .I1 ({Output_s1[37], Output_s0[37]}), .I2 ({Output_s1[38], Output_s0[38]}), .I3 ({Output_s1[39], Output_s0[39]}), .clk (clk), .r (Fresh[31]), .O ({new_AGEMA_signal_790, Feedback[31]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[8].SboxInst/y_0 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r (Fresh[32]), .O ({new_AGEMA_signal_795, Feedback[32]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[8].SboxInst/y_1 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r (Fresh[33]), .O ({new_AGEMA_signal_796, Feedback[33]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[8].SboxInst/y_2 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r (Fresh[34]), .O ({new_AGEMA_signal_797, Feedback[34]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[8].SboxInst/y_3 ( .I0 ({Output_s1[16], Output_s0[16]}), .I1 ({Output_s1[17], Output_s0[17]}), .I2 ({Output_s1[18], Output_s0[18]}), .I3 ({Output_s1[19], Output_s0[19]}), .clk (clk), .r (Fresh[35]), .O ({new_AGEMA_signal_798, Feedback[35]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[9].SboxInst/y_0 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r (Fresh[36]), .O ({new_AGEMA_signal_803, Feedback[36]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[9].SboxInst/y_1 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r (Fresh[37]), .O ({new_AGEMA_signal_804, Feedback[37]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[9].SboxInst/y_2 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r (Fresh[38]), .O ({new_AGEMA_signal_805, Feedback[38]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[9].SboxInst/y_3 ( .I0 ({Output_s1[28], Output_s0[28]}), .I1 ({Output_s1[29], Output_s0[29]}), .I2 ({Output_s1[30], Output_s0[30]}), .I3 ({Output_s1[31], Output_s0[31]}), .clk (clk), .r (Fresh[39]), .O ({new_AGEMA_signal_806, Feedback[39]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[10].SboxInst/y_0 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r (Fresh[40]), .O ({new_AGEMA_signal_811, Feedback[40]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[10].SboxInst/y_1 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r (Fresh[41]), .O ({new_AGEMA_signal_812, Feedback[41]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[10].SboxInst/y_2 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r (Fresh[42]), .O ({new_AGEMA_signal_813, Feedback[42]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[10].SboxInst/y_3 ( .I0 ({Output_s1[24], Output_s0[24]}), .I1 ({Output_s1[25], Output_s0[25]}), .I2 ({Output_s1[26], Output_s0[26]}), .I3 ({Output_s1[27], Output_s0[27]}), .clk (clk), .r (Fresh[43]), .O ({new_AGEMA_signal_814, Feedback[43]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[11].SboxInst/y_0 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r (Fresh[44]), .O ({new_AGEMA_signal_819, Feedback[44]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[11].SboxInst/y_1 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r (Fresh[45]), .O ({new_AGEMA_signal_820, Feedback[45]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[11].SboxInst/y_2 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r (Fresh[46]), .O ({new_AGEMA_signal_821, Feedback[46]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[11].SboxInst/y_3 ( .I0 ({Output_s1[20], Output_s0[20]}), .I1 ({Output_s1[21], Output_s0[21]}), .I2 ({Output_s1[22], Output_s0[22]}), .I3 ({Output_s1[23], Output_s0[23]}), .clk (clk), .r (Fresh[47]), .O ({new_AGEMA_signal_822, Feedback[47]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[12].SboxInst/y_0 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r (Fresh[48]), .O ({new_AGEMA_signal_827, Feedback[48]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[12].SboxInst/y_1 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r (Fresh[49]), .O ({new_AGEMA_signal_828, Feedback[49]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[12].SboxInst/y_2 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r (Fresh[50]), .O ({new_AGEMA_signal_829, Feedback[50]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[12].SboxInst/y_3 ( .I0 ({Output_s1[4], Output_s0[4]}), .I1 ({Output_s1[5], Output_s0[5]}), .I2 ({Output_s1[6], Output_s0[6]}), .I3 ({Output_s1[7], Output_s0[7]}), .clk (clk), .r (Fresh[51]), .O ({new_AGEMA_signal_830, Feedback[51]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[13].SboxInst/y_0 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r (Fresh[52]), .O ({new_AGEMA_signal_835, Feedback[52]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[13].SboxInst/y_1 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r (Fresh[53]), .O ({new_AGEMA_signal_836, Feedback[53]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[13].SboxInst/y_2 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r (Fresh[54]), .O ({new_AGEMA_signal_837, Feedback[54]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[13].SboxInst/y_3 ( .I0 ({Output_s1[8], Output_s0[8]}), .I1 ({Output_s1[9], Output_s0[9]}), .I2 ({Output_s1[10], Output_s0[10]}), .I3 ({Output_s1[11], Output_s0[11]}), .clk (clk), .r (Fresh[55]), .O ({new_AGEMA_signal_838, Feedback[55]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[14].SboxInst/y_0 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r (Fresh[56]), .O ({new_AGEMA_signal_843, Feedback[56]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[14].SboxInst/y_1 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r (Fresh[57]), .O ({new_AGEMA_signal_844, Feedback[57]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[14].SboxInst/y_2 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r (Fresh[58]), .O ({new_AGEMA_signal_845, Feedback[58]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[14].SboxInst/y_3 ( .I0 ({Output_s1[12], Output_s0[12]}), .I1 ({Output_s1[13], Output_s0[13]}), .I2 ({Output_s1[14], Output_s0[14]}), .I3 ({Output_s1[15], Output_s0[15]}), .clk (clk), .r (Fresh[59]), .O ({new_AGEMA_signal_846, Feedback[59]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0EEC ) ) \SubCellInst/GEN[15].SboxInst/y_0 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r (Fresh[60]), .O ({new_AGEMA_signal_851, Feedback[60]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hA0FA ) ) \SubCellInst/GEN[15].SboxInst/y_1 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r (Fresh[61]), .O ({new_AGEMA_signal_852, Feedback[61]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'hC8D5 ) ) \SubCellInst/GEN[15].SboxInst/y_2 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r (Fresh[62]), .O ({new_AGEMA_signal_853, Feedback[62]}) ) ;
    LUT4_GHPC #(.low_latency(0), .pipeline(0),  .INIT ( 16'h0377 ) ) \SubCellInst/GEN[15].SboxInst/y_3 ( .I0 ({Output_s1[0], Output_s0[0]}), .I1 ({Output_s1[1], Output_s0[1]}), .I2 ({Output_s1[2], Output_s0[2]}), .I3 ({Output_s1[3], Output_s0[3]}), .clk (clk), .r (Fresh[63]), .O ({new_AGEMA_signal_854, Feedback[63]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[0], Input_s0[0]}), .I1 ({Key_s1[0], Key_s0[0]}), .I2 ({Key_s1[64], Key_s0[64]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_731, Feedback[0]}), .O ({new_AGEMA_signal_1031, AddRoundKeyOutput[0]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[10], Input_s0[10]}), .I1 ({Key_s1[10], Key_s0[10]}), .I2 ({Key_s1[74], Key_s0[74]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_749, Feedback[10]}), .O ({new_AGEMA_signal_1034, AddRoundKeyOutput[10]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[11], Input_s0[11]}), .I1 ({Key_s1[11], Key_s0[11]}), .I2 ({Key_s1[75], Key_s0[75]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_750, Feedback[11]}), .O ({new_AGEMA_signal_1037, AddRoundKeyOutput[11]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[12], Input_s0[12]}), .I1 ({Key_s1[12], Key_s0[12]}), .I2 ({Key_s1[76], Key_s0[76]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_755, Feedback[12]}), .O ({new_AGEMA_signal_1040, AddRoundKeyOutput[12]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[13], Input_s0[13]}), .I1 ({Key_s1[13], Key_s0[13]}), .I2 ({Key_s1[77], Key_s0[77]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_756, Feedback[13]}), .O ({new_AGEMA_signal_1043, AddRoundKeyOutput[13]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[14], Input_s0[14]}), .I1 ({Key_s1[14], Key_s0[14]}), .I2 ({Key_s1[78], Key_s0[78]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_757, Feedback[14]}), .O ({new_AGEMA_signal_1046, AddRoundKeyOutput[14]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[3].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[15], Input_s0[15]}), .I1 ({Key_s1[15], Key_s0[15]}), .I2 ({Key_s1[79], Key_s0[79]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_758, Feedback[15]}), .O ({new_AGEMA_signal_1049, AddRoundKeyOutput[15]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[16], Input_s0[16]}), .I1 ({Key_s1[16], Key_s0[16]}), .I2 ({Key_s1[80], Key_s0[80]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_763, Feedback[16]}), .O ({new_AGEMA_signal_1052, AddRoundKeyOutput[16]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[17], Input_s0[17]}), .I1 ({Key_s1[17], Key_s0[17]}), .I2 ({Key_s1[81], Key_s0[81]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_764, Feedback[17]}), .O ({new_AGEMA_signal_1055, AddRoundKeyOutput[17]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[18], Input_s0[18]}), .I1 ({Key_s1[18], Key_s0[18]}), .I2 ({Key_s1[82], Key_s0[82]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_765, Feedback[18]}), .O ({new_AGEMA_signal_1058, AddRoundKeyOutput[18]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[4].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[19], Input_s0[19]}), .I1 ({Key_s1[19], Key_s0[19]}), .I2 ({Key_s1[83], Key_s0[83]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_766, Feedback[19]}), .O ({new_AGEMA_signal_1061, AddRoundKeyOutput[19]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[1], Input_s0[1]}), .I1 ({Key_s1[1], Key_s0[1]}), .I2 ({Key_s1[65], Key_s0[65]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_732, Feedback[1]}), .O ({new_AGEMA_signal_1064, AddRoundKeyOutput[1]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[20], Input_s0[20]}), .I1 ({Key_s1[20], Key_s0[20]}), .I2 ({Key_s1[84], Key_s0[84]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_771, Feedback[20]}), .O ({new_AGEMA_signal_1067, AddRoundKeyOutput[20]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[21], Input_s0[21]}), .I1 ({Key_s1[21], Key_s0[21]}), .I2 ({Key_s1[85], Key_s0[85]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_772, Feedback[21]}), .O ({new_AGEMA_signal_1070, AddRoundKeyOutput[21]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[22], Input_s0[22]}), .I1 ({Key_s1[22], Key_s0[22]}), .I2 ({Key_s1[86], Key_s0[86]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_773, Feedback[22]}), .O ({new_AGEMA_signal_1073, AddRoundKeyOutput[22]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[5].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[23], Input_s0[23]}), .I1 ({Key_s1[23], Key_s0[23]}), .I2 ({Key_s1[87], Key_s0[87]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_774, Feedback[23]}), .O ({new_AGEMA_signal_1076, AddRoundKeyOutput[23]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[24], Input_s0[24]}), .I1 ({Key_s1[24], Key_s0[24]}), .I2 ({Key_s1[88], Key_s0[88]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_779, Feedback[24]}), .O ({new_AGEMA_signal_1079, AddRoundKeyOutput[24]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[25], Input_s0[25]}), .I1 ({Key_s1[25], Key_s0[25]}), .I2 ({Key_s1[89], Key_s0[89]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_780, Feedback[25]}), .O ({new_AGEMA_signal_1082, AddRoundKeyOutput[25]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[26], Input_s0[26]}), .I1 ({Key_s1[26], Key_s0[26]}), .I2 ({Key_s1[90], Key_s0[90]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_781, Feedback[26]}), .O ({new_AGEMA_signal_1085, AddRoundKeyOutput[26]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[6].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[27], Input_s0[27]}), .I1 ({Key_s1[27], Key_s0[27]}), .I2 ({Key_s1[91], Key_s0[91]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_782, Feedback[27]}), .O ({new_AGEMA_signal_1088, AddRoundKeyOutput[27]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[28], Input_s0[28]}), .I1 ({Key_s1[28], Key_s0[28]}), .I2 ({Key_s1[92], Key_s0[92]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_787, Feedback[28]}), .O ({new_AGEMA_signal_1091, AddRoundKeyOutput[28]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[29], Input_s0[29]}), .I1 ({Key_s1[29], Key_s0[29]}), .I2 ({Key_s1[93], Key_s0[93]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_788, Feedback[29]}), .O ({new_AGEMA_signal_1094, AddRoundKeyOutput[29]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[2], Input_s0[2]}), .I1 ({Key_s1[2], Key_s0[2]}), .I2 ({Key_s1[66], Key_s0[66]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_733, Feedback[2]}), .O ({new_AGEMA_signal_1097, AddRoundKeyOutput[2]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[30], Input_s0[30]}), .I1 ({Key_s1[30], Key_s0[30]}), .I2 ({Key_s1[94], Key_s0[94]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_789, Feedback[30]}), .O ({new_AGEMA_signal_1100, AddRoundKeyOutput[30]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[7].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[31], Input_s0[31]}), .I1 ({Key_s1[31], Key_s0[31]}), .I2 ({Key_s1[95], Key_s0[95]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_790, Feedback[31]}), .O ({new_AGEMA_signal_1103, AddRoundKeyOutput[31]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[3], Input_s0[3]}), .I1 ({Key_s1[3], Key_s0[3]}), .I2 ({Key_s1[67], Key_s0[67]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_734, Feedback[3]}), .O ({new_AGEMA_signal_1106, AddRoundKeyOutput[3]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[4], Input_s0[4]}), .I1 ({Key_s1[4], Key_s0[4]}), .I2 ({Key_s1[68], Key_s0[68]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_739, Feedback[4]}), .O ({new_AGEMA_signal_1109, AddRoundKeyOutput[4]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[5], Input_s0[5]}), .I1 ({Key_s1[5], Key_s0[5]}), .I2 ({Key_s1[69], Key_s0[69]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_740, Feedback[5]}), .O ({new_AGEMA_signal_1112, AddRoundKeyOutput[5]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[6], Input_s0[6]}), .I1 ({Key_s1[6], Key_s0[6]}), .I2 ({Key_s1[70], Key_s0[70]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_741, Feedback[6]}), .O ({new_AGEMA_signal_1115, AddRoundKeyOutput[6]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[7], Input_s0[7]}), .I1 ({Key_s1[7], Key_s0[7]}), .I2 ({Key_s1[71], Key_s0[71]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_742, Feedback[7]}), .O ({new_AGEMA_signal_1118, AddRoundKeyOutput[7]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[8], Input_s0[8]}), .I1 ({Key_s1[8], Key_s0[8]}), .I2 ({Key_s1[72], Key_s0[72]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_747, Feedback[8]}), .O ({new_AGEMA_signal_1121, AddRoundKeyOutput[8]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h5A335A0F5ACC5AF0 ) , .MASK ( 6'b011000 ), .INIT2 ( 64'h5A335A0F5ACC5AF0 ) ) \AddKeyXOR2/GEN1[2].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[9], Input_s0[9]}), .I1 ({Key_s1[9], Key_s0[9]}), .I2 ({Key_s1[73], Key_s0[73]}), .I3 ({1'b0, rst}), .I4 ({1'b0, \selectsRegInst/s_current_state [0]}), .I5 ({new_AGEMA_signal_748, Feedback[9]}), .O ({new_AGEMA_signal_1124, AddRoundKeyOutput[9]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_935, N55}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [5]}), .I3 ({new_AGEMA_signal_932, N54}), .I4 ({new_AGEMA_signal_821, Feedback[46]}), .I5 ({new_AGEMA_signal_757, Feedback[14]}), .O ({new_AGEMA_signal_1125, AddRoundKeyOutput[46]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_941, N58}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [4]}), .I3 ({new_AGEMA_signal_938, N57}), .I4 ({new_AGEMA_signal_820, Feedback[45]}), .I5 ({new_AGEMA_signal_756, Feedback[13]}), .O ({new_AGEMA_signal_1126, AddRoundKeyOutput[45]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[32], Input_s0[32]}), .I1 ({Input_s1[0], Input_s0[0]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_857, N4}), .I4 ({new_AGEMA_signal_795, Feedback[32]}), .I5 ({new_AGEMA_signal_731, Feedback[0]}), .O ({new_AGEMA_signal_1128, AddRoundKeyOutput[32]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[33], Input_s0[33]}), .I1 ({Input_s1[1], Input_s0[1]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_860, N6}), .I4 ({new_AGEMA_signal_796, Feedback[33]}), .I5 ({new_AGEMA_signal_732, Feedback[1]}), .O ({new_AGEMA_signal_1130, AddRoundKeyOutput[33]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[34], Input_s0[34]}), .I1 ({Input_s1[2], Input_s0[2]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_863, N8}), .I4 ({new_AGEMA_signal_797, Feedback[34]}), .I5 ({new_AGEMA_signal_733, Feedback[2]}), .O ({new_AGEMA_signal_1132, AddRoundKeyOutput[34]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[8].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[35], Input_s0[35]}), .I1 ({Input_s1[3], Input_s0[3]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_866, N10}), .I4 ({new_AGEMA_signal_798, Feedback[35]}), .I5 ({new_AGEMA_signal_734, Feedback[3]}), .O ({new_AGEMA_signal_1134, AddRoundKeyOutput[35]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[36], Input_s0[36]}), .I1 ({Input_s1[4], Input_s0[4]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_869, N12}), .I4 ({new_AGEMA_signal_803, Feedback[36]}), .I5 ({new_AGEMA_signal_739, Feedback[4]}), .O ({new_AGEMA_signal_1136, AddRoundKeyOutput[36]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[37], Input_s0[37]}), .I1 ({Input_s1[5], Input_s0[5]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_872, N14}), .I4 ({new_AGEMA_signal_804, Feedback[37]}), .I5 ({new_AGEMA_signal_740, Feedback[5]}), .O ({new_AGEMA_signal_1138, AddRoundKeyOutput[37]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[38], Input_s0[38]}), .I1 ({Input_s1[6], Input_s0[6]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_875, N16}), .I4 ({new_AGEMA_signal_805, Feedback[38]}), .I5 ({new_AGEMA_signal_741, Feedback[6]}), .O ({new_AGEMA_signal_1140, AddRoundKeyOutput[38]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyXOR2/GEN1[9].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[39], Input_s0[39]}), .I1 ({Input_s1[7], Input_s0[7]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_878, N18}), .I4 ({new_AGEMA_signal_806, Feedback[39]}), .I5 ({new_AGEMA_signal_742, Feedback[7]}), .O ({new_AGEMA_signal_1142, AddRoundKeyOutput[39]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h609F6F906F90609F ) , .MASK ( 6'b000100 ), .INIT2 ( 64'h9F60906F906F9F60 ) ) \AddKeyConstXOR/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({Input_s1[43], Input_s0[43]}), .I1 ({Input_s1[11], Input_s0[11]}), .I2 ({1'b0, rst}), .I3 ({new_AGEMA_signal_881, N20}), .I4 ({new_AGEMA_signal_814, Feedback[43]}), .I5 ({new_AGEMA_signal_750, Feedback[11]}), .O ({new_AGEMA_signal_1144, AddRoundKeyOutput[43]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_975, N75}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_884, N22}), .I3 ({new_AGEMA_signal_827, Feedback[48]}), .I4 ({new_AGEMA_signal_763, Feedback[16]}), .I5 ({new_AGEMA_signal_731, Feedback[0]}), .O ({new_AGEMA_signal_1145, AddRoundKeyOutput[48]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_979, N77}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_887, N24}), .I3 ({new_AGEMA_signal_828, Feedback[49]}), .I4 ({new_AGEMA_signal_764, Feedback[17]}), .I5 ({new_AGEMA_signal_732, Feedback[1]}), .O ({new_AGEMA_signal_1146, AddRoundKeyOutput[49]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_983, N79}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_890, N26}), .I3 ({new_AGEMA_signal_829, Feedback[50]}), .I4 ({new_AGEMA_signal_765, Feedback[18]}), .I5 ({new_AGEMA_signal_733, Feedback[2]}), .O ({new_AGEMA_signal_1147, AddRoundKeyOutput[50]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[0].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_987, N81}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_893, N28}), .I3 ({new_AGEMA_signal_830, Feedback[51]}), .I4 ({new_AGEMA_signal_766, Feedback[19]}), .I5 ({new_AGEMA_signal_734, Feedback[3]}), .O ({new_AGEMA_signal_1148, AddRoundKeyOutput[51]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_991, N83}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_896, N30}), .I3 ({new_AGEMA_signal_835, Feedback[52]}), .I4 ({new_AGEMA_signal_771, Feedback[20]}), .I5 ({new_AGEMA_signal_739, Feedback[4]}), .O ({new_AGEMA_signal_1149, AddRoundKeyOutput[52]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_995, N85}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_899, N32}), .I3 ({new_AGEMA_signal_836, Feedback[53]}), .I4 ({new_AGEMA_signal_772, Feedback[21]}), .I5 ({new_AGEMA_signal_740, Feedback[5]}), .O ({new_AGEMA_signal_1150, AddRoundKeyOutput[53]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_999, N87}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_902, N34}), .I3 ({new_AGEMA_signal_837, Feedback[54]}), .I4 ({new_AGEMA_signal_773, Feedback[22]}), .I5 ({new_AGEMA_signal_741, Feedback[6]}), .O ({new_AGEMA_signal_1151, AddRoundKeyOutput[54]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1003, N89}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_905, N36}), .I3 ({new_AGEMA_signal_838, Feedback[55]}), .I4 ({new_AGEMA_signal_774, Feedback[23]}), .I5 ({new_AGEMA_signal_742, Feedback[7]}), .O ({new_AGEMA_signal_1152, AddRoundKeyOutput[55]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1006, N91}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_908, N38}), .I3 ({new_AGEMA_signal_843, Feedback[56]}), .I4 ({new_AGEMA_signal_779, Feedback[24]}), .I5 ({new_AGEMA_signal_747, Feedback[8]}), .O ({new_AGEMA_signal_1153, AddRoundKeyOutput[56]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1009, N93}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_911, N40}), .I3 ({new_AGEMA_signal_844, Feedback[57]}), .I4 ({new_AGEMA_signal_780, Feedback[25]}), .I5 ({new_AGEMA_signal_748, Feedback[9]}), .O ({new_AGEMA_signal_1154, AddRoundKeyOutput[57]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1012, N95}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_914, N42}), .I3 ({new_AGEMA_signal_845, Feedback[58]}), .I4 ({new_AGEMA_signal_781, Feedback[26]}), .I5 ({new_AGEMA_signal_749, Feedback[10]}), .O ({new_AGEMA_signal_1155, AddRoundKeyOutput[58]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[2].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1016, N97}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_917, N44}), .I3 ({new_AGEMA_signal_846, Feedback[59]}), .I4 ({new_AGEMA_signal_782, Feedback[27]}), .I5 ({new_AGEMA_signal_750, Feedback[11]}), .O ({new_AGEMA_signal_1156, AddRoundKeyOutput[59]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1019, N99}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_920, N46}), .I3 ({new_AGEMA_signal_851, Feedback[60]}), .I4 ({new_AGEMA_signal_787, Feedback[28]}), .I5 ({new_AGEMA_signal_755, Feedback[12]}), .O ({new_AGEMA_signal_1157, AddRoundKeyOutput[60]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1022, N101}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_923, N48}), .I3 ({new_AGEMA_signal_852, Feedback[61]}), .I4 ({new_AGEMA_signal_788, Feedback[29]}), .I5 ({new_AGEMA_signal_756, Feedback[13]}), .O ({new_AGEMA_signal_1158, AddRoundKeyOutput[61]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1025, N103}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_926, N50}), .I3 ({new_AGEMA_signal_853, Feedback[62]}), .I4 ({new_AGEMA_signal_789, Feedback[30]}), .I5 ({new_AGEMA_signal_757, Feedback[14]}), .O ({new_AGEMA_signal_1159, AddRoundKeyOutput[62]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'hB48787B487B4B487 ) , .MASK ( 6'b000010 ), .INIT2 ( 64'h4B78784B784B4B78 ) ) \AddKeyXOR1/GEN1[3].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_1028, N105}), .I1 ({1'b0, rst}), .I2 ({new_AGEMA_signal_929, N52}), .I3 ({new_AGEMA_signal_854, Feedback[63]}), .I4 ({new_AGEMA_signal_790, Feedback[31]}), .I5 ({new_AGEMA_signal_758, Feedback[15]}), .O ({new_AGEMA_signal_1160, AddRoundKeyOutput[63]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[3].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_947, N61}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [6]}), .I3 ({new_AGEMA_signal_944, N60}), .I4 ({new_AGEMA_signal_822, Feedback[47]}), .I5 ({new_AGEMA_signal_758, Feedback[15]}), .O ({new_AGEMA_signal_1161, AddRoundKeyOutput[47]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4774744774474774 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[1].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_953, N64}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [3]}), .I3 ({new_AGEMA_signal_950, N63}), .I4 ({new_AGEMA_signal_819, Feedback[44]}), .I5 ({new_AGEMA_signal_755, Feedback[12]}), .O ({new_AGEMA_signal_1162, AddRoundKeyOutput[44]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[0].GEN2[2].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_959, N67}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [2]}), .I3 ({new_AGEMA_signal_956, N66}), .I4 ({new_AGEMA_signal_813, Feedback[42]}), .I5 ({new_AGEMA_signal_749, Feedback[10]}), .O ({new_AGEMA_signal_1163, AddRoundKeyOutput[42]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h8BB8B88BB88B8BB8 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[0].GEN2[1].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_965, N70}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [1]}), .I3 ({new_AGEMA_signal_962, N69}), .I4 ({new_AGEMA_signal_812, Feedback[41]}), .I5 ({new_AGEMA_signal_748, Feedback[9]}), .O ({new_AGEMA_signal_1164, AddRoundKeyOutput[41]}) ) ;
    LUT6_masked #(.low_latency(0), .pipeline(0),  .INIT ( 64'h4774744774474774 ) , .MASK ( 6'b000110 ), .INIT2 ( 64'hBB8888BB88BBBB88 ) ) \AddKeyConstXOR/GEN1[0].GEN2[0].XORInst/Mxor_Q_xo<0>1 ( .I0 ({new_AGEMA_signal_971, N73}), .I1 ({1'b0, rst}), .I2 ({1'b0, \FSMRegInst/s_current_state [0]}), .I3 ({new_AGEMA_signal_968, N72}), .I4 ({new_AGEMA_signal_811, Feedback[40]}), .I5 ({new_AGEMA_signal_747, Feedback[8]}), .O ({new_AGEMA_signal_1165, AddRoundKeyOutput[40]}) ) ;

    /* register cells */
    FD done_2 ( .D (done_internal), .C (clk_gated), .Q (done) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_6 ( .D (\FSMUpdate [6]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [6]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_5 ( .D (\FSM [6]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [5]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_4 ( .D (\FSM [5]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [4]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_3 ( .D (\FSM [4]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [3]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_2 ( .D (\FSMUpdate [2]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [2]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_1 ( .D (\FSM [2]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [1]) ) ;
    FD #( .INIT ( 1'b0 ) ) \FSMRegInst/s_current_state_0 ( .D (\FSM [1]), .C (clk_gated), .Q (\FSMRegInst/s_current_state [0]) ) ;
    FD #( .INIT ( 1'b0 ) ) \selectsRegInst/s_current_state_0 ( .D (selectsNext[0]), .C (clk_gated), .Q (\selectsRegInst/s_current_state [0]) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_63 ( .D ({new_AGEMA_signal_1160, AddRoundKeyOutput[63]}), .clk (clk_gated), .Q ({Output_s1[63], Output_s0[63]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_62 ( .D ({new_AGEMA_signal_1159, AddRoundKeyOutput[62]}), .clk (clk_gated), .Q ({Output_s1[62], Output_s0[62]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_61 ( .D ({new_AGEMA_signal_1158, AddRoundKeyOutput[61]}), .clk (clk_gated), .Q ({Output_s1[61], Output_s0[61]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_60 ( .D ({new_AGEMA_signal_1157, AddRoundKeyOutput[60]}), .clk (clk_gated), .Q ({Output_s1[60], Output_s0[60]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_59 ( .D ({new_AGEMA_signal_1156, AddRoundKeyOutput[59]}), .clk (clk_gated), .Q ({Output_s1[59], Output_s0[59]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_58 ( .D ({new_AGEMA_signal_1155, AddRoundKeyOutput[58]}), .clk (clk_gated), .Q ({Output_s1[58], Output_s0[58]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_57 ( .D ({new_AGEMA_signal_1154, AddRoundKeyOutput[57]}), .clk (clk_gated), .Q ({Output_s1[57], Output_s0[57]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_56 ( .D ({new_AGEMA_signal_1153, AddRoundKeyOutput[56]}), .clk (clk_gated), .Q ({Output_s1[56], Output_s0[56]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_55 ( .D ({new_AGEMA_signal_1152, AddRoundKeyOutput[55]}), .clk (clk_gated), .Q ({Output_s1[55], Output_s0[55]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_54 ( .D ({new_AGEMA_signal_1151, AddRoundKeyOutput[54]}), .clk (clk_gated), .Q ({Output_s1[54], Output_s0[54]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_53 ( .D ({new_AGEMA_signal_1150, AddRoundKeyOutput[53]}), .clk (clk_gated), .Q ({Output_s1[53], Output_s0[53]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_52 ( .D ({new_AGEMA_signal_1149, AddRoundKeyOutput[52]}), .clk (clk_gated), .Q ({Output_s1[52], Output_s0[52]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_51 ( .D ({new_AGEMA_signal_1148, AddRoundKeyOutput[51]}), .clk (clk_gated), .Q ({Output_s1[51], Output_s0[51]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_50 ( .D ({new_AGEMA_signal_1147, AddRoundKeyOutput[50]}), .clk (clk_gated), .Q ({Output_s1[50], Output_s0[50]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_49 ( .D ({new_AGEMA_signal_1146, AddRoundKeyOutput[49]}), .clk (clk_gated), .Q ({Output_s1[49], Output_s0[49]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_48 ( .D ({new_AGEMA_signal_1145, AddRoundKeyOutput[48]}), .clk (clk_gated), .Q ({Output_s1[48], Output_s0[48]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_47 ( .D ({new_AGEMA_signal_1161, AddRoundKeyOutput[47]}), .clk (clk_gated), .Q ({Output_s1[47], Output_s0[47]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_46 ( .D ({new_AGEMA_signal_1125, AddRoundKeyOutput[46]}), .clk (clk_gated), .Q ({Output_s1[46], Output_s0[46]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_45 ( .D ({new_AGEMA_signal_1126, AddRoundKeyOutput[45]}), .clk (clk_gated), .Q ({Output_s1[45], Output_s0[45]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_44 ( .D ({new_AGEMA_signal_1162, AddRoundKeyOutput[44]}), .clk (clk_gated), .Q ({Output_s1[44], Output_s0[44]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_43 ( .D ({new_AGEMA_signal_1144, AddRoundKeyOutput[43]}), .clk (clk_gated), .Q ({Output_s1[43], Output_s0[43]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_42 ( .D ({new_AGEMA_signal_1163, AddRoundKeyOutput[42]}), .clk (clk_gated), .Q ({Output_s1[42], Output_s0[42]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_41 ( .D ({new_AGEMA_signal_1164, AddRoundKeyOutput[41]}), .clk (clk_gated), .Q ({Output_s1[41], Output_s0[41]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_40 ( .D ({new_AGEMA_signal_1165, AddRoundKeyOutput[40]}), .clk (clk_gated), .Q ({Output_s1[40], Output_s0[40]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_39 ( .D ({new_AGEMA_signal_1142, AddRoundKeyOutput[39]}), .clk (clk_gated), .Q ({Output_s1[39], Output_s0[39]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_38 ( .D ({new_AGEMA_signal_1140, AddRoundKeyOutput[38]}), .clk (clk_gated), .Q ({Output_s1[38], Output_s0[38]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_37 ( .D ({new_AGEMA_signal_1138, AddRoundKeyOutput[37]}), .clk (clk_gated), .Q ({Output_s1[37], Output_s0[37]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_36 ( .D ({new_AGEMA_signal_1136, AddRoundKeyOutput[36]}), .clk (clk_gated), .Q ({Output_s1[36], Output_s0[36]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_35 ( .D ({new_AGEMA_signal_1134, AddRoundKeyOutput[35]}), .clk (clk_gated), .Q ({Output_s1[35], Output_s0[35]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_34 ( .D ({new_AGEMA_signal_1132, AddRoundKeyOutput[34]}), .clk (clk_gated), .Q ({Output_s1[34], Output_s0[34]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_33 ( .D ({new_AGEMA_signal_1130, AddRoundKeyOutput[33]}), .clk (clk_gated), .Q ({Output_s1[33], Output_s0[33]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_32 ( .D ({new_AGEMA_signal_1128, AddRoundKeyOutput[32]}), .clk (clk_gated), .Q ({Output_s1[32], Output_s0[32]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_31 ( .D ({new_AGEMA_signal_1103, AddRoundKeyOutput[31]}), .clk (clk_gated), .Q ({Output_s1[31], Output_s0[31]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_30 ( .D ({new_AGEMA_signal_1100, AddRoundKeyOutput[30]}), .clk (clk_gated), .Q ({Output_s1[30], Output_s0[30]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_29 ( .D ({new_AGEMA_signal_1094, AddRoundKeyOutput[29]}), .clk (clk_gated), .Q ({Output_s1[29], Output_s0[29]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_28 ( .D ({new_AGEMA_signal_1091, AddRoundKeyOutput[28]}), .clk (clk_gated), .Q ({Output_s1[28], Output_s0[28]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_27 ( .D ({new_AGEMA_signal_1088, AddRoundKeyOutput[27]}), .clk (clk_gated), .Q ({Output_s1[27], Output_s0[27]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_26 ( .D ({new_AGEMA_signal_1085, AddRoundKeyOutput[26]}), .clk (clk_gated), .Q ({Output_s1[26], Output_s0[26]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_25 ( .D ({new_AGEMA_signal_1082, AddRoundKeyOutput[25]}), .clk (clk_gated), .Q ({Output_s1[25], Output_s0[25]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_24 ( .D ({new_AGEMA_signal_1079, AddRoundKeyOutput[24]}), .clk (clk_gated), .Q ({Output_s1[24], Output_s0[24]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_23 ( .D ({new_AGEMA_signal_1076, AddRoundKeyOutput[23]}), .clk (clk_gated), .Q ({Output_s1[23], Output_s0[23]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_22 ( .D ({new_AGEMA_signal_1073, AddRoundKeyOutput[22]}), .clk (clk_gated), .Q ({Output_s1[22], Output_s0[22]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_21 ( .D ({new_AGEMA_signal_1070, AddRoundKeyOutput[21]}), .clk (clk_gated), .Q ({Output_s1[21], Output_s0[21]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_20 ( .D ({new_AGEMA_signal_1067, AddRoundKeyOutput[20]}), .clk (clk_gated), .Q ({Output_s1[20], Output_s0[20]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_19 ( .D ({new_AGEMA_signal_1061, AddRoundKeyOutput[19]}), .clk (clk_gated), .Q ({Output_s1[19], Output_s0[19]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_18 ( .D ({new_AGEMA_signal_1058, AddRoundKeyOutput[18]}), .clk (clk_gated), .Q ({Output_s1[18], Output_s0[18]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_17 ( .D ({new_AGEMA_signal_1055, AddRoundKeyOutput[17]}), .clk (clk_gated), .Q ({Output_s1[17], Output_s0[17]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_16 ( .D ({new_AGEMA_signal_1052, AddRoundKeyOutput[16]}), .clk (clk_gated), .Q ({Output_s1[16], Output_s0[16]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_15 ( .D ({new_AGEMA_signal_1049, AddRoundKeyOutput[15]}), .clk (clk_gated), .Q ({Output_s1[15], Output_s0[15]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_14 ( .D ({new_AGEMA_signal_1046, AddRoundKeyOutput[14]}), .clk (clk_gated), .Q ({Output_s1[14], Output_s0[14]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_13 ( .D ({new_AGEMA_signal_1043, AddRoundKeyOutput[13]}), .clk (clk_gated), .Q ({Output_s1[13], Output_s0[13]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_12 ( .D ({new_AGEMA_signal_1040, AddRoundKeyOutput[12]}), .clk (clk_gated), .Q ({Output_s1[12], Output_s0[12]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_11 ( .D ({new_AGEMA_signal_1037, AddRoundKeyOutput[11]}), .clk (clk_gated), .Q ({Output_s1[11], Output_s0[11]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_10 ( .D ({new_AGEMA_signal_1034, AddRoundKeyOutput[10]}), .clk (clk_gated), .Q ({Output_s1[10], Output_s0[10]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_9 ( .D ({new_AGEMA_signal_1124, AddRoundKeyOutput[9]}), .clk (clk_gated), .Q ({Output_s1[9], Output_s0[9]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_8 ( .D ({new_AGEMA_signal_1121, AddRoundKeyOutput[8]}), .clk (clk_gated), .Q ({Output_s1[8], Output_s0[8]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_7 ( .D ({new_AGEMA_signal_1118, AddRoundKeyOutput[7]}), .clk (clk_gated), .Q ({Output_s1[7], Output_s0[7]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_6 ( .D ({new_AGEMA_signal_1115, AddRoundKeyOutput[6]}), .clk (clk_gated), .Q ({Output_s1[6], Output_s0[6]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_5 ( .D ({new_AGEMA_signal_1112, AddRoundKeyOutput[5]}), .clk (clk_gated), .Q ({Output_s1[5], Output_s0[5]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_4 ( .D ({new_AGEMA_signal_1109, AddRoundKeyOutput[4]}), .clk (clk_gated), .Q ({Output_s1[4], Output_s0[4]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_3 ( .D ({new_AGEMA_signal_1106, AddRoundKeyOutput[3]}), .clk (clk_gated), .Q ({Output_s1[3], Output_s0[3]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_2 ( .D ({new_AGEMA_signal_1097, AddRoundKeyOutput[2]}), .clk (clk_gated), .Q ({Output_s1[2], Output_s0[2]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_1 ( .D ({new_AGEMA_signal_1064, AddRoundKeyOutput[1]}), .clk (clk_gated), .Q ({Output_s1[1], Output_s0[1]}) ) ;
    FD_masked #(.low_latency(0), .pipeline(0),  .INIT ( 1'b0 ) ) \StateReg/s_current_state_0 ( .D ({new_AGEMA_signal_1031, AddRoundKeyOutput[0]}), .clk (clk_gated), .Q ({Output_s1[0], Output_s0[0]}) ) ;
endmodule
