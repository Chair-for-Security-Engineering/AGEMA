/* modified netlist. Source: module AES in file AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_HPC3_Pipeline_d2 (plaintext_s0, key_s0, clk, reset, plaintext_s1, plaintext_s2, key_s1, key_s2, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [815:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    wire AKSRnotDone ;
    wire LastRoundorDone ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire n55 ;
    wire n56 ;
    wire n57 ;
    wire n58 ;
    wire n59 ;
    wire n60 ;
    wire n61 ;
    wire n62 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire MuxSboxIn_n7 ;
    wire MuxSboxIn_n6 ;
    wire MuxSboxIn_n5 ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire MixColumnsIns_n64 ;
    wire MixColumnsIns_n63 ;
    wire MixColumnsIns_n62 ;
    wire MixColumnsIns_n61 ;
    wire MixColumnsIns_n60 ;
    wire MixColumnsIns_n59 ;
    wire MixColumnsIns_n58 ;
    wire MixColumnsIns_n57 ;
    wire MixColumnsIns_n56 ;
    wire MixColumnsIns_n55 ;
    wire MixColumnsIns_n54 ;
    wire MixColumnsIns_n53 ;
    wire MixColumnsIns_n52 ;
    wire MixColumnsIns_n51 ;
    wire MixColumnsIns_n50 ;
    wire MixColumnsIns_n49 ;
    wire MixColumnsIns_n48 ;
    wire MixColumnsIns_n47 ;
    wire MixColumnsIns_n46 ;
    wire MixColumnsIns_n45 ;
    wire MixColumnsIns_n44 ;
    wire MixColumnsIns_n43 ;
    wire MixColumnsIns_n42 ;
    wire MixColumnsIns_n41 ;
    wire MixColumnsIns_n40 ;
    wire MixColumnsIns_n39 ;
    wire MixColumnsIns_n38 ;
    wire MixColumnsIns_n37 ;
    wire MixColumnsIns_n36 ;
    wire MixColumnsIns_n35 ;
    wire MixColumnsIns_n34 ;
    wire MixColumnsIns_n33 ;
    wire MixColumnsIns_n32 ;
    wire MixColumnsIns_n31 ;
    wire MixColumnsIns_n30 ;
    wire MixColumnsIns_n29 ;
    wire MixColumnsIns_n28 ;
    wire MixColumnsIns_n27 ;
    wire MixColumnsIns_n26 ;
    wire MixColumnsIns_n25 ;
    wire MixColumnsIns_n24 ;
    wire MixColumnsIns_n23 ;
    wire MixColumnsIns_n22 ;
    wire MixColumnsIns_n21 ;
    wire MixColumnsIns_n20 ;
    wire MixColumnsIns_n19 ;
    wire MixColumnsIns_n18 ;
    wire MixColumnsIns_n17 ;
    wire MixColumnsIns_n16 ;
    wire MixColumnsIns_n15 ;
    wire MixColumnsIns_n14 ;
    wire MixColumnsIns_n13 ;
    wire MixColumnsIns_n12 ;
    wire MixColumnsIns_n11 ;
    wire MixColumnsIns_n10 ;
    wire MixColumnsIns_n9 ;
    wire MixColumnsIns_n8 ;
    wire MixColumnsIns_n7 ;
    wire MixColumnsIns_n6 ;
    wire MixColumnsIns_n5 ;
    wire MixColumnsIns_n4 ;
    wire MixColumnsIns_n3 ;
    wire MixColumnsIns_n2 ;
    wire MixColumnsIns_n1 ;
    wire MuxMCOut_n6 ;
    wire MuxMCOut_n5 ;
    wire MuxMCOut_n4 ;
    wire MuxRound_n19 ;
    wire MuxRound_n18 ;
    wire MuxRound_n17 ;
    wire MuxRound_n16 ;
    wire MuxRound_n15 ;
    wire MuxRound_n14 ;
    wire MuxRound_n13 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire MuxKeyExpansion_n21 ;
    wire MuxKeyExpansion_n20 ;
    wire MuxKeyExpansion_n19 ;
    wire MuxKeyExpansion_n18 ;
    wire MuxKeyExpansion_n17 ;
    wire MuxKeyExpansion_n16 ;
    wire MuxKeyExpansion_n15 ;
    wire MuxKeyExpansion_n14 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n42 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n44 ;
    wire RoundCounterIns_n45 ;
    wire InRoundCounterIns_n12 ;
    wire InRoundCounterIns_n11 ;
    wire InRoundCounterIns_n10 ;
    wire InRoundCounterIns_n9 ;
    wire InRoundCounterIns_n8 ;
    wire InRoundCounterIns_n7 ;
    wire InRoundCounterIns_n5 ;
    wire InRoundCounterIns_n4 ;
    wire InRoundCounterIns_n3 ;
    wire InRoundCounterIns_n2 ;
    wire InRoundCounterIns_n1 ;
    wire InRoundCounterIns_n6 ;
    wire InRoundCounterIns_n39 ;
    wire InRoundCounterIns_n40 ;
    wire InRoundCounterIns_n41 ;
    wire [127:0] RoundOutput ;
    wire [127:0] ShiftRowsOutput ;
    wire [31:0] KSSubBytesInput ;
    wire [31:0] SubBytesInput ;
    wire [3:0] SubBytesOutput ;
    wire [31:0] MixColumnsOutput ;
    wire [31:0] ColumnOutput ;
    wire [127:0] RoundKeyOutput ;
    wire [127:32] RoundKey ;
    wire [7:0] Rcon ;
    wire [127:0] KeyExpansionOutput ;
    wire [3:0] RoundCounter ;
    wire [2:0] InRoundCounter ;
    wire [28:0] MixColumnsIns_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;

    /* cells in depth 0 */
    AND2_X1 U323 ( .A1 (n45), .A2 (n44), .ZN (AKSRnotDone) ) ;
    NOR2_X1 U324 ( .A1 (n60), .A2 (n49), .ZN (LastRoundorDone) ) ;
    AND2_X1 U325 ( .A1 (RoundCounter[0]), .A2 (LastRoundorDone), .ZN (done) ) ;
    INV_X1 U326 ( .A (RoundCounter[3]), .ZN (n60) ) ;
    NOR2_X1 U327 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (n45) ) ;
    INV_X1 U328 ( .A (RoundCounter[2]), .ZN (n46) ) ;
    NAND2_X1 U329 ( .A1 (RoundCounter[1]), .A2 (n46), .ZN (n49) ) ;
    NOR2_X1 U330 ( .A1 (done), .A2 (InRoundCounter[2]), .ZN (n44) ) ;
    INV_X1 U331 ( .A (RoundCounter[1]), .ZN (n55) ) ;
    NAND2_X1 U332 ( .A1 (n55), .A2 (n46), .ZN (n47) ) ;
    NOR2_X1 U333 ( .A1 (RoundCounter[0]), .A2 (n47), .ZN (Rcon[0]) ) ;
    NOR2_X1 U334 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n58) ) ;
    NOR2_X1 U335 ( .A1 (n58), .A2 (n47), .ZN (Rcon[1]) ) ;
    NOR2_X1 U336 ( .A1 (RoundCounter[3]), .A2 (n49), .ZN (n48) ) ;
    NOR2_X1 U337 ( .A1 (n60), .A2 (n47), .ZN (n54) ) ;
    MUX2_X1 U338 ( .S (RoundCounter[0]), .A (n48), .B (n54), .Z (Rcon[2]) ) ;
    INV_X1 U339 ( .A (RoundCounter[0]), .ZN (n50) ) ;
    NOR2_X1 U340 ( .A1 (n50), .A2 (n49), .ZN (n51) ) ;
    MUX2_X1 U341 ( .S (RoundCounter[3]), .A (n51), .B (Rcon[0]), .Z (Rcon[3]) ) ;
    NAND2_X1 U342 ( .A1 (RoundCounter[2]), .A2 (n58), .ZN (n52) ) ;
    NOR2_X1 U343 ( .A1 (RoundCounter[1]), .A2 (n52), .ZN (n53) ) ;
    OR2_X1 U344 ( .A1 (n54), .A2 (n53), .ZN (Rcon[4]) ) ;
    XNOR2_X1 U345 ( .A (RoundCounter[2]), .B (RoundCounter[3]), .ZN (n57) ) ;
    NAND2_X1 U346 ( .A1 (RoundCounter[0]), .A2 (n55), .ZN (n56) ) ;
    NOR2_X1 U347 ( .A1 (n57), .A2 (n56), .ZN (Rcon[5]) ) ;
    INV_X1 U348 ( .A (n58), .ZN (n59) ) ;
    NAND2_X1 U349 ( .A1 (RoundCounter[1]), .A2 (RoundCounter[2]), .ZN (n61) ) ;
    NOR2_X1 U350 ( .A1 (n59), .A2 (n61), .ZN (Rcon[6]) ) ;
    NAND2_X1 U351 ( .A1 (RoundCounter[0]), .A2 (n60), .ZN (n62) ) ;
    NOR2_X1 U352 ( .A1 (n62), .A2 (n61), .ZN (Rcon[7]) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U353 ( .a ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, ShiftRowsOutput[96]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U354 ( .a ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, RoundKey[100]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, ShiftRowsOutput[68]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U355 ( .a ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, RoundKey[101]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, ShiftRowsOutput[69]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U356 ( .a ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, RoundKey[102]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, ShiftRowsOutput[70]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U357 ( .a ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, RoundKey[103]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, ShiftRowsOutput[71]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U358 ( .a ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, RoundKey[104]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, ShiftRowsOutput[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U359 ( .a ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, RoundKey[105]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U360 ( .a ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, RoundKey[106]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, ShiftRowsOutput[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U361 ( .a ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, RoundKey[107]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U362 ( .a ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, RoundKey[108]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, ShiftRowsOutput[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U363 ( .a ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, RoundKey[109]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U364 ( .a ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, ShiftRowsOutput[74]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U365 ( .a ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, RoundKey[110]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, ShiftRowsOutput[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U366 ( .a ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, RoundKey[111]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, ShiftRowsOutput[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U367 ( .a ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, RoundKey[112]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, ShiftRowsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U368 ( .a ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, RoundKey[113]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, ShiftRowsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U369 ( .a ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, RoundKey[114]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, ShiftRowsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U370 ( .a ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, RoundKey[115]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, ShiftRowsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U371 ( .a ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, RoundKey[116]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, ShiftRowsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U372 ( .a ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, RoundKey[117]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, ShiftRowsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U373 ( .a ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, RoundKey[118]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, ShiftRowsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U374 ( .a ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, RoundKey[119]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, ShiftRowsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U375 ( .a ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, ShiftRowsOutput[75]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U376 ( .a ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, RoundKey[120]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, ShiftRowsOutput[120]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U377 ( .a ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, RoundKey[121]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, ShiftRowsOutput[121]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U378 ( .a ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, RoundKey[122]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[122]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U379 ( .a ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, RoundKey[123]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[123]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U380 ( .a ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, RoundKey[124]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, ShiftRowsOutput[124]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U381 ( .a ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, RoundKey[125]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, ShiftRowsOutput[125]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U382 ( .a ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, RoundKey[126]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, ShiftRowsOutput[126]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U383 ( .a ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, RoundKey[127]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, ShiftRowsOutput[127]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U384 ( .a ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, ShiftRowsOutput[76]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U385 ( .a ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[77]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U386 ( .a ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, ShiftRowsOutput[78]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U387 ( .a ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, ShiftRowsOutput[79]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U388 ( .a ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, ShiftRowsOutput[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U389 ( .a ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, ShiftRowsOutput[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U390 ( .a ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, ShiftRowsOutput[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U391 ( .a ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, ShiftRowsOutput[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U392 ( .a ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, ShiftRowsOutput[97]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U393 ( .a ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, ShiftRowsOutput[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U394 ( .a ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, ShiftRowsOutput[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U395 ( .a ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U396 ( .a ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, ShiftRowsOutput[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U397 ( .a ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, ShiftRowsOutput[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U398 ( .a ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, ShiftRowsOutput[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U399 ( .a ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, ShiftRowsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U400 ( .a ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, ShiftRowsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U401 ( .a ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, ShiftRowsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U402 ( .a ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, ShiftRowsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U403 ( .a ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, ShiftRowsOutput[98]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U404 ( .a ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, ShiftRowsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U405 ( .a ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, ShiftRowsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U406 ( .a ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, RoundKey[32]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, ShiftRowsOutput[0]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U407 ( .a ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, RoundKey[33]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, ShiftRowsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U408 ( .a ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, RoundKey[34]}), .c ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, ShiftRowsOutput[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U409 ( .a ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, RoundKey[35]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, ShiftRowsOutput[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U410 ( .a ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, RoundKey[36]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, ShiftRowsOutput[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U411 ( .a ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, RoundKey[37]}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, ShiftRowsOutput[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U412 ( .a ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, RoundKey[38]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, ShiftRowsOutput[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U413 ( .a ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, RoundKey[39]}), .c ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, ShiftRowsOutput[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U414 ( .a ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, ShiftRowsOutput[99]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U415 ( .a ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, RoundKey[40]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, ShiftRowsOutput[104]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U416 ( .a ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, RoundKey[41]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, ShiftRowsOutput[105]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U417 ( .a ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, RoundKey[42]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, ShiftRowsOutput[106]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U418 ( .a ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, RoundKey[43]}), .c ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, ShiftRowsOutput[107]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U419 ( .a ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, RoundKey[44]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[108]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U420 ( .a ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, RoundKey[45]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, ShiftRowsOutput[109]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U421 ( .a ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, RoundKey[46]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, ShiftRowsOutput[110]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U422 ( .a ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, RoundKey[47]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, ShiftRowsOutput[111]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U423 ( .a ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, RoundKey[48]}), .c ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, ShiftRowsOutput[80]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U424 ( .a ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, RoundKey[49]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, ShiftRowsOutput[81]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U425 ( .a ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, ShiftRowsOutput[100]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U426 ( .a ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, RoundKey[50]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, ShiftRowsOutput[82]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U427 ( .a ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, RoundKey[51]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, ShiftRowsOutput[83]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U428 ( .a ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, RoundKey[52]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, ShiftRowsOutput[84]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U429 ( .a ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, RoundKey[53]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, ShiftRowsOutput[85]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U430 ( .a ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, RoundKey[54]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, ShiftRowsOutput[86]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U431 ( .a ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, RoundKey[55]}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, ShiftRowsOutput[87]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U432 ( .a ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, RoundKey[56]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, ShiftRowsOutput[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U433 ( .a ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, RoundKey[57]}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, ShiftRowsOutput[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U434 ( .a ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, RoundKey[58]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, ShiftRowsOutput[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U435 ( .a ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, RoundKey[59]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, ShiftRowsOutput[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U436 ( .a ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, ShiftRowsOutput[101]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U437 ( .a ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, RoundKey[60]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, ShiftRowsOutput[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U438 ( .a ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, RoundKey[61]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, ShiftRowsOutput[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U439 ( .a ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, RoundKey[62]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, ShiftRowsOutput[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U440 ( .a ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, RoundKey[63]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, ShiftRowsOutput[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U441 ( .a ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, RoundKey[64]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, ShiftRowsOutput[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U442 ( .a ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, RoundKey[65]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, ShiftRowsOutput[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U443 ( .a ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, RoundKey[66]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, ShiftRowsOutput[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U444 ( .a ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, RoundKey[67]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, ShiftRowsOutput[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U445 ( .a ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, RoundKey[68]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, ShiftRowsOutput[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U446 ( .a ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, RoundKey[69]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, ShiftRowsOutput[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U447 ( .a ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, ShiftRowsOutput[102]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U448 ( .a ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, RoundKey[70]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, ShiftRowsOutput[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U449 ( .a ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, RoundKey[71]}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, ShiftRowsOutput[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U450 ( .a ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, RoundKey[72]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, ShiftRowsOutput[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U451 ( .a ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, RoundKey[73]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, ShiftRowsOutput[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U452 ( .a ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, RoundKey[74]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, ShiftRowsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U453 ( .a ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, RoundKey[75]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, ShiftRowsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U454 ( .a ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, RoundKey[76]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, ShiftRowsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U455 ( .a ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, RoundKey[77]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, ShiftRowsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U456 ( .a ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, RoundKey[78]}), .c ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, ShiftRowsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U457 ( .a ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, RoundKey[79]}), .c ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, ShiftRowsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U458 ( .a ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, ShiftRowsOutput[103]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U459 ( .a ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, RoundKey[80]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, ShiftRowsOutput[112]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U460 ( .a ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, RoundKey[81]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, ShiftRowsOutput[113]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U461 ( .a ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, RoundKey[82]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, ShiftRowsOutput[114]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U462 ( .a ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, RoundKey[83]}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, ShiftRowsOutput[115]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U463 ( .a ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, RoundKey[84]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, ShiftRowsOutput[116]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U464 ( .a ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, RoundKey[85]}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, ShiftRowsOutput[117]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U465 ( .a ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, RoundKey[86]}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, ShiftRowsOutput[118]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U466 ( .a ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, RoundKey[87]}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, ShiftRowsOutput[119]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U467 ( .a ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, RoundKey[88]}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, ShiftRowsOutput[88]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U468 ( .a ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, RoundKey[89]}), .c ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, ShiftRowsOutput[89]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U469 ( .a ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, ShiftRowsOutput[72]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U470 ( .a ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, RoundKey[90]}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, ShiftRowsOutput[90]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U471 ( .a ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, RoundKey[91]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, ShiftRowsOutput[91]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U472 ( .a ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, RoundKey[92]}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, ShiftRowsOutput[92]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U473 ( .a ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, RoundKey[93]}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, ShiftRowsOutput[93]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U474 ( .a ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, RoundKey[94]}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, ShiftRowsOutput[94]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U475 ( .a ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, RoundKey[95]}), .c ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, ShiftRowsOutput[95]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U476 ( .a ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, RoundKey[96]}), .c ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, ShiftRowsOutput[64]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U477 ( .a ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, RoundKey[97]}), .c ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, ShiftRowsOutput[65]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U478 ( .a ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, RoundKey[98]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, ShiftRowsOutput[66]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U479 ( .a ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, RoundKey[99]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, ShiftRowsOutput[67]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) U480 ( .a ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, ShiftRowsOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, RoundOutput[32]}), .a ({plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, RoundOutput[33]}), .a ({plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, RoundOutput[34]}), .a ({plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, RoundOutput[35]}), .a ({plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, RoundOutput[36]}), .a ({plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, RoundOutput[37]}), .a ({plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, RoundOutput[38]}), .a ({plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, RoundOutput[39]}), .a ({plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, RoundOutput[40]}), .a ({plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, RoundOutput[41]}), .a ({plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, RoundOutput[42]}), .a ({plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, RoundOutput[43]}), .a ({plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, RoundOutput[44]}), .a ({plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, RoundOutput[45]}), .a ({plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, RoundOutput[46]}), .a ({plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, RoundOutput[47]}), .a ({plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, RoundOutput[48]}), .a ({plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, RoundOutput[49]}), .a ({plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, RoundOutput[50]}), .a ({plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, RoundOutput[51]}), .a ({plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, RoundOutput[52]}), .a ({plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, RoundOutput[53]}), .a ({plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, RoundOutput[54]}), .a ({plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, RoundOutput[55]}), .a ({plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, RoundOutput[56]}), .a ({plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, RoundOutput[57]}), .a ({plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, RoundOutput[58]}), .a ({plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, RoundOutput[59]}), .a ({plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, RoundOutput[60]}), .a ({plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, RoundOutput[61]}), .a ({plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, RoundOutput[62]}), .a ({plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, RoundOutput[63]}), .a ({plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, RoundOutput[64]}), .a ({plaintext_s2[64], plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, RoundOutput[65]}), .a ({plaintext_s2[65], plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, RoundOutput[66]}), .a ({plaintext_s2[66], plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, RoundOutput[67]}), .a ({plaintext_s2[67], plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, RoundOutput[68]}), .a ({plaintext_s2[68], plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, RoundOutput[69]}), .a ({plaintext_s2[69], plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, RoundOutput[70]}), .a ({plaintext_s2[70], plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, RoundOutput[71]}), .a ({plaintext_s2[71], plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, RoundOutput[72]}), .a ({plaintext_s2[72], plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, RoundOutput[73]}), .a ({plaintext_s2[73], plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, RoundOutput[74]}), .a ({plaintext_s2[74], plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, RoundOutput[75]}), .a ({plaintext_s2[75], plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, RoundOutput[76]}), .a ({plaintext_s2[76], plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, RoundOutput[77]}), .a ({plaintext_s2[77], plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, RoundOutput[78]}), .a ({plaintext_s2[78], plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, RoundOutput[79]}), .a ({plaintext_s2[79], plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, RoundOutput[80]}), .a ({plaintext_s2[80], plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, RoundOutput[81]}), .a ({plaintext_s2[81], plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, RoundOutput[82]}), .a ({plaintext_s2[82], plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, RoundOutput[83]}), .a ({plaintext_s2[83], plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, RoundOutput[84]}), .a ({plaintext_s2[84], plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, RoundOutput[85]}), .a ({plaintext_s2[85], plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, RoundOutput[86]}), .a ({plaintext_s2[86], plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, RoundOutput[87]}), .a ({plaintext_s2[87], plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, RoundOutput[88]}), .a ({plaintext_s2[88], plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, RoundOutput[89]}), .a ({plaintext_s2[89], plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, RoundOutput[90]}), .a ({plaintext_s2[90], plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, RoundOutput[91]}), .a ({plaintext_s2[91], plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, RoundOutput[92]}), .a ({plaintext_s2[92], plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, RoundOutput[93]}), .a ({plaintext_s2[93], plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, RoundOutput[94]}), .a ({plaintext_s2[94], plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, RoundOutput[95]}), .a ({plaintext_s2[95], plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, RoundOutput[96]}), .a ({plaintext_s2[96], plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, RoundOutput[97]}), .a ({plaintext_s2[97], plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, RoundOutput[98]}), .a ({plaintext_s2[98], plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, RoundOutput[99]}), .a ({plaintext_s2[99], plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, RoundOutput[100]}), .a ({plaintext_s2[100], plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, RoundOutput[101]}), .a ({plaintext_s2[101], plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, RoundOutput[102]}), .a ({plaintext_s2[102], plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, RoundOutput[103]}), .a ({plaintext_s2[103], plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, RoundOutput[104]}), .a ({plaintext_s2[104], plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, RoundOutput[105]}), .a ({plaintext_s2[105], plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, RoundOutput[106]}), .a ({plaintext_s2[106], plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, RoundOutput[107]}), .a ({plaintext_s2[107], plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, RoundOutput[108]}), .a ({plaintext_s2[108], plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, RoundOutput[109]}), .a ({plaintext_s2[109], plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, RoundOutput[110]}), .a ({plaintext_s2[110], plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, RoundOutput[111]}), .a ({plaintext_s2[111], plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, RoundOutput[112]}), .a ({plaintext_s2[112], plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, RoundOutput[113]}), .a ({plaintext_s2[113], plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, RoundOutput[114]}), .a ({plaintext_s2[114], plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, RoundOutput[115]}), .a ({plaintext_s2[115], plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, RoundOutput[116]}), .a ({plaintext_s2[116], plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, RoundOutput[117]}), .a ({plaintext_s2[117], plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, RoundOutput[118]}), .a ({plaintext_s2[118], plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, RoundOutput[119]}), .a ({plaintext_s2[119], plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, RoundOutput[120]}), .a ({plaintext_s2[120], plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, RoundOutput[121]}), .a ({plaintext_s2[121], plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, RoundOutput[122]}), .a ({plaintext_s2[122], plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, RoundOutput[123]}), .a ({plaintext_s2[123], plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, RoundOutput[124]}), .a ({plaintext_s2[124], plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, RoundOutput[125]}), .a ({plaintext_s2[125], plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, RoundOutput[126]}), .a ({plaintext_s2[126], plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, RoundOutput[127]}), .a ({plaintext_s2[127], plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    INV_X1 MuxSboxIn_U3 ( .A (AKSRnotDone), .ZN (MuxSboxIn_n7) ) ;
    INV_X1 MuxSboxIn_U2 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n5) ) ;
    INV_X1 MuxSboxIn_U1 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n6) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_0_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .a ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_1_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_2_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_3_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, SubBytesInput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_4_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_5_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, SubBytesInput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_6_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .a ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, SubBytesInput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_7_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_8_U1 ( .s (AKSRnotDone), .b ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_9_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_10_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .a ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_11_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, SubBytesInput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_12_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .a ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_13_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, SubBytesInput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_14_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .a ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, SubBytesInput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_15_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_16_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .a ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_17_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .a ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_18_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_19_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .a ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, SubBytesInput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_20_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .a ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_21_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, SubBytesInput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_22_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .a ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, SubBytesInput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_23_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .a ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_24_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .a ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_25_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_26_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_27_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, SubBytesInput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_28_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .a ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_29_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, SubBytesInput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_30_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, SubBytesInput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxSboxIn_mux_inst_31_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .a ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}), .b ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, SubBytesInput[7]}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}), .c ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, SubBytesInput[3]}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, SubBytesInput[6]}), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, SubBytesInput[5]}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .b ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .b ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, SubBytesInput[6]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, SubBytesInput[5]}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, SubBytesInput[2]}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, SubBytesInput[4]}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .c ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, SubBytesInput[1]}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, SubBytesInput[15]}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, SubBytesInput[11]}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, SubBytesInput[14]}), .b ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, SubBytesInput[13]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, SubBytesInput[14]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, SubBytesInput[13]}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, SubBytesInput[10]}), .c ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, SubBytesInput[12]}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, SubBytesInput[9]}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .c ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}), .b ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}), .c ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, SubBytesInput[23]}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}), .c ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, SubBytesInput[19]}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, SubBytesInput[22]}), .b ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, SubBytesInput[21]}), .c ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .b ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, SubBytesInput[22]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, SubBytesInput[21]}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, SubBytesInput[18]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, SubBytesInput[20]}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .c ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, SubBytesInput[17]}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .c ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_4031, new_AGEMA_signal_4030, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, SubBytesInput[31]}), .b ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, SubBytesInput[27]}), .b ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}), .c ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, SubBytesInput[30]}), .b ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, SubBytesInput[29]}), .c ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, SubBytesInput[30]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, SubBytesInput[29]}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, SubBytesInput[26]}), .c ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, SubBytesInput[28]}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .c ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, SubBytesInput[25]}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    INV_X1 MuxMCOut_U3 ( .A (LastRoundorDone), .ZN (MuxMCOut_n6) ) ;
    INV_X1 MuxMCOut_U2 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n5) ) ;
    INV_X1 MuxMCOut_U1 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n4) ) ;
    INV_X1 MuxRound_U7 ( .A (AKSRnotDone), .ZN (MuxRound_n19) ) ;
    INV_X1 MuxRound_U6 ( .A (MuxRound_n19), .ZN (MuxRound_n16) ) ;
    INV_X1 MuxRound_U5 ( .A (MuxRound_n19), .ZN (MuxRound_n14) ) ;
    INV_X1 MuxRound_U4 ( .A (MuxRound_n19), .ZN (MuxRound_n13) ) ;
    INV_X1 MuxRound_U3 ( .A (MuxRound_n19), .ZN (MuxRound_n15) ) ;
    INV_X1 MuxRound_U2 ( .A (MuxRound_n19), .ZN (MuxRound_n18) ) ;
    INV_X1 MuxRound_U1 ( .A (MuxRound_n19), .ZN (MuxRound_n17) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_32_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_33_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .a ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_34_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .a ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_35_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .a ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_36_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_37_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .a ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_38_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .a ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_39_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_40_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .a ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_41_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_42_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .a ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_43_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_44_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .a ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_45_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_46_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_47_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .a ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_48_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .a ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, ShiftRowsOutput[48]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_49_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, ShiftRowsOutput[49]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_50_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .a ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, ShiftRowsOutput[50]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_51_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .a ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, ShiftRowsOutput[51]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_52_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .a ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, ShiftRowsOutput[52]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_53_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .a ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, ShiftRowsOutput[53]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_54_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, ShiftRowsOutput[54]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_55_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, ShiftRowsOutput[55]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_56_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, ShiftRowsOutput[56]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_57_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, ShiftRowsOutput[57]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_58_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, ShiftRowsOutput[58]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_59_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, ShiftRowsOutput[59]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_60_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, ShiftRowsOutput[60]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_61_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, ShiftRowsOutput[61]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_62_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, ShiftRowsOutput[62]}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_63_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, ShiftRowsOutput[63]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_64_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .a ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, ShiftRowsOutput[64]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_65_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, ShiftRowsOutput[65]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_66_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, ShiftRowsOutput[66]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_67_U1 ( .s (MuxRound_n18), .b ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, ShiftRowsOutput[67]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_68_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .a ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, ShiftRowsOutput[68]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_69_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .a ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, ShiftRowsOutput[69]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_70_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .a ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, ShiftRowsOutput[70]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_71_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .a ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, ShiftRowsOutput[71]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_72_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .a ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, ShiftRowsOutput[72]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_73_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, ShiftRowsOutput[73]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_74_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .a ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, ShiftRowsOutput[74]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_75_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, ShiftRowsOutput[75]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_76_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .a ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, ShiftRowsOutput[76]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_77_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .a ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, ShiftRowsOutput[77]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_78_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .a ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, ShiftRowsOutput[78]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_79_U1 ( .s (MuxRound_n17), .b ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, ShiftRowsOutput[79]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_80_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .a ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, ShiftRowsOutput[80]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_81_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .a ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, ShiftRowsOutput[81]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_82_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .a ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, ShiftRowsOutput[82]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_83_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .a ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, ShiftRowsOutput[83]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_84_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .a ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, ShiftRowsOutput[84]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_85_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .a ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, ShiftRowsOutput[85]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_86_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .a ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, ShiftRowsOutput[86]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_87_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .a ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, ShiftRowsOutput[87]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_88_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, ShiftRowsOutput[88]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_89_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, ShiftRowsOutput[89]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_90_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, ShiftRowsOutput[90]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_91_U1 ( .s (MuxRound_n16), .b ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, ShiftRowsOutput[91]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_92_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, ShiftRowsOutput[92]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_93_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, ShiftRowsOutput[93]}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_94_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, ShiftRowsOutput[94]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_95_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, ShiftRowsOutput[95]}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_96_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .a ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, ShiftRowsOutput[96]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_97_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, ShiftRowsOutput[97]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_98_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .a ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, ShiftRowsOutput[98]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_99_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .a ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, ShiftRowsOutput[99]}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_100_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .a ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, ShiftRowsOutput[100]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_101_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .a ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, ShiftRowsOutput[101]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_102_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .a ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, ShiftRowsOutput[102]}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_103_U1 ( .s (MuxRound_n15), .b ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .a ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, ShiftRowsOutput[103]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_104_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .a ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, ShiftRowsOutput[104]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_105_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .a ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, ShiftRowsOutput[105]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_106_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .a ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, ShiftRowsOutput[106]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_107_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .a ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, ShiftRowsOutput[107]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_108_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .a ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, ShiftRowsOutput[108]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_109_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .a ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, ShiftRowsOutput[109]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_110_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .a ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, ShiftRowsOutput[110]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_111_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .a ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, ShiftRowsOutput[111]}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_112_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .a ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, ShiftRowsOutput[112]}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_113_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .a ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, ShiftRowsOutput[113]}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_114_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, ShiftRowsOutput[114]}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_115_U1 ( .s (MuxRound_n14), .b ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .a ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, ShiftRowsOutput[115]}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_116_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .a ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, ShiftRowsOutput[116]}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_117_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .a ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, ShiftRowsOutput[117]}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_118_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .a ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, ShiftRowsOutput[118]}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_119_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .a ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, ShiftRowsOutput[119]}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_120_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, ShiftRowsOutput[120]}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_121_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, ShiftRowsOutput[121]}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_122_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, ShiftRowsOutput[122]}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_123_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, ShiftRowsOutput[123]}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_124_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, ShiftRowsOutput[124]}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_125_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, ShiftRowsOutput[125]}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_126_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, ShiftRowsOutput[126]}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_127_U1 ( .s (MuxRound_n13), .b ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, ShiftRowsOutput[127]}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, RoundOutput[127]}) ) ;
    INV_X1 MuxKeyExpansion_U8 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n14) ) ;
    INV_X1 MuxKeyExpansion_U7 ( .A (AKSRnotDone), .ZN (MuxKeyExpansion_n21) ) ;
    INV_X1 MuxKeyExpansion_U6 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n16) ) ;
    INV_X1 MuxKeyExpansion_U5 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n17) ) ;
    INV_X1 MuxKeyExpansion_U4 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n18) ) ;
    INV_X1 MuxKeyExpansion_U3 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n19) ) ;
    INV_X1 MuxKeyExpansion_U2 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n20) ) ;
    INV_X1 MuxKeyExpansion_U1 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n15) ) ;
    NOR2_X1 RoundCounterIns_U11 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_n45) ) ;
    XNOR2_X1 RoundCounterIns_U10 ( .A (RoundCounter[0]), .B (AKSRnotDone), .ZN (RoundCounterIns_n10) ) ;
    NOR2_X1 RoundCounterIns_U9 ( .A1 (reset), .A2 (RoundCounterIns_n9), .ZN (RoundCounterIns_n44) ) ;
    XOR2_X1 RoundCounterIns_U8 ( .A (RoundCounter[1]), .B (RoundCounterIns_n8), .Z (RoundCounterIns_n9) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (reset), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n42) ) ;
    XOR2_X1 RoundCounterIns_U6 ( .A (RoundCounter[3]), .B (RoundCounterIns_n6), .Z (RoundCounterIns_n7) ) ;
    NAND2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounter[2]), .ZN (RoundCounterIns_n6) ) ;
    NOR2_X1 RoundCounterIns_U4 ( .A1 (reset), .A2 (RoundCounterIns_n4), .ZN (RoundCounterIns_n1) ) ;
    XNOR2_X1 RoundCounterIns_U3 ( .A (RoundCounter[2]), .B (RoundCounterIns_n5), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (RoundCounterIns_n2), .A2 (RoundCounterIns_n8), .ZN (RoundCounterIns_n5) ) ;
    NAND2_X1 RoundCounterIns_U1 ( .A1 (AKSRnotDone), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_n8) ) ;
    INV_X1 RoundCounterIns_count_reg_1__U1 ( .A (RoundCounter[1]), .ZN (RoundCounterIns_n2) ) ;
    NOR2_X1 InRoundCounterIns_U13 ( .A1 (reset), .A2 (InRoundCounterIns_n12), .ZN (InRoundCounterIns_n41) ) ;
    XOR2_X1 InRoundCounterIns_U12 ( .A (InRoundCounter[0]), .B (InRoundCounterIns_n11), .Z (InRoundCounterIns_n12) ) ;
    NAND2_X1 InRoundCounterIns_U11 ( .A1 (InRoundCounterIns_n10), .A2 (1'b1), .ZN (InRoundCounterIns_n11) ) ;
    NAND2_X1 InRoundCounterIns_U10 ( .A1 (InRoundCounterIns_n9), .A2 (InRoundCounter[2]), .ZN (InRoundCounterIns_n10) ) ;
    NAND2_X1 InRoundCounterIns_U9 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (InRoundCounterIns_n9) ) ;
    NOR2_X1 InRoundCounterIns_U8 ( .A1 (reset), .A2 (InRoundCounterIns_n8), .ZN (InRoundCounterIns_n40) ) ;
    MUX2_X1 InRoundCounterIns_U7 ( .S (InRoundCounter[1]), .A (InRoundCounterIns_n7), .B (InRoundCounterIns_n5), .Z (InRoundCounterIns_n8) ) ;
    NOR2_X1 InRoundCounterIns_U6 ( .A1 (reset), .A2 (InRoundCounterIns_n4), .ZN (InRoundCounterIns_n39) ) ;
    NOR2_X1 InRoundCounterIns_U5 ( .A1 (InRoundCounterIns_n3), .A2 (InRoundCounterIns_n2), .ZN (InRoundCounterIns_n4) ) ;
    NOR2_X1 InRoundCounterIns_U4 ( .A1 (InRoundCounterIns_n1), .A2 (InRoundCounterIns_n7), .ZN (InRoundCounterIns_n2) ) ;
    NAND2_X1 InRoundCounterIns_U3 ( .A1 (InRoundCounterIns_n5), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n7) ) ;
    AND2_X1 InRoundCounterIns_U2 ( .A1 (InRoundCounter[0]), .A2 (1'b1), .ZN (InRoundCounterIns_n5) ) ;
    NOR2_X1 InRoundCounterIns_U1 ( .A1 (1'b1), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n3) ) ;
    INV_X1 InRoundCounterIns_count_reg_1__U1 ( .A (InRoundCounter[1]), .ZN (InRoundCounterIns_n1) ) ;
    INV_X1 InRoundCounterIns_count_reg_2__U1 ( .A (InRoundCounter[2]), .ZN (InRoundCounterIns_n6) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_7100, new_AGEMA_signal_7099, new_AGEMA_signal_7098}), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, SubBytesIns_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, SubBytesInput[0]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_4003, new_AGEMA_signal_4002, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_7103, new_AGEMA_signal_7102, new_AGEMA_signal_7101}), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_4067, new_AGEMA_signal_4066, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_4003, new_AGEMA_signal_4002, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_7106, new_AGEMA_signal_7105, new_AGEMA_signal_7104}), .c ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_4075, new_AGEMA_signal_4074, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_4067, new_AGEMA_signal_4066, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_4075, new_AGEMA_signal_4074, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_7109, new_AGEMA_signal_7108, new_AGEMA_signal_7107}), .c ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_7112, new_AGEMA_signal_7111, new_AGEMA_signal_7110}), .b ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, SubBytesIns_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, SubBytesInput[8]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_7115, new_AGEMA_signal_7114, new_AGEMA_signal_7113}), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_7118, new_AGEMA_signal_7117, new_AGEMA_signal_7116}), .c ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_7121, new_AGEMA_signal_7120, new_AGEMA_signal_7119}), .c ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_7124, new_AGEMA_signal_7123, new_AGEMA_signal_7122}), .b ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, SubBytesIns_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, SubBytesInput[16]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_4039, new_AGEMA_signal_4038, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_7127, new_AGEMA_signal_7126, new_AGEMA_signal_7125}), .b ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_3967, new_AGEMA_signal_3966, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_3967, new_AGEMA_signal_3966, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_4039, new_AGEMA_signal_4038, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_7130, new_AGEMA_signal_7129, new_AGEMA_signal_7128}), .c ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_7133, new_AGEMA_signal_7132, new_AGEMA_signal_7131}), .c ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_7136, new_AGEMA_signal_7135, new_AGEMA_signal_7134}), .b ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, SubBytesIns_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, SubBytesInput[24]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_7139, new_AGEMA_signal_7138, new_AGEMA_signal_7137}), .b ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_7142, new_AGEMA_signal_7141, new_AGEMA_signal_7140}), .c ({new_AGEMA_signal_4103, new_AGEMA_signal_4102, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_4103, new_AGEMA_signal_4102, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_7145, new_AGEMA_signal_7144, new_AGEMA_signal_7143}), .c ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2061 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_7098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_3894), .Q (new_AGEMA_signal_7099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_3895), .Q (new_AGEMA_signal_7100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2064 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_7101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_7102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_3903), .Q (new_AGEMA_signal_7103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2067 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_7104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_7105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_3995), .Q (new_AGEMA_signal_7106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2070 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_7107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_7108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_3997), .Q (new_AGEMA_signal_7109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2073 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_7110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_7111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_3921), .Q (new_AGEMA_signal_7112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2076 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_7113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_7114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_3929), .Q (new_AGEMA_signal_7115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2079 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_7116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_7117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_4013), .Q (new_AGEMA_signal_7118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2082 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_7119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_4014), .Q (new_AGEMA_signal_7120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_7121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2085 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_7122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_7123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_3947), .Q (new_AGEMA_signal_7124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2088 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_7125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_3954), .Q (new_AGEMA_signal_7126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_3955), .Q (new_AGEMA_signal_7127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2091 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_7128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_7129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_7130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2094 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_7131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_4032), .Q (new_AGEMA_signal_7132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_7133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2097 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_7134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_7135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_3973), .Q (new_AGEMA_signal_7136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2100 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_7137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_7138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_3981), .Q (new_AGEMA_signal_7139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2103 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_7140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_7141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_4049), .Q (new_AGEMA_signal_7142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2106 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_7143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_4050), .Q (new_AGEMA_signal_7144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_7145) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_7242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2209 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_7246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2213 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_7250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2217 ( .C (clk), .D (plaintext_s2[0]), .Q (new_AGEMA_signal_7254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2221 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_7258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2225 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_7262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2229 ( .C (clk), .D (plaintext_s2[1]), .Q (new_AGEMA_signal_7266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2233 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_7270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2237 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_7274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2241 ( .C (clk), .D (plaintext_s2[2]), .Q (new_AGEMA_signal_7278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2245 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_7282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2249 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_7286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2253 ( .C (clk), .D (plaintext_s2[3]), .Q (new_AGEMA_signal_7290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2257 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_7294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2261 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_7298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2265 ( .C (clk), .D (plaintext_s2[4]), .Q (new_AGEMA_signal_7302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2269 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_7306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2273 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_7310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2277 ( .C (clk), .D (plaintext_s2[5]), .Q (new_AGEMA_signal_7314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2281 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_7318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2285 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_7322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2289 ( .C (clk), .D (plaintext_s2[6]), .Q (new_AGEMA_signal_7326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2293 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_7330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2297 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_7334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2301 ( .C (clk), .D (plaintext_s2[7]), .Q (new_AGEMA_signal_7338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2305 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_7342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2309 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_7346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2313 ( .C (clk), .D (plaintext_s2[8]), .Q (new_AGEMA_signal_7350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2317 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_7354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2321 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_7358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2325 ( .C (clk), .D (plaintext_s2[9]), .Q (new_AGEMA_signal_7362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2329 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_7366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2333 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_7370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2337 ( .C (clk), .D (plaintext_s2[10]), .Q (new_AGEMA_signal_7374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2341 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_7378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2345 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_7382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2349 ( .C (clk), .D (plaintext_s2[11]), .Q (new_AGEMA_signal_7386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2353 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_7390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2357 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_7394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2361 ( .C (clk), .D (plaintext_s2[12]), .Q (new_AGEMA_signal_7398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2365 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_7402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2369 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_7406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2373 ( .C (clk), .D (plaintext_s2[13]), .Q (new_AGEMA_signal_7410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2377 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_7414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2381 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_7418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2385 ( .C (clk), .D (plaintext_s2[14]), .Q (new_AGEMA_signal_7422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2389 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_7426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2393 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_7430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2397 ( .C (clk), .D (plaintext_s2[15]), .Q (new_AGEMA_signal_7434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2401 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_7438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2405 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_7442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2409 ( .C (clk), .D (plaintext_s2[16]), .Q (new_AGEMA_signal_7446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2413 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_7450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2417 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_7454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2421 ( .C (clk), .D (plaintext_s2[17]), .Q (new_AGEMA_signal_7458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2425 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_7462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2429 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_7466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2433 ( .C (clk), .D (plaintext_s2[18]), .Q (new_AGEMA_signal_7470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2437 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_7474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2441 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_7478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2445 ( .C (clk), .D (plaintext_s2[19]), .Q (new_AGEMA_signal_7482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2449 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_7486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2453 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_7490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2457 ( .C (clk), .D (plaintext_s2[20]), .Q (new_AGEMA_signal_7494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2461 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_7498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2465 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_7502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2469 ( .C (clk), .D (plaintext_s2[21]), .Q (new_AGEMA_signal_7506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2473 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_7510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2477 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_7514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2481 ( .C (clk), .D (plaintext_s2[22]), .Q (new_AGEMA_signal_7518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2485 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_7522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2489 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_7526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2493 ( .C (clk), .D (plaintext_s2[23]), .Q (new_AGEMA_signal_7530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2497 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_7534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2501 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_7538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2505 ( .C (clk), .D (plaintext_s2[24]), .Q (new_AGEMA_signal_7542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2509 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_7546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2513 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_7550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2517 ( .C (clk), .D (plaintext_s2[25]), .Q (new_AGEMA_signal_7554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2521 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_7558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2525 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_7562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2529 ( .C (clk), .D (plaintext_s2[26]), .Q (new_AGEMA_signal_7566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2533 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_7570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2537 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_7574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2541 ( .C (clk), .D (plaintext_s2[27]), .Q (new_AGEMA_signal_7578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2545 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_7582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2549 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_7586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2553 ( .C (clk), .D (plaintext_s2[28]), .Q (new_AGEMA_signal_7590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2557 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_7594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2561 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_7598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2565 ( .C (clk), .D (plaintext_s2[29]), .Q (new_AGEMA_signal_7602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2569 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_7606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2573 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_7610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2577 ( .C (clk), .D (plaintext_s2[30]), .Q (new_AGEMA_signal_7614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2581 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_7618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2585 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_7622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2589 ( .C (clk), .D (plaintext_s2[31]), .Q (new_AGEMA_signal_7626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2593 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_7630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_3826), .Q (new_AGEMA_signal_7633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_3827), .Q (new_AGEMA_signal_7636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2602 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_7639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_3890), .Q (new_AGEMA_signal_7642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_3891), .Q (new_AGEMA_signal_7645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2611 ( .C (clk), .D (SubBytesInput[0]), .Q (new_AGEMA_signal_7648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_7651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_3109), .Q (new_AGEMA_signal_7654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2620 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_7657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_3834), .Q (new_AGEMA_signal_7660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_3835), .Q (new_AGEMA_signal_7663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2629 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_7666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_3828), .Q (new_AGEMA_signal_7669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_3829), .Q (new_AGEMA_signal_7672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2638 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_7675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_7678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_3897), .Q (new_AGEMA_signal_7681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2647 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_7684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_3832), .Q (new_AGEMA_signal_7687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_3833), .Q (new_AGEMA_signal_7690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2656 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_7693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_7696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_3841), .Q (new_AGEMA_signal_7699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2665 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_7702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_3892), .Q (new_AGEMA_signal_7705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_3893), .Q (new_AGEMA_signal_7708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2674 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_7711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_3830), .Q (new_AGEMA_signal_7714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_3831), .Q (new_AGEMA_signal_7717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2683 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_7720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_7723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_3901), .Q (new_AGEMA_signal_7726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2692 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_7729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_7732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_3837), .Q (new_AGEMA_signal_7735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2701 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_7738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_7741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_7744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2710 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_7747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_7750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_3839), .Q (new_AGEMA_signal_7753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2719 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_7756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_3898), .Q (new_AGEMA_signal_7759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_3899), .Q (new_AGEMA_signal_7762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2728 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_7765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_3746), .Q (new_AGEMA_signal_7768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_7771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2737 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_7774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_7777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_7780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2746 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_7783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_3748), .Q (new_AGEMA_signal_7786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_3749), .Q (new_AGEMA_signal_7789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2755 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_7792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_3842), .Q (new_AGEMA_signal_7795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_3843), .Q (new_AGEMA_signal_7798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2764 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_7801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_7804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_3917), .Q (new_AGEMA_signal_7807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2773 ( .C (clk), .D (SubBytesInput[8]), .Q (new_AGEMA_signal_7810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_3106), .Q (new_AGEMA_signal_7813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_3107), .Q (new_AGEMA_signal_7816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2782 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_7819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_3850), .Q (new_AGEMA_signal_7822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_3851), .Q (new_AGEMA_signal_7825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2791 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_7828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_3844), .Q (new_AGEMA_signal_7831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_3845), .Q (new_AGEMA_signal_7834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2800 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_7837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_3922), .Q (new_AGEMA_signal_7840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_3923), .Q (new_AGEMA_signal_7843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2809 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_7846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_3848), .Q (new_AGEMA_signal_7849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_3849), .Q (new_AGEMA_signal_7852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2818 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_7855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_3856), .Q (new_AGEMA_signal_7858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_3857), .Q (new_AGEMA_signal_7861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2827 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_7864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_7867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_3919), .Q (new_AGEMA_signal_7870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2836 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_7873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_3846), .Q (new_AGEMA_signal_7876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_3847), .Q (new_AGEMA_signal_7879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2845 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_7882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_7885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_3927), .Q (new_AGEMA_signal_7888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2854 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_7891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_7894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_3853), .Q (new_AGEMA_signal_7897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2863 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_7900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_3770), .Q (new_AGEMA_signal_7903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_3771), .Q (new_AGEMA_signal_7906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2872 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_7909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_7912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_3855), .Q (new_AGEMA_signal_7915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2881 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_7918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_7921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_3925), .Q (new_AGEMA_signal_7924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2890 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_7927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_3766), .Q (new_AGEMA_signal_7930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_3767), .Q (new_AGEMA_signal_7933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2899 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_7936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_3772), .Q (new_AGEMA_signal_7939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_3773), .Q (new_AGEMA_signal_7942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2908 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_7945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_7948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_7951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2917 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_7954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_3858), .Q (new_AGEMA_signal_7957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_3859), .Q (new_AGEMA_signal_7960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2926 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_7963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_7966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_7969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2935 ( .C (clk), .D (SubBytesInput[16]), .Q (new_AGEMA_signal_7972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_3138), .Q (new_AGEMA_signal_7975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_3139), .Q (new_AGEMA_signal_7978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2944 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_7981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_3866), .Q (new_AGEMA_signal_7984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_3867), .Q (new_AGEMA_signal_7987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2953 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_7990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_7993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_3861), .Q (new_AGEMA_signal_7996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2962 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_7999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_8002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_3949), .Q (new_AGEMA_signal_8005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2971 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_8008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_8011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_3865), .Q (new_AGEMA_signal_8014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2980 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_8017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_3872), .Q (new_AGEMA_signal_8020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_3873), .Q (new_AGEMA_signal_8023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2989 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_8026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_8029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_3945), .Q (new_AGEMA_signal_8032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2998 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_8035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_8038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_3863), .Q (new_AGEMA_signal_8041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3007 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_8044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_8047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_3953), .Q (new_AGEMA_signal_8050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3016 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_8053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_3868), .Q (new_AGEMA_signal_8056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_3869), .Q (new_AGEMA_signal_8059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3025 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_8062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_3790), .Q (new_AGEMA_signal_8065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_3791), .Q (new_AGEMA_signal_8068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3034 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_8071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_3870), .Q (new_AGEMA_signal_8074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_3871), .Q (new_AGEMA_signal_8077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3043 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_8080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_8083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_3951), .Q (new_AGEMA_signal_8086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3052 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_8089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_3786), .Q (new_AGEMA_signal_8092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_3787), .Q (new_AGEMA_signal_8095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3061 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_8098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_3792), .Q (new_AGEMA_signal_8101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_3793), .Q (new_AGEMA_signal_8104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3070 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_8107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_3788), .Q (new_AGEMA_signal_8110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_3789), .Q (new_AGEMA_signal_8113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3079 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_8116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_3874), .Q (new_AGEMA_signal_8119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_3875), .Q (new_AGEMA_signal_8122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3088 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_8125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_8128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_3969), .Q (new_AGEMA_signal_8131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3097 ( .C (clk), .D (SubBytesInput[24]), .Q (new_AGEMA_signal_8134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_3154), .Q (new_AGEMA_signal_8137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_3155), .Q (new_AGEMA_signal_8140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3106 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_8143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_3882), .Q (new_AGEMA_signal_8146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_3883), .Q (new_AGEMA_signal_8149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3115 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_8152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_3876), .Q (new_AGEMA_signal_8155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_3877), .Q (new_AGEMA_signal_8158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3124 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_8161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_8164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_3975), .Q (new_AGEMA_signal_8167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3133 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_8170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_3880), .Q (new_AGEMA_signal_8173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_3881), .Q (new_AGEMA_signal_8176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3142 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_8179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_8182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_3889), .Q (new_AGEMA_signal_8185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3151 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_8188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_3970), .Q (new_AGEMA_signal_8191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_3971), .Q (new_AGEMA_signal_8194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3160 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_8197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_8200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_3879), .Q (new_AGEMA_signal_8203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3169 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_8206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_3978), .Q (new_AGEMA_signal_8209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_8212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3178 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_8215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_8218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_3885), .Q (new_AGEMA_signal_8221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3187 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_8224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_3810), .Q (new_AGEMA_signal_8227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_3811), .Q (new_AGEMA_signal_8230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3196 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_8233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_8236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_3887), .Q (new_AGEMA_signal_8239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3205 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_8242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_8245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_3977), .Q (new_AGEMA_signal_8248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3214 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_8251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_3806), .Q (new_AGEMA_signal_8254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_3807), .Q (new_AGEMA_signal_8257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3223 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_8260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_8263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_3813), .Q (new_AGEMA_signal_8266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3232 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_8269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_3808), .Q (new_AGEMA_signal_8272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_3809), .Q (new_AGEMA_signal_8275) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (MuxMCOut_n5), .Q (new_AGEMA_signal_8278) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (LastRoundorDone), .Q (new_AGEMA_signal_8282) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (MuxMCOut_n4), .Q (new_AGEMA_signal_8286) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (AKSRnotDone), .Q (new_AGEMA_signal_8290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3257 ( .C (clk), .D (ShiftRowsOutput[0]), .Q (new_AGEMA_signal_8294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_8298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_2661), .Q (new_AGEMA_signal_8302) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (MuxRound_n13), .Q (new_AGEMA_signal_8306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3273 ( .C (clk), .D (ShiftRowsOutput[1]), .Q (new_AGEMA_signal_8310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_8314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_2667), .Q (new_AGEMA_signal_8318) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (MuxRound_n14), .Q (new_AGEMA_signal_8322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3289 ( .C (clk), .D (ShiftRowsOutput[2]), .Q (new_AGEMA_signal_8326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_8330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_2673), .Q (new_AGEMA_signal_8334) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (MuxRound_n15), .Q (new_AGEMA_signal_8338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3305 ( .C (clk), .D (ShiftRowsOutput[3]), .Q (new_AGEMA_signal_8342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_2678), .Q (new_AGEMA_signal_8346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_2679), .Q (new_AGEMA_signal_8350) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (MuxRound_n16), .Q (new_AGEMA_signal_8354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3321 ( .C (clk), .D (ShiftRowsOutput[4]), .Q (new_AGEMA_signal_8358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_8362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_2685), .Q (new_AGEMA_signal_8366) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (MuxRound_n17), .Q (new_AGEMA_signal_8370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3337 ( .C (clk), .D (ShiftRowsOutput[5]), .Q (new_AGEMA_signal_8374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_2690), .Q (new_AGEMA_signal_8378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_2691), .Q (new_AGEMA_signal_8382) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (MuxRound_n18), .Q (new_AGEMA_signal_8386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3353 ( .C (clk), .D (ShiftRowsOutput[6]), .Q (new_AGEMA_signal_8390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_2696), .Q (new_AGEMA_signal_8394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_2697), .Q (new_AGEMA_signal_8398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3365 ( .C (clk), .D (ShiftRowsOutput[7]), .Q (new_AGEMA_signal_8402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_8406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_2703), .Q (new_AGEMA_signal_8410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3377 ( .C (clk), .D (ShiftRowsOutput[8]), .Q (new_AGEMA_signal_8414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_2924), .Q (new_AGEMA_signal_8418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_2925), .Q (new_AGEMA_signal_8422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3389 ( .C (clk), .D (ShiftRowsOutput[9]), .Q (new_AGEMA_signal_8426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_2930), .Q (new_AGEMA_signal_8430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_2931), .Q (new_AGEMA_signal_8434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3401 ( .C (clk), .D (ShiftRowsOutput[10]), .Q (new_AGEMA_signal_8438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_2936), .Q (new_AGEMA_signal_8442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_2937), .Q (new_AGEMA_signal_8446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3413 ( .C (clk), .D (ShiftRowsOutput[11]), .Q (new_AGEMA_signal_8450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_2942), .Q (new_AGEMA_signal_8454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_2943), .Q (new_AGEMA_signal_8458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3425 ( .C (clk), .D (ShiftRowsOutput[12]), .Q (new_AGEMA_signal_8462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_2948), .Q (new_AGEMA_signal_8466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_2949), .Q (new_AGEMA_signal_8470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3437 ( .C (clk), .D (ShiftRowsOutput[13]), .Q (new_AGEMA_signal_8474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_2954), .Q (new_AGEMA_signal_8478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_2955), .Q (new_AGEMA_signal_8482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3449 ( .C (clk), .D (ShiftRowsOutput[14]), .Q (new_AGEMA_signal_8486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_2960), .Q (new_AGEMA_signal_8490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_2961), .Q (new_AGEMA_signal_8494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3461 ( .C (clk), .D (ShiftRowsOutput[15]), .Q (new_AGEMA_signal_8498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_2966), .Q (new_AGEMA_signal_8502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_2967), .Q (new_AGEMA_signal_8506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3473 ( .C (clk), .D (ShiftRowsOutput[16]), .Q (new_AGEMA_signal_8510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_2426), .Q (new_AGEMA_signal_8514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_2427), .Q (new_AGEMA_signal_8518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3485 ( .C (clk), .D (ShiftRowsOutput[17]), .Q (new_AGEMA_signal_8522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_2432), .Q (new_AGEMA_signal_8526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_2433), .Q (new_AGEMA_signal_8530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3497 ( .C (clk), .D (ShiftRowsOutput[18]), .Q (new_AGEMA_signal_8534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3501 ( .C (clk), .D (new_AGEMA_signal_2438), .Q (new_AGEMA_signal_8538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_2439), .Q (new_AGEMA_signal_8542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3509 ( .C (clk), .D (ShiftRowsOutput[19]), .Q (new_AGEMA_signal_8546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_2444), .Q (new_AGEMA_signal_8550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_2445), .Q (new_AGEMA_signal_8554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3521 ( .C (clk), .D (ShiftRowsOutput[20]), .Q (new_AGEMA_signal_8558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_2450), .Q (new_AGEMA_signal_8562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_2451), .Q (new_AGEMA_signal_8566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3533 ( .C (clk), .D (ShiftRowsOutput[21]), .Q (new_AGEMA_signal_8570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3537 ( .C (clk), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_8574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_2457), .Q (new_AGEMA_signal_8578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3545 ( .C (clk), .D (ShiftRowsOutput[22]), .Q (new_AGEMA_signal_8582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_2462), .Q (new_AGEMA_signal_8586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_2463), .Q (new_AGEMA_signal_8590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3557 ( .C (clk), .D (ShiftRowsOutput[23]), .Q (new_AGEMA_signal_8594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_8598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_2469), .Q (new_AGEMA_signal_8602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3569 ( .C (clk), .D (ShiftRowsOutput[24]), .Q (new_AGEMA_signal_8606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3573 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_8610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_2607), .Q (new_AGEMA_signal_8614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3581 ( .C (clk), .D (ShiftRowsOutput[25]), .Q (new_AGEMA_signal_8618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3585 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_8622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_2613), .Q (new_AGEMA_signal_8626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3593 ( .C (clk), .D (ShiftRowsOutput[26]), .Q (new_AGEMA_signal_8630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_8634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_2619), .Q (new_AGEMA_signal_8638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3605 ( .C (clk), .D (ShiftRowsOutput[27]), .Q (new_AGEMA_signal_8642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3609 ( .C (clk), .D (new_AGEMA_signal_2624), .Q (new_AGEMA_signal_8646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_2625), .Q (new_AGEMA_signal_8650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3617 ( .C (clk), .D (ShiftRowsOutput[28]), .Q (new_AGEMA_signal_8654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3621 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_8658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_2631), .Q (new_AGEMA_signal_8662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3629 ( .C (clk), .D (ShiftRowsOutput[29]), .Q (new_AGEMA_signal_8666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_8670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_2637), .Q (new_AGEMA_signal_8674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3641 ( .C (clk), .D (ShiftRowsOutput[30]), .Q (new_AGEMA_signal_8678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3645 ( .C (clk), .D (new_AGEMA_signal_2648), .Q (new_AGEMA_signal_8682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_2649), .Q (new_AGEMA_signal_8686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3653 ( .C (clk), .D (ShiftRowsOutput[31]), .Q (new_AGEMA_signal_8690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_8694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_2655), .Q (new_AGEMA_signal_8698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3665 ( .C (clk), .D (key_s0[0]), .Q (new_AGEMA_signal_8702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3669 ( .C (clk), .D (key_s1[0]), .Q (new_AGEMA_signal_8706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3673 ( .C (clk), .D (key_s2[0]), .Q (new_AGEMA_signal_8710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3677 ( .C (clk), .D (key_s0[1]), .Q (new_AGEMA_signal_8714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3681 ( .C (clk), .D (key_s1[1]), .Q (new_AGEMA_signal_8718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3685 ( .C (clk), .D (key_s2[1]), .Q (new_AGEMA_signal_8722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3689 ( .C (clk), .D (key_s0[2]), .Q (new_AGEMA_signal_8726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3693 ( .C (clk), .D (key_s1[2]), .Q (new_AGEMA_signal_8730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3697 ( .C (clk), .D (key_s2[2]), .Q (new_AGEMA_signal_8734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3701 ( .C (clk), .D (key_s0[3]), .Q (new_AGEMA_signal_8738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3705 ( .C (clk), .D (key_s1[3]), .Q (new_AGEMA_signal_8742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3709 ( .C (clk), .D (key_s2[3]), .Q (new_AGEMA_signal_8746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3713 ( .C (clk), .D (key_s0[4]), .Q (new_AGEMA_signal_8750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3717 ( .C (clk), .D (key_s1[4]), .Q (new_AGEMA_signal_8754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3721 ( .C (clk), .D (key_s2[4]), .Q (new_AGEMA_signal_8758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3725 ( .C (clk), .D (key_s0[5]), .Q (new_AGEMA_signal_8762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3729 ( .C (clk), .D (key_s1[5]), .Q (new_AGEMA_signal_8766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3733 ( .C (clk), .D (key_s2[5]), .Q (new_AGEMA_signal_8770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3737 ( .C (clk), .D (key_s0[6]), .Q (new_AGEMA_signal_8774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3741 ( .C (clk), .D (key_s1[6]), .Q (new_AGEMA_signal_8778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3745 ( .C (clk), .D (key_s2[6]), .Q (new_AGEMA_signal_8782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3749 ( .C (clk), .D (key_s0[7]), .Q (new_AGEMA_signal_8786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3753 ( .C (clk), .D (key_s1[7]), .Q (new_AGEMA_signal_8790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3757 ( .C (clk), .D (key_s2[7]), .Q (new_AGEMA_signal_8794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3761 ( .C (clk), .D (key_s0[8]), .Q (new_AGEMA_signal_8798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3765 ( .C (clk), .D (key_s1[8]), .Q (new_AGEMA_signal_8802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3769 ( .C (clk), .D (key_s2[8]), .Q (new_AGEMA_signal_8806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3773 ( .C (clk), .D (key_s0[9]), .Q (new_AGEMA_signal_8810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3777 ( .C (clk), .D (key_s1[9]), .Q (new_AGEMA_signal_8814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3781 ( .C (clk), .D (key_s2[9]), .Q (new_AGEMA_signal_8818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3785 ( .C (clk), .D (key_s0[10]), .Q (new_AGEMA_signal_8822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3789 ( .C (clk), .D (key_s1[10]), .Q (new_AGEMA_signal_8826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3793 ( .C (clk), .D (key_s2[10]), .Q (new_AGEMA_signal_8830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3797 ( .C (clk), .D (key_s0[11]), .Q (new_AGEMA_signal_8834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3801 ( .C (clk), .D (key_s1[11]), .Q (new_AGEMA_signal_8838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3805 ( .C (clk), .D (key_s2[11]), .Q (new_AGEMA_signal_8842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3809 ( .C (clk), .D (key_s0[12]), .Q (new_AGEMA_signal_8846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3813 ( .C (clk), .D (key_s1[12]), .Q (new_AGEMA_signal_8850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3817 ( .C (clk), .D (key_s2[12]), .Q (new_AGEMA_signal_8854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3821 ( .C (clk), .D (key_s0[13]), .Q (new_AGEMA_signal_8858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3825 ( .C (clk), .D (key_s1[13]), .Q (new_AGEMA_signal_8862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3829 ( .C (clk), .D (key_s2[13]), .Q (new_AGEMA_signal_8866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3833 ( .C (clk), .D (key_s0[14]), .Q (new_AGEMA_signal_8870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3837 ( .C (clk), .D (key_s1[14]), .Q (new_AGEMA_signal_8874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3841 ( .C (clk), .D (key_s2[14]), .Q (new_AGEMA_signal_8878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3845 ( .C (clk), .D (key_s0[15]), .Q (new_AGEMA_signal_8882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3849 ( .C (clk), .D (key_s1[15]), .Q (new_AGEMA_signal_8886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3853 ( .C (clk), .D (key_s2[15]), .Q (new_AGEMA_signal_8890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3857 ( .C (clk), .D (key_s0[16]), .Q (new_AGEMA_signal_8894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3861 ( .C (clk), .D (key_s1[16]), .Q (new_AGEMA_signal_8898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3865 ( .C (clk), .D (key_s2[16]), .Q (new_AGEMA_signal_8902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3869 ( .C (clk), .D (key_s0[17]), .Q (new_AGEMA_signal_8906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3873 ( .C (clk), .D (key_s1[17]), .Q (new_AGEMA_signal_8910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3877 ( .C (clk), .D (key_s2[17]), .Q (new_AGEMA_signal_8914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3881 ( .C (clk), .D (key_s0[18]), .Q (new_AGEMA_signal_8918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3885 ( .C (clk), .D (key_s1[18]), .Q (new_AGEMA_signal_8922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3889 ( .C (clk), .D (key_s2[18]), .Q (new_AGEMA_signal_8926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3893 ( .C (clk), .D (key_s0[19]), .Q (new_AGEMA_signal_8930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3897 ( .C (clk), .D (key_s1[19]), .Q (new_AGEMA_signal_8934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3901 ( .C (clk), .D (key_s2[19]), .Q (new_AGEMA_signal_8938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3905 ( .C (clk), .D (key_s0[20]), .Q (new_AGEMA_signal_8942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3909 ( .C (clk), .D (key_s1[20]), .Q (new_AGEMA_signal_8946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3913 ( .C (clk), .D (key_s2[20]), .Q (new_AGEMA_signal_8950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3917 ( .C (clk), .D (key_s0[21]), .Q (new_AGEMA_signal_8954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3921 ( .C (clk), .D (key_s1[21]), .Q (new_AGEMA_signal_8958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3925 ( .C (clk), .D (key_s2[21]), .Q (new_AGEMA_signal_8962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3929 ( .C (clk), .D (key_s0[22]), .Q (new_AGEMA_signal_8966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3933 ( .C (clk), .D (key_s1[22]), .Q (new_AGEMA_signal_8970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3937 ( .C (clk), .D (key_s2[22]), .Q (new_AGEMA_signal_8974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3941 ( .C (clk), .D (key_s0[23]), .Q (new_AGEMA_signal_8978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3945 ( .C (clk), .D (key_s1[23]), .Q (new_AGEMA_signal_8982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3949 ( .C (clk), .D (key_s2[23]), .Q (new_AGEMA_signal_8986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3953 ( .C (clk), .D (key_s0[24]), .Q (new_AGEMA_signal_8990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3957 ( .C (clk), .D (key_s1[24]), .Q (new_AGEMA_signal_8994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3961 ( .C (clk), .D (key_s2[24]), .Q (new_AGEMA_signal_8998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3965 ( .C (clk), .D (key_s0[25]), .Q (new_AGEMA_signal_9002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3969 ( .C (clk), .D (key_s1[25]), .Q (new_AGEMA_signal_9006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3973 ( .C (clk), .D (key_s2[25]), .Q (new_AGEMA_signal_9010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3977 ( .C (clk), .D (key_s0[26]), .Q (new_AGEMA_signal_9014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3981 ( .C (clk), .D (key_s1[26]), .Q (new_AGEMA_signal_9018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3985 ( .C (clk), .D (key_s2[26]), .Q (new_AGEMA_signal_9022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3989 ( .C (clk), .D (key_s0[27]), .Q (new_AGEMA_signal_9026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3993 ( .C (clk), .D (key_s1[27]), .Q (new_AGEMA_signal_9030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3997 ( .C (clk), .D (key_s2[27]), .Q (new_AGEMA_signal_9034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4001 ( .C (clk), .D (key_s0[28]), .Q (new_AGEMA_signal_9038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4005 ( .C (clk), .D (key_s1[28]), .Q (new_AGEMA_signal_9042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4009 ( .C (clk), .D (key_s2[28]), .Q (new_AGEMA_signal_9046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4013 ( .C (clk), .D (key_s0[29]), .Q (new_AGEMA_signal_9050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4017 ( .C (clk), .D (key_s1[29]), .Q (new_AGEMA_signal_9054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4021 ( .C (clk), .D (key_s2[29]), .Q (new_AGEMA_signal_9058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4025 ( .C (clk), .D (key_s0[30]), .Q (new_AGEMA_signal_9062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4029 ( .C (clk), .D (key_s1[30]), .Q (new_AGEMA_signal_9066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4033 ( .C (clk), .D (key_s2[30]), .Q (new_AGEMA_signal_9070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4037 ( .C (clk), .D (key_s0[31]), .Q (new_AGEMA_signal_9074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4041 ( .C (clk), .D (key_s1[31]), .Q (new_AGEMA_signal_9078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4045 ( .C (clk), .D (key_s2[31]), .Q (new_AGEMA_signal_9082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4049 ( .C (clk), .D (key_s0[32]), .Q (new_AGEMA_signal_9086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4053 ( .C (clk), .D (key_s1[32]), .Q (new_AGEMA_signal_9090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4057 ( .C (clk), .D (key_s2[32]), .Q (new_AGEMA_signal_9094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4061 ( .C (clk), .D (key_s0[33]), .Q (new_AGEMA_signal_9098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4065 ( .C (clk), .D (key_s1[33]), .Q (new_AGEMA_signal_9102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4069 ( .C (clk), .D (key_s2[33]), .Q (new_AGEMA_signal_9106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4073 ( .C (clk), .D (key_s0[34]), .Q (new_AGEMA_signal_9110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4077 ( .C (clk), .D (key_s1[34]), .Q (new_AGEMA_signal_9114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4081 ( .C (clk), .D (key_s2[34]), .Q (new_AGEMA_signal_9118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4085 ( .C (clk), .D (key_s0[35]), .Q (new_AGEMA_signal_9122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4089 ( .C (clk), .D (key_s1[35]), .Q (new_AGEMA_signal_9126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4093 ( .C (clk), .D (key_s2[35]), .Q (new_AGEMA_signal_9130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4097 ( .C (clk), .D (key_s0[36]), .Q (new_AGEMA_signal_9134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4101 ( .C (clk), .D (key_s1[36]), .Q (new_AGEMA_signal_9138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4105 ( .C (clk), .D (key_s2[36]), .Q (new_AGEMA_signal_9142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4109 ( .C (clk), .D (key_s0[37]), .Q (new_AGEMA_signal_9146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4113 ( .C (clk), .D (key_s1[37]), .Q (new_AGEMA_signal_9150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4117 ( .C (clk), .D (key_s2[37]), .Q (new_AGEMA_signal_9154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4121 ( .C (clk), .D (key_s0[38]), .Q (new_AGEMA_signal_9158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4125 ( .C (clk), .D (key_s1[38]), .Q (new_AGEMA_signal_9162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4129 ( .C (clk), .D (key_s2[38]), .Q (new_AGEMA_signal_9166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4133 ( .C (clk), .D (key_s0[39]), .Q (new_AGEMA_signal_9170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4137 ( .C (clk), .D (key_s1[39]), .Q (new_AGEMA_signal_9174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4141 ( .C (clk), .D (key_s2[39]), .Q (new_AGEMA_signal_9178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4145 ( .C (clk), .D (key_s0[40]), .Q (new_AGEMA_signal_9182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4149 ( .C (clk), .D (key_s1[40]), .Q (new_AGEMA_signal_9186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4153 ( .C (clk), .D (key_s2[40]), .Q (new_AGEMA_signal_9190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4157 ( .C (clk), .D (key_s0[41]), .Q (new_AGEMA_signal_9194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4161 ( .C (clk), .D (key_s1[41]), .Q (new_AGEMA_signal_9198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4165 ( .C (clk), .D (key_s2[41]), .Q (new_AGEMA_signal_9202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4169 ( .C (clk), .D (key_s0[42]), .Q (new_AGEMA_signal_9206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4173 ( .C (clk), .D (key_s1[42]), .Q (new_AGEMA_signal_9210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4177 ( .C (clk), .D (key_s2[42]), .Q (new_AGEMA_signal_9214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4181 ( .C (clk), .D (key_s0[43]), .Q (new_AGEMA_signal_9218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4185 ( .C (clk), .D (key_s1[43]), .Q (new_AGEMA_signal_9222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4189 ( .C (clk), .D (key_s2[43]), .Q (new_AGEMA_signal_9226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4193 ( .C (clk), .D (key_s0[44]), .Q (new_AGEMA_signal_9230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4197 ( .C (clk), .D (key_s1[44]), .Q (new_AGEMA_signal_9234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4201 ( .C (clk), .D (key_s2[44]), .Q (new_AGEMA_signal_9238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4205 ( .C (clk), .D (key_s0[45]), .Q (new_AGEMA_signal_9242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4209 ( .C (clk), .D (key_s1[45]), .Q (new_AGEMA_signal_9246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4213 ( .C (clk), .D (key_s2[45]), .Q (new_AGEMA_signal_9250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4217 ( .C (clk), .D (key_s0[46]), .Q (new_AGEMA_signal_9254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4221 ( .C (clk), .D (key_s1[46]), .Q (new_AGEMA_signal_9258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4225 ( .C (clk), .D (key_s2[46]), .Q (new_AGEMA_signal_9262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4229 ( .C (clk), .D (key_s0[47]), .Q (new_AGEMA_signal_9266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4233 ( .C (clk), .D (key_s1[47]), .Q (new_AGEMA_signal_9270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4237 ( .C (clk), .D (key_s2[47]), .Q (new_AGEMA_signal_9274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4241 ( .C (clk), .D (key_s0[48]), .Q (new_AGEMA_signal_9278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4245 ( .C (clk), .D (key_s1[48]), .Q (new_AGEMA_signal_9282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4249 ( .C (clk), .D (key_s2[48]), .Q (new_AGEMA_signal_9286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4253 ( .C (clk), .D (key_s0[49]), .Q (new_AGEMA_signal_9290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4257 ( .C (clk), .D (key_s1[49]), .Q (new_AGEMA_signal_9294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4261 ( .C (clk), .D (key_s2[49]), .Q (new_AGEMA_signal_9298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4265 ( .C (clk), .D (key_s0[50]), .Q (new_AGEMA_signal_9302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4269 ( .C (clk), .D (key_s1[50]), .Q (new_AGEMA_signal_9306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4273 ( .C (clk), .D (key_s2[50]), .Q (new_AGEMA_signal_9310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4277 ( .C (clk), .D (key_s0[51]), .Q (new_AGEMA_signal_9314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4281 ( .C (clk), .D (key_s1[51]), .Q (new_AGEMA_signal_9318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4285 ( .C (clk), .D (key_s2[51]), .Q (new_AGEMA_signal_9322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4289 ( .C (clk), .D (key_s0[52]), .Q (new_AGEMA_signal_9326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4293 ( .C (clk), .D (key_s1[52]), .Q (new_AGEMA_signal_9330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4297 ( .C (clk), .D (key_s2[52]), .Q (new_AGEMA_signal_9334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4301 ( .C (clk), .D (key_s0[53]), .Q (new_AGEMA_signal_9338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4305 ( .C (clk), .D (key_s1[53]), .Q (new_AGEMA_signal_9342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4309 ( .C (clk), .D (key_s2[53]), .Q (new_AGEMA_signal_9346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4313 ( .C (clk), .D (key_s0[54]), .Q (new_AGEMA_signal_9350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4317 ( .C (clk), .D (key_s1[54]), .Q (new_AGEMA_signal_9354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4321 ( .C (clk), .D (key_s2[54]), .Q (new_AGEMA_signal_9358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4325 ( .C (clk), .D (key_s0[55]), .Q (new_AGEMA_signal_9362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4329 ( .C (clk), .D (key_s1[55]), .Q (new_AGEMA_signal_9366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4333 ( .C (clk), .D (key_s2[55]), .Q (new_AGEMA_signal_9370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4337 ( .C (clk), .D (key_s0[56]), .Q (new_AGEMA_signal_9374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4341 ( .C (clk), .D (key_s1[56]), .Q (new_AGEMA_signal_9378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4345 ( .C (clk), .D (key_s2[56]), .Q (new_AGEMA_signal_9382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4349 ( .C (clk), .D (key_s0[57]), .Q (new_AGEMA_signal_9386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4353 ( .C (clk), .D (key_s1[57]), .Q (new_AGEMA_signal_9390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4357 ( .C (clk), .D (key_s2[57]), .Q (new_AGEMA_signal_9394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4361 ( .C (clk), .D (key_s0[58]), .Q (new_AGEMA_signal_9398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4365 ( .C (clk), .D (key_s1[58]), .Q (new_AGEMA_signal_9402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4369 ( .C (clk), .D (key_s2[58]), .Q (new_AGEMA_signal_9406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4373 ( .C (clk), .D (key_s0[59]), .Q (new_AGEMA_signal_9410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4377 ( .C (clk), .D (key_s1[59]), .Q (new_AGEMA_signal_9414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4381 ( .C (clk), .D (key_s2[59]), .Q (new_AGEMA_signal_9418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4385 ( .C (clk), .D (key_s0[60]), .Q (new_AGEMA_signal_9422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4389 ( .C (clk), .D (key_s1[60]), .Q (new_AGEMA_signal_9426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4393 ( .C (clk), .D (key_s2[60]), .Q (new_AGEMA_signal_9430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4397 ( .C (clk), .D (key_s0[61]), .Q (new_AGEMA_signal_9434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4401 ( .C (clk), .D (key_s1[61]), .Q (new_AGEMA_signal_9438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4405 ( .C (clk), .D (key_s2[61]), .Q (new_AGEMA_signal_9442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4409 ( .C (clk), .D (key_s0[62]), .Q (new_AGEMA_signal_9446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4413 ( .C (clk), .D (key_s1[62]), .Q (new_AGEMA_signal_9450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4417 ( .C (clk), .D (key_s2[62]), .Q (new_AGEMA_signal_9454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4421 ( .C (clk), .D (key_s0[63]), .Q (new_AGEMA_signal_9458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4425 ( .C (clk), .D (key_s1[63]), .Q (new_AGEMA_signal_9462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4429 ( .C (clk), .D (key_s2[63]), .Q (new_AGEMA_signal_9466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4433 ( .C (clk), .D (key_s0[64]), .Q (new_AGEMA_signal_9470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4437 ( .C (clk), .D (key_s1[64]), .Q (new_AGEMA_signal_9474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4441 ( .C (clk), .D (key_s2[64]), .Q (new_AGEMA_signal_9478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4445 ( .C (clk), .D (key_s0[65]), .Q (new_AGEMA_signal_9482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4449 ( .C (clk), .D (key_s1[65]), .Q (new_AGEMA_signal_9486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4453 ( .C (clk), .D (key_s2[65]), .Q (new_AGEMA_signal_9490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4457 ( .C (clk), .D (key_s0[66]), .Q (new_AGEMA_signal_9494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4461 ( .C (clk), .D (key_s1[66]), .Q (new_AGEMA_signal_9498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4465 ( .C (clk), .D (key_s2[66]), .Q (new_AGEMA_signal_9502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4469 ( .C (clk), .D (key_s0[67]), .Q (new_AGEMA_signal_9506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4473 ( .C (clk), .D (key_s1[67]), .Q (new_AGEMA_signal_9510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4477 ( .C (clk), .D (key_s2[67]), .Q (new_AGEMA_signal_9514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4481 ( .C (clk), .D (key_s0[68]), .Q (new_AGEMA_signal_9518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4485 ( .C (clk), .D (key_s1[68]), .Q (new_AGEMA_signal_9522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4489 ( .C (clk), .D (key_s2[68]), .Q (new_AGEMA_signal_9526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4493 ( .C (clk), .D (key_s0[69]), .Q (new_AGEMA_signal_9530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4497 ( .C (clk), .D (key_s1[69]), .Q (new_AGEMA_signal_9534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4501 ( .C (clk), .D (key_s2[69]), .Q (new_AGEMA_signal_9538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4505 ( .C (clk), .D (key_s0[70]), .Q (new_AGEMA_signal_9542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4509 ( .C (clk), .D (key_s1[70]), .Q (new_AGEMA_signal_9546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4513 ( .C (clk), .D (key_s2[70]), .Q (new_AGEMA_signal_9550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4517 ( .C (clk), .D (key_s0[71]), .Q (new_AGEMA_signal_9554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4521 ( .C (clk), .D (key_s1[71]), .Q (new_AGEMA_signal_9558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4525 ( .C (clk), .D (key_s2[71]), .Q (new_AGEMA_signal_9562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4529 ( .C (clk), .D (key_s0[72]), .Q (new_AGEMA_signal_9566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4533 ( .C (clk), .D (key_s1[72]), .Q (new_AGEMA_signal_9570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4537 ( .C (clk), .D (key_s2[72]), .Q (new_AGEMA_signal_9574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4541 ( .C (clk), .D (key_s0[73]), .Q (new_AGEMA_signal_9578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4545 ( .C (clk), .D (key_s1[73]), .Q (new_AGEMA_signal_9582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4549 ( .C (clk), .D (key_s2[73]), .Q (new_AGEMA_signal_9586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4553 ( .C (clk), .D (key_s0[74]), .Q (new_AGEMA_signal_9590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4557 ( .C (clk), .D (key_s1[74]), .Q (new_AGEMA_signal_9594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4561 ( .C (clk), .D (key_s2[74]), .Q (new_AGEMA_signal_9598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4565 ( .C (clk), .D (key_s0[75]), .Q (new_AGEMA_signal_9602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4569 ( .C (clk), .D (key_s1[75]), .Q (new_AGEMA_signal_9606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4573 ( .C (clk), .D (key_s2[75]), .Q (new_AGEMA_signal_9610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4577 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_9614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4581 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_9618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4585 ( .C (clk), .D (key_s2[76]), .Q (new_AGEMA_signal_9622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4589 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_9626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4593 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_9630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4597 ( .C (clk), .D (key_s2[77]), .Q (new_AGEMA_signal_9634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4601 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_9638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4605 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_9642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4609 ( .C (clk), .D (key_s2[78]), .Q (new_AGEMA_signal_9646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4613 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_9650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4617 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_9654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4621 ( .C (clk), .D (key_s2[79]), .Q (new_AGEMA_signal_9658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4625 ( .C (clk), .D (key_s0[80]), .Q (new_AGEMA_signal_9662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4629 ( .C (clk), .D (key_s1[80]), .Q (new_AGEMA_signal_9666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4633 ( .C (clk), .D (key_s2[80]), .Q (new_AGEMA_signal_9670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4637 ( .C (clk), .D (key_s0[81]), .Q (new_AGEMA_signal_9674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4641 ( .C (clk), .D (key_s1[81]), .Q (new_AGEMA_signal_9678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4645 ( .C (clk), .D (key_s2[81]), .Q (new_AGEMA_signal_9682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4649 ( .C (clk), .D (key_s0[82]), .Q (new_AGEMA_signal_9686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4653 ( .C (clk), .D (key_s1[82]), .Q (new_AGEMA_signal_9690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4657 ( .C (clk), .D (key_s2[82]), .Q (new_AGEMA_signal_9694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4661 ( .C (clk), .D (key_s0[83]), .Q (new_AGEMA_signal_9698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4665 ( .C (clk), .D (key_s1[83]), .Q (new_AGEMA_signal_9702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4669 ( .C (clk), .D (key_s2[83]), .Q (new_AGEMA_signal_9706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4673 ( .C (clk), .D (key_s0[84]), .Q (new_AGEMA_signal_9710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4677 ( .C (clk), .D (key_s1[84]), .Q (new_AGEMA_signal_9714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4681 ( .C (clk), .D (key_s2[84]), .Q (new_AGEMA_signal_9718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4685 ( .C (clk), .D (key_s0[85]), .Q (new_AGEMA_signal_9722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4689 ( .C (clk), .D (key_s1[85]), .Q (new_AGEMA_signal_9726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4693 ( .C (clk), .D (key_s2[85]), .Q (new_AGEMA_signal_9730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4697 ( .C (clk), .D (key_s0[86]), .Q (new_AGEMA_signal_9734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4701 ( .C (clk), .D (key_s1[86]), .Q (new_AGEMA_signal_9738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4705 ( .C (clk), .D (key_s2[86]), .Q (new_AGEMA_signal_9742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4709 ( .C (clk), .D (key_s0[87]), .Q (new_AGEMA_signal_9746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4713 ( .C (clk), .D (key_s1[87]), .Q (new_AGEMA_signal_9750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4717 ( .C (clk), .D (key_s2[87]), .Q (new_AGEMA_signal_9754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4721 ( .C (clk), .D (key_s0[88]), .Q (new_AGEMA_signal_9758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4725 ( .C (clk), .D (key_s1[88]), .Q (new_AGEMA_signal_9762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4729 ( .C (clk), .D (key_s2[88]), .Q (new_AGEMA_signal_9766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4733 ( .C (clk), .D (key_s0[89]), .Q (new_AGEMA_signal_9770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4737 ( .C (clk), .D (key_s1[89]), .Q (new_AGEMA_signal_9774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4741 ( .C (clk), .D (key_s2[89]), .Q (new_AGEMA_signal_9778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4745 ( .C (clk), .D (key_s0[90]), .Q (new_AGEMA_signal_9782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4749 ( .C (clk), .D (key_s1[90]), .Q (new_AGEMA_signal_9786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4753 ( .C (clk), .D (key_s2[90]), .Q (new_AGEMA_signal_9790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4757 ( .C (clk), .D (key_s0[91]), .Q (new_AGEMA_signal_9794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4761 ( .C (clk), .D (key_s1[91]), .Q (new_AGEMA_signal_9798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4765 ( .C (clk), .D (key_s2[91]), .Q (new_AGEMA_signal_9802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4769 ( .C (clk), .D (key_s0[92]), .Q (new_AGEMA_signal_9806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4773 ( .C (clk), .D (key_s1[92]), .Q (new_AGEMA_signal_9810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4777 ( .C (clk), .D (key_s2[92]), .Q (new_AGEMA_signal_9814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4781 ( .C (clk), .D (key_s0[93]), .Q (new_AGEMA_signal_9818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4785 ( .C (clk), .D (key_s1[93]), .Q (new_AGEMA_signal_9822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4789 ( .C (clk), .D (key_s2[93]), .Q (new_AGEMA_signal_9826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4793 ( .C (clk), .D (key_s0[94]), .Q (new_AGEMA_signal_9830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4797 ( .C (clk), .D (key_s1[94]), .Q (new_AGEMA_signal_9834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4801 ( .C (clk), .D (key_s2[94]), .Q (new_AGEMA_signal_9838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4805 ( .C (clk), .D (key_s0[95]), .Q (new_AGEMA_signal_9842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4809 ( .C (clk), .D (key_s1[95]), .Q (new_AGEMA_signal_9846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4813 ( .C (clk), .D (key_s2[95]), .Q (new_AGEMA_signal_9850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4817 ( .C (clk), .D (key_s0[96]), .Q (new_AGEMA_signal_9854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4821 ( .C (clk), .D (key_s1[96]), .Q (new_AGEMA_signal_9858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4825 ( .C (clk), .D (key_s2[96]), .Q (new_AGEMA_signal_9862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4829 ( .C (clk), .D (key_s0[97]), .Q (new_AGEMA_signal_9866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4833 ( .C (clk), .D (key_s1[97]), .Q (new_AGEMA_signal_9870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4837 ( .C (clk), .D (key_s2[97]), .Q (new_AGEMA_signal_9874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4841 ( .C (clk), .D (key_s0[98]), .Q (new_AGEMA_signal_9878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4845 ( .C (clk), .D (key_s1[98]), .Q (new_AGEMA_signal_9882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4849 ( .C (clk), .D (key_s2[98]), .Q (new_AGEMA_signal_9886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4853 ( .C (clk), .D (key_s0[99]), .Q (new_AGEMA_signal_9890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4857 ( .C (clk), .D (key_s1[99]), .Q (new_AGEMA_signal_9894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4861 ( .C (clk), .D (key_s2[99]), .Q (new_AGEMA_signal_9898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4865 ( .C (clk), .D (key_s0[100]), .Q (new_AGEMA_signal_9902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4869 ( .C (clk), .D (key_s1[100]), .Q (new_AGEMA_signal_9906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4873 ( .C (clk), .D (key_s2[100]), .Q (new_AGEMA_signal_9910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4877 ( .C (clk), .D (key_s0[101]), .Q (new_AGEMA_signal_9914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4881 ( .C (clk), .D (key_s1[101]), .Q (new_AGEMA_signal_9918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4885 ( .C (clk), .D (key_s2[101]), .Q (new_AGEMA_signal_9922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4889 ( .C (clk), .D (key_s0[102]), .Q (new_AGEMA_signal_9926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4893 ( .C (clk), .D (key_s1[102]), .Q (new_AGEMA_signal_9930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4897 ( .C (clk), .D (key_s2[102]), .Q (new_AGEMA_signal_9934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4901 ( .C (clk), .D (key_s0[103]), .Q (new_AGEMA_signal_9938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4905 ( .C (clk), .D (key_s1[103]), .Q (new_AGEMA_signal_9942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4909 ( .C (clk), .D (key_s2[103]), .Q (new_AGEMA_signal_9946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4913 ( .C (clk), .D (key_s0[104]), .Q (new_AGEMA_signal_9950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4917 ( .C (clk), .D (key_s1[104]), .Q (new_AGEMA_signal_9954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4921 ( .C (clk), .D (key_s2[104]), .Q (new_AGEMA_signal_9958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4925 ( .C (clk), .D (key_s0[105]), .Q (new_AGEMA_signal_9962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4929 ( .C (clk), .D (key_s1[105]), .Q (new_AGEMA_signal_9966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4933 ( .C (clk), .D (key_s2[105]), .Q (new_AGEMA_signal_9970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4937 ( .C (clk), .D (key_s0[106]), .Q (new_AGEMA_signal_9974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4941 ( .C (clk), .D (key_s1[106]), .Q (new_AGEMA_signal_9978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4945 ( .C (clk), .D (key_s2[106]), .Q (new_AGEMA_signal_9982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4949 ( .C (clk), .D (key_s0[107]), .Q (new_AGEMA_signal_9986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4953 ( .C (clk), .D (key_s1[107]), .Q (new_AGEMA_signal_9990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4957 ( .C (clk), .D (key_s2[107]), .Q (new_AGEMA_signal_9994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4961 ( .C (clk), .D (key_s0[108]), .Q (new_AGEMA_signal_9998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4965 ( .C (clk), .D (key_s1[108]), .Q (new_AGEMA_signal_10002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4969 ( .C (clk), .D (key_s2[108]), .Q (new_AGEMA_signal_10006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4973 ( .C (clk), .D (key_s0[109]), .Q (new_AGEMA_signal_10010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4977 ( .C (clk), .D (key_s1[109]), .Q (new_AGEMA_signal_10014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4981 ( .C (clk), .D (key_s2[109]), .Q (new_AGEMA_signal_10018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4985 ( .C (clk), .D (key_s0[110]), .Q (new_AGEMA_signal_10022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4989 ( .C (clk), .D (key_s1[110]), .Q (new_AGEMA_signal_10026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4993 ( .C (clk), .D (key_s2[110]), .Q (new_AGEMA_signal_10030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4997 ( .C (clk), .D (key_s0[111]), .Q (new_AGEMA_signal_10034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5001 ( .C (clk), .D (key_s1[111]), .Q (new_AGEMA_signal_10038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5005 ( .C (clk), .D (key_s2[111]), .Q (new_AGEMA_signal_10042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5009 ( .C (clk), .D (key_s0[112]), .Q (new_AGEMA_signal_10046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5013 ( .C (clk), .D (key_s1[112]), .Q (new_AGEMA_signal_10050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5017 ( .C (clk), .D (key_s2[112]), .Q (new_AGEMA_signal_10054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5021 ( .C (clk), .D (key_s0[113]), .Q (new_AGEMA_signal_10058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5025 ( .C (clk), .D (key_s1[113]), .Q (new_AGEMA_signal_10062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5029 ( .C (clk), .D (key_s2[113]), .Q (new_AGEMA_signal_10066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5033 ( .C (clk), .D (key_s0[114]), .Q (new_AGEMA_signal_10070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5037 ( .C (clk), .D (key_s1[114]), .Q (new_AGEMA_signal_10074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5041 ( .C (clk), .D (key_s2[114]), .Q (new_AGEMA_signal_10078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5045 ( .C (clk), .D (key_s0[115]), .Q (new_AGEMA_signal_10082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5049 ( .C (clk), .D (key_s1[115]), .Q (new_AGEMA_signal_10086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5053 ( .C (clk), .D (key_s2[115]), .Q (new_AGEMA_signal_10090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5057 ( .C (clk), .D (key_s0[116]), .Q (new_AGEMA_signal_10094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5061 ( .C (clk), .D (key_s1[116]), .Q (new_AGEMA_signal_10098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5065 ( .C (clk), .D (key_s2[116]), .Q (new_AGEMA_signal_10102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5069 ( .C (clk), .D (key_s0[117]), .Q (new_AGEMA_signal_10106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5073 ( .C (clk), .D (key_s1[117]), .Q (new_AGEMA_signal_10110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5077 ( .C (clk), .D (key_s2[117]), .Q (new_AGEMA_signal_10114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5081 ( .C (clk), .D (key_s0[118]), .Q (new_AGEMA_signal_10118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5085 ( .C (clk), .D (key_s1[118]), .Q (new_AGEMA_signal_10122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5089 ( .C (clk), .D (key_s2[118]), .Q (new_AGEMA_signal_10126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5093 ( .C (clk), .D (key_s0[119]), .Q (new_AGEMA_signal_10130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5097 ( .C (clk), .D (key_s1[119]), .Q (new_AGEMA_signal_10134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5101 ( .C (clk), .D (key_s2[119]), .Q (new_AGEMA_signal_10138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5105 ( .C (clk), .D (key_s0[120]), .Q (new_AGEMA_signal_10142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5109 ( .C (clk), .D (key_s1[120]), .Q (new_AGEMA_signal_10146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5113 ( .C (clk), .D (key_s2[120]), .Q (new_AGEMA_signal_10150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5117 ( .C (clk), .D (key_s0[121]), .Q (new_AGEMA_signal_10154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5121 ( .C (clk), .D (key_s1[121]), .Q (new_AGEMA_signal_10158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5125 ( .C (clk), .D (key_s2[121]), .Q (new_AGEMA_signal_10162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5129 ( .C (clk), .D (key_s0[122]), .Q (new_AGEMA_signal_10166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5133 ( .C (clk), .D (key_s1[122]), .Q (new_AGEMA_signal_10170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5137 ( .C (clk), .D (key_s2[122]), .Q (new_AGEMA_signal_10174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5141 ( .C (clk), .D (key_s0[123]), .Q (new_AGEMA_signal_10178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5145 ( .C (clk), .D (key_s1[123]), .Q (new_AGEMA_signal_10182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5149 ( .C (clk), .D (key_s2[123]), .Q (new_AGEMA_signal_10186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5153 ( .C (clk), .D (key_s0[124]), .Q (new_AGEMA_signal_10190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5157 ( .C (clk), .D (key_s1[124]), .Q (new_AGEMA_signal_10194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5161 ( .C (clk), .D (key_s2[124]), .Q (new_AGEMA_signal_10198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5165 ( .C (clk), .D (key_s0[125]), .Q (new_AGEMA_signal_10202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5169 ( .C (clk), .D (key_s1[125]), .Q (new_AGEMA_signal_10206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5173 ( .C (clk), .D (key_s2[125]), .Q (new_AGEMA_signal_10210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5177 ( .C (clk), .D (key_s0[126]), .Q (new_AGEMA_signal_10214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5181 ( .C (clk), .D (key_s1[126]), .Q (new_AGEMA_signal_10218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5185 ( .C (clk), .D (key_s2[126]), .Q (new_AGEMA_signal_10222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5189 ( .C (clk), .D (key_s0[127]), .Q (new_AGEMA_signal_10226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5193 ( .C (clk), .D (key_s1[127]), .Q (new_AGEMA_signal_10230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5197 ( .C (clk), .D (key_s2[127]), .Q (new_AGEMA_signal_10234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5201 ( .C (clk), .D (KSSubBytesInput[9]), .Q (new_AGEMA_signal_10238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5205 ( .C (clk), .D (new_AGEMA_signal_3102), .Q (new_AGEMA_signal_10242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5209 ( .C (clk), .D (new_AGEMA_signal_3103), .Q (new_AGEMA_signal_10246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5213 ( .C (clk), .D (KSSubBytesInput[8]), .Q (new_AGEMA_signal_10250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5217 ( .C (clk), .D (new_AGEMA_signal_3036), .Q (new_AGEMA_signal_10254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5221 ( .C (clk), .D (new_AGEMA_signal_3037), .Q (new_AGEMA_signal_10258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5225 ( .C (clk), .D (KSSubBytesInput[23]), .Q (new_AGEMA_signal_10262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5229 ( .C (clk), .D (new_AGEMA_signal_2970), .Q (new_AGEMA_signal_10266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5233 ( .C (clk), .D (new_AGEMA_signal_2971), .Q (new_AGEMA_signal_10270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5237 ( .C (clk), .D (KSSubBytesInput[22]), .Q (new_AGEMA_signal_10274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5241 ( .C (clk), .D (new_AGEMA_signal_2904), .Q (new_AGEMA_signal_10278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5245 ( .C (clk), .D (new_AGEMA_signal_2905), .Q (new_AGEMA_signal_10282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5249 ( .C (clk), .D (KSSubBytesInput[21]), .Q (new_AGEMA_signal_10286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5253 ( .C (clk), .D (new_AGEMA_signal_2838), .Q (new_AGEMA_signal_10290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5257 ( .C (clk), .D (new_AGEMA_signal_2839), .Q (new_AGEMA_signal_10294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5261 ( .C (clk), .D (KSSubBytesInput[20]), .Q (new_AGEMA_signal_10298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5265 ( .C (clk), .D (new_AGEMA_signal_2772), .Q (new_AGEMA_signal_10302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5269 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_10306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5273 ( .C (clk), .D (RoundKey[41]), .Q (new_AGEMA_signal_10310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5277 ( .C (clk), .D (new_AGEMA_signal_2718), .Q (new_AGEMA_signal_10314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5281 ( .C (clk), .D (new_AGEMA_signal_2719), .Q (new_AGEMA_signal_10318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5285 ( .C (clk), .D (RoundKey[73]), .Q (new_AGEMA_signal_10322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5289 ( .C (clk), .D (new_AGEMA_signal_2928), .Q (new_AGEMA_signal_10326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5293 ( .C (clk), .D (new_AGEMA_signal_2929), .Q (new_AGEMA_signal_10330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5297 ( .C (clk), .D (RoundKey[40]), .Q (new_AGEMA_signal_10334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5301 ( .C (clk), .D (new_AGEMA_signal_2712), .Q (new_AGEMA_signal_10338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5305 ( .C (clk), .D (new_AGEMA_signal_2713), .Q (new_AGEMA_signal_10342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5309 ( .C (clk), .D (RoundKey[72]), .Q (new_AGEMA_signal_10346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5313 ( .C (clk), .D (new_AGEMA_signal_2922), .Q (new_AGEMA_signal_10350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5317 ( .C (clk), .D (new_AGEMA_signal_2923), .Q (new_AGEMA_signal_10354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5321 ( .C (clk), .D (KSSubBytesInput[19]), .Q (new_AGEMA_signal_10358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5325 ( .C (clk), .D (new_AGEMA_signal_2706), .Q (new_AGEMA_signal_10362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5329 ( .C (clk), .D (new_AGEMA_signal_2707), .Q (new_AGEMA_signal_10366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5333 ( .C (clk), .D (RoundKey[39]), .Q (new_AGEMA_signal_10370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5337 ( .C (clk), .D (new_AGEMA_signal_2700), .Q (new_AGEMA_signal_10374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5341 ( .C (clk), .D (new_AGEMA_signal_2701), .Q (new_AGEMA_signal_10378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5345 ( .C (clk), .D (RoundKey[71]), .Q (new_AGEMA_signal_10382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5349 ( .C (clk), .D (new_AGEMA_signal_2916), .Q (new_AGEMA_signal_10386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5353 ( .C (clk), .D (new_AGEMA_signal_2917), .Q (new_AGEMA_signal_10390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5357 ( .C (clk), .D (RoundKey[38]), .Q (new_AGEMA_signal_10394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5361 ( .C (clk), .D (new_AGEMA_signal_2694), .Q (new_AGEMA_signal_10398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5365 ( .C (clk), .D (new_AGEMA_signal_2695), .Q (new_AGEMA_signal_10402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5369 ( .C (clk), .D (RoundKey[70]), .Q (new_AGEMA_signal_10406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5373 ( .C (clk), .D (new_AGEMA_signal_2910), .Q (new_AGEMA_signal_10410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5377 ( .C (clk), .D (new_AGEMA_signal_2911), .Q (new_AGEMA_signal_10414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5381 ( .C (clk), .D (RoundKey[37]), .Q (new_AGEMA_signal_10418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5385 ( .C (clk), .D (new_AGEMA_signal_2688), .Q (new_AGEMA_signal_10422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5389 ( .C (clk), .D (new_AGEMA_signal_2689), .Q (new_AGEMA_signal_10426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5393 ( .C (clk), .D (RoundKey[69]), .Q (new_AGEMA_signal_10430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5397 ( .C (clk), .D (new_AGEMA_signal_2898), .Q (new_AGEMA_signal_10434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5401 ( .C (clk), .D (new_AGEMA_signal_2899), .Q (new_AGEMA_signal_10438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5405 ( .C (clk), .D (RoundKey[36]), .Q (new_AGEMA_signal_10442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5409 ( .C (clk), .D (new_AGEMA_signal_2682), .Q (new_AGEMA_signal_10446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5413 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_10450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5417 ( .C (clk), .D (RoundKey[68]), .Q (new_AGEMA_signal_10454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5421 ( .C (clk), .D (new_AGEMA_signal_2892), .Q (new_AGEMA_signal_10458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5425 ( .C (clk), .D (new_AGEMA_signal_2893), .Q (new_AGEMA_signal_10462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5429 ( .C (clk), .D (RoundKey[35]), .Q (new_AGEMA_signal_10466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5433 ( .C (clk), .D (new_AGEMA_signal_2676), .Q (new_AGEMA_signal_10470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5437 ( .C (clk), .D (new_AGEMA_signal_2677), .Q (new_AGEMA_signal_10474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5441 ( .C (clk), .D (RoundKey[67]), .Q (new_AGEMA_signal_10478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5445 ( .C (clk), .D (new_AGEMA_signal_2886), .Q (new_AGEMA_signal_10482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5449 ( .C (clk), .D (new_AGEMA_signal_2887), .Q (new_AGEMA_signal_10486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5453 ( .C (clk), .D (RoundKey[99]), .Q (new_AGEMA_signal_10490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5457 ( .C (clk), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_10494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5461 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_10498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5465 ( .C (clk), .D (KSSubBytesInput[31]), .Q (new_AGEMA_signal_10502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5469 ( .C (clk), .D (new_AGEMA_signal_2652), .Q (new_AGEMA_signal_10506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5473 ( .C (clk), .D (new_AGEMA_signal_2653), .Q (new_AGEMA_signal_10510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5477 ( .C (clk), .D (RoundKey[63]), .Q (new_AGEMA_signal_10514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5481 ( .C (clk), .D (new_AGEMA_signal_2862), .Q (new_AGEMA_signal_10518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5485 ( .C (clk), .D (new_AGEMA_signal_2863), .Q (new_AGEMA_signal_10522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5489 ( .C (clk), .D (RoundKey[95]), .Q (new_AGEMA_signal_10526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5493 ( .C (clk), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_10530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5497 ( .C (clk), .D (new_AGEMA_signal_3073), .Q (new_AGEMA_signal_10534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5501 ( .C (clk), .D (KSSubBytesInput[30]), .Q (new_AGEMA_signal_10538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5505 ( .C (clk), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_10542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5509 ( .C (clk), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_10546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5513 ( .C (clk), .D (RoundKey[62]), .Q (new_AGEMA_signal_10550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5517 ( .C (clk), .D (new_AGEMA_signal_2856), .Q (new_AGEMA_signal_10554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5521 ( .C (clk), .D (new_AGEMA_signal_2857), .Q (new_AGEMA_signal_10558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5525 ( .C (clk), .D (RoundKey[94]), .Q (new_AGEMA_signal_10562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5529 ( .C (clk), .D (new_AGEMA_signal_3066), .Q (new_AGEMA_signal_10566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5533 ( .C (clk), .D (new_AGEMA_signal_3067), .Q (new_AGEMA_signal_10570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5537 ( .C (clk), .D (KSSubBytesInput[18]), .Q (new_AGEMA_signal_10574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5541 ( .C (clk), .D (new_AGEMA_signal_2640), .Q (new_AGEMA_signal_10578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5545 ( .C (clk), .D (new_AGEMA_signal_2641), .Q (new_AGEMA_signal_10582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5549 ( .C (clk), .D (RoundKey[34]), .Q (new_AGEMA_signal_10586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5553 ( .C (clk), .D (new_AGEMA_signal_2670), .Q (new_AGEMA_signal_10590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5557 ( .C (clk), .D (new_AGEMA_signal_2671), .Q (new_AGEMA_signal_10594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5561 ( .C (clk), .D (RoundKey[66]), .Q (new_AGEMA_signal_10598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5565 ( .C (clk), .D (new_AGEMA_signal_2880), .Q (new_AGEMA_signal_10602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5569 ( .C (clk), .D (new_AGEMA_signal_2881), .Q (new_AGEMA_signal_10606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5573 ( .C (clk), .D (RoundKey[98]), .Q (new_AGEMA_signal_10610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5577 ( .C (clk), .D (new_AGEMA_signal_3090), .Q (new_AGEMA_signal_10614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5581 ( .C (clk), .D (new_AGEMA_signal_3091), .Q (new_AGEMA_signal_10618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5585 ( .C (clk), .D (KSSubBytesInput[29]), .Q (new_AGEMA_signal_10622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5589 ( .C (clk), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_10626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5593 ( .C (clk), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_10630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5597 ( .C (clk), .D (RoundKey[61]), .Q (new_AGEMA_signal_10634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5601 ( .C (clk), .D (new_AGEMA_signal_2850), .Q (new_AGEMA_signal_10638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5605 ( .C (clk), .D (new_AGEMA_signal_2851), .Q (new_AGEMA_signal_10642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5609 ( .C (clk), .D (RoundKey[93]), .Q (new_AGEMA_signal_10646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5613 ( .C (clk), .D (new_AGEMA_signal_3060), .Q (new_AGEMA_signal_10650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5617 ( .C (clk), .D (new_AGEMA_signal_3061), .Q (new_AGEMA_signal_10654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5621 ( .C (clk), .D (KSSubBytesInput[28]), .Q (new_AGEMA_signal_10658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5625 ( .C (clk), .D (new_AGEMA_signal_2628), .Q (new_AGEMA_signal_10662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5629 ( .C (clk), .D (new_AGEMA_signal_2629), .Q (new_AGEMA_signal_10666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5633 ( .C (clk), .D (RoundKey[60]), .Q (new_AGEMA_signal_10670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5637 ( .C (clk), .D (new_AGEMA_signal_2844), .Q (new_AGEMA_signal_10674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5641 ( .C (clk), .D (new_AGEMA_signal_2845), .Q (new_AGEMA_signal_10678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5645 ( .C (clk), .D (RoundKey[92]), .Q (new_AGEMA_signal_10682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5649 ( .C (clk), .D (new_AGEMA_signal_3054), .Q (new_AGEMA_signal_10686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5653 ( .C (clk), .D (new_AGEMA_signal_3055), .Q (new_AGEMA_signal_10690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5657 ( .C (clk), .D (KSSubBytesInput[27]), .Q (new_AGEMA_signal_10694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5661 ( .C (clk), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_10698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5665 ( .C (clk), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_10702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5669 ( .C (clk), .D (RoundKey[59]), .Q (new_AGEMA_signal_10706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5673 ( .C (clk), .D (new_AGEMA_signal_2832), .Q (new_AGEMA_signal_10710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5677 ( .C (clk), .D (new_AGEMA_signal_2833), .Q (new_AGEMA_signal_10714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5681 ( .C (clk), .D (RoundKey[91]), .Q (new_AGEMA_signal_10718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5685 ( .C (clk), .D (new_AGEMA_signal_3048), .Q (new_AGEMA_signal_10722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5689 ( .C (clk), .D (new_AGEMA_signal_3049), .Q (new_AGEMA_signal_10726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5693 ( .C (clk), .D (KSSubBytesInput[26]), .Q (new_AGEMA_signal_10730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5697 ( .C (clk), .D (new_AGEMA_signal_2616), .Q (new_AGEMA_signal_10734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5701 ( .C (clk), .D (new_AGEMA_signal_2617), .Q (new_AGEMA_signal_10738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5705 ( .C (clk), .D (RoundKey[58]), .Q (new_AGEMA_signal_10742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5709 ( .C (clk), .D (new_AGEMA_signal_2826), .Q (new_AGEMA_signal_10746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5713 ( .C (clk), .D (new_AGEMA_signal_2827), .Q (new_AGEMA_signal_10750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5717 ( .C (clk), .D (RoundKey[90]), .Q (new_AGEMA_signal_10754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5721 ( .C (clk), .D (new_AGEMA_signal_3042), .Q (new_AGEMA_signal_10758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5725 ( .C (clk), .D (new_AGEMA_signal_3043), .Q (new_AGEMA_signal_10762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5729 ( .C (clk), .D (KSSubBytesInput[25]), .Q (new_AGEMA_signal_10766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5733 ( .C (clk), .D (new_AGEMA_signal_2610), .Q (new_AGEMA_signal_10770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5737 ( .C (clk), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_10774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5741 ( .C (clk), .D (RoundKey[57]), .Q (new_AGEMA_signal_10778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5745 ( .C (clk), .D (new_AGEMA_signal_2820), .Q (new_AGEMA_signal_10782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5749 ( .C (clk), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_10786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5753 ( .C (clk), .D (RoundKey[89]), .Q (new_AGEMA_signal_10790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5757 ( .C (clk), .D (new_AGEMA_signal_3030), .Q (new_AGEMA_signal_10794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5761 ( .C (clk), .D (new_AGEMA_signal_3031), .Q (new_AGEMA_signal_10798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5765 ( .C (clk), .D (KSSubBytesInput[24]), .Q (new_AGEMA_signal_10802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5769 ( .C (clk), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_10806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5773 ( .C (clk), .D (new_AGEMA_signal_2605), .Q (new_AGEMA_signal_10810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5777 ( .C (clk), .D (RoundKey[56]), .Q (new_AGEMA_signal_10814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5781 ( .C (clk), .D (new_AGEMA_signal_2814), .Q (new_AGEMA_signal_10818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5785 ( .C (clk), .D (new_AGEMA_signal_2815), .Q (new_AGEMA_signal_10822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5789 ( .C (clk), .D (RoundKey[88]), .Q (new_AGEMA_signal_10826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5793 ( .C (clk), .D (new_AGEMA_signal_3024), .Q (new_AGEMA_signal_10830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5797 ( .C (clk), .D (new_AGEMA_signal_3025), .Q (new_AGEMA_signal_10834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5801 ( .C (clk), .D (KSSubBytesInput[7]), .Q (new_AGEMA_signal_10838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5805 ( .C (clk), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_10842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5809 ( .C (clk), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_10846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5813 ( .C (clk), .D (RoundKey[55]), .Q (new_AGEMA_signal_10850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5817 ( .C (clk), .D (new_AGEMA_signal_2808), .Q (new_AGEMA_signal_10854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5821 ( .C (clk), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_10858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5825 ( .C (clk), .D (RoundKey[87]), .Q (new_AGEMA_signal_10862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5829 ( .C (clk), .D (new_AGEMA_signal_3018), .Q (new_AGEMA_signal_10866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5833 ( .C (clk), .D (new_AGEMA_signal_3019), .Q (new_AGEMA_signal_10870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5837 ( .C (clk), .D (KSSubBytesInput[6]), .Q (new_AGEMA_signal_10874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5841 ( .C (clk), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_10878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5845 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_10882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5849 ( .C (clk), .D (RoundKey[54]), .Q (new_AGEMA_signal_10886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5853 ( .C (clk), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_10890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5857 ( .C (clk), .D (new_AGEMA_signal_2803), .Q (new_AGEMA_signal_10894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5861 ( .C (clk), .D (RoundKey[86]), .Q (new_AGEMA_signal_10898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5865 ( .C (clk), .D (new_AGEMA_signal_3012), .Q (new_AGEMA_signal_10902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5869 ( .C (clk), .D (new_AGEMA_signal_3013), .Q (new_AGEMA_signal_10906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5873 ( .C (clk), .D (KSSubBytesInput[5]), .Q (new_AGEMA_signal_10910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5877 ( .C (clk), .D (new_AGEMA_signal_2586), .Q (new_AGEMA_signal_10914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5881 ( .C (clk), .D (new_AGEMA_signal_2587), .Q (new_AGEMA_signal_10918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5885 ( .C (clk), .D (RoundKey[53]), .Q (new_AGEMA_signal_10922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5889 ( .C (clk), .D (new_AGEMA_signal_2796), .Q (new_AGEMA_signal_10926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5893 ( .C (clk), .D (new_AGEMA_signal_2797), .Q (new_AGEMA_signal_10930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5897 ( .C (clk), .D (RoundKey[85]), .Q (new_AGEMA_signal_10934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5901 ( .C (clk), .D (new_AGEMA_signal_3006), .Q (new_AGEMA_signal_10938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5905 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (new_AGEMA_signal_10942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5909 ( .C (clk), .D (KSSubBytesInput[4]), .Q (new_AGEMA_signal_10946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5913 ( .C (clk), .D (new_AGEMA_signal_2580), .Q (new_AGEMA_signal_10950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5917 ( .C (clk), .D (new_AGEMA_signal_2581), .Q (new_AGEMA_signal_10954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5921 ( .C (clk), .D (RoundKey[52]), .Q (new_AGEMA_signal_10958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5925 ( .C (clk), .D (new_AGEMA_signal_2790), .Q (new_AGEMA_signal_10962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5929 ( .C (clk), .D (new_AGEMA_signal_2791), .Q (new_AGEMA_signal_10966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5933 ( .C (clk), .D (RoundKey[84]), .Q (new_AGEMA_signal_10970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5937 ( .C (clk), .D (new_AGEMA_signal_3000), .Q (new_AGEMA_signal_10974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5941 ( .C (clk), .D (new_AGEMA_signal_3001), .Q (new_AGEMA_signal_10978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5945 ( .C (clk), .D (KSSubBytesInput[17]), .Q (new_AGEMA_signal_10982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5949 ( .C (clk), .D (new_AGEMA_signal_2574), .Q (new_AGEMA_signal_10986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5953 ( .C (clk), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_10990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5957 ( .C (clk), .D (RoundKey[33]), .Q (new_AGEMA_signal_10994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5961 ( .C (clk), .D (new_AGEMA_signal_2664), .Q (new_AGEMA_signal_10998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5965 ( .C (clk), .D (new_AGEMA_signal_2665), .Q (new_AGEMA_signal_11002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5969 ( .C (clk), .D (RoundKey[65]), .Q (new_AGEMA_signal_11006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5973 ( .C (clk), .D (new_AGEMA_signal_2874), .Q (new_AGEMA_signal_11010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5977 ( .C (clk), .D (new_AGEMA_signal_2875), .Q (new_AGEMA_signal_11014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5981 ( .C (clk), .D (RoundKey[97]), .Q (new_AGEMA_signal_11018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5985 ( .C (clk), .D (new_AGEMA_signal_3084), .Q (new_AGEMA_signal_11022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5989 ( .C (clk), .D (new_AGEMA_signal_3085), .Q (new_AGEMA_signal_11026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5993 ( .C (clk), .D (KSSubBytesInput[3]), .Q (new_AGEMA_signal_11030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5997 ( .C (clk), .D (new_AGEMA_signal_2568), .Q (new_AGEMA_signal_11034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6001 ( .C (clk), .D (new_AGEMA_signal_2569), .Q (new_AGEMA_signal_11038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6005 ( .C (clk), .D (RoundKey[51]), .Q (new_AGEMA_signal_11042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6009 ( .C (clk), .D (new_AGEMA_signal_2784), .Q (new_AGEMA_signal_11046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6013 ( .C (clk), .D (new_AGEMA_signal_2785), .Q (new_AGEMA_signal_11050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6017 ( .C (clk), .D (RoundKey[83]), .Q (new_AGEMA_signal_11054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6021 ( .C (clk), .D (new_AGEMA_signal_2994), .Q (new_AGEMA_signal_11058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6025 ( .C (clk), .D (new_AGEMA_signal_2995), .Q (new_AGEMA_signal_11062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6029 ( .C (clk), .D (KSSubBytesInput[2]), .Q (new_AGEMA_signal_11066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6033 ( .C (clk), .D (new_AGEMA_signal_2562), .Q (new_AGEMA_signal_11070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6037 ( .C (clk), .D (new_AGEMA_signal_2563), .Q (new_AGEMA_signal_11074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6041 ( .C (clk), .D (RoundKey[50]), .Q (new_AGEMA_signal_11078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6045 ( .C (clk), .D (new_AGEMA_signal_2778), .Q (new_AGEMA_signal_11082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6049 ( .C (clk), .D (new_AGEMA_signal_2779), .Q (new_AGEMA_signal_11086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6053 ( .C (clk), .D (RoundKey[82]), .Q (new_AGEMA_signal_11090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6057 ( .C (clk), .D (new_AGEMA_signal_2988), .Q (new_AGEMA_signal_11094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6061 ( .C (clk), .D (new_AGEMA_signal_2989), .Q (new_AGEMA_signal_11098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6065 ( .C (clk), .D (KSSubBytesInput[1]), .Q (new_AGEMA_signal_11102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6069 ( .C (clk), .D (new_AGEMA_signal_2556), .Q (new_AGEMA_signal_11106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6073 ( .C (clk), .D (new_AGEMA_signal_2557), .Q (new_AGEMA_signal_11110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6077 ( .C (clk), .D (RoundKey[49]), .Q (new_AGEMA_signal_11114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6081 ( .C (clk), .D (new_AGEMA_signal_2766), .Q (new_AGEMA_signal_11118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6085 ( .C (clk), .D (new_AGEMA_signal_2767), .Q (new_AGEMA_signal_11122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6089 ( .C (clk), .D (RoundKey[81]), .Q (new_AGEMA_signal_11126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6093 ( .C (clk), .D (new_AGEMA_signal_2982), .Q (new_AGEMA_signal_11130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6097 ( .C (clk), .D (new_AGEMA_signal_2983), .Q (new_AGEMA_signal_11134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6101 ( .C (clk), .D (KSSubBytesInput[0]), .Q (new_AGEMA_signal_11138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6105 ( .C (clk), .D (new_AGEMA_signal_2550), .Q (new_AGEMA_signal_11142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6109 ( .C (clk), .D (new_AGEMA_signal_2551), .Q (new_AGEMA_signal_11146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6113 ( .C (clk), .D (RoundKey[48]), .Q (new_AGEMA_signal_11150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6117 ( .C (clk), .D (new_AGEMA_signal_2760), .Q (new_AGEMA_signal_11154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6121 ( .C (clk), .D (new_AGEMA_signal_2761), .Q (new_AGEMA_signal_11158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6125 ( .C (clk), .D (RoundKey[80]), .Q (new_AGEMA_signal_11162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6129 ( .C (clk), .D (new_AGEMA_signal_2976), .Q (new_AGEMA_signal_11166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6133 ( .C (clk), .D (new_AGEMA_signal_2977), .Q (new_AGEMA_signal_11170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6137 ( .C (clk), .D (KSSubBytesInput[15]), .Q (new_AGEMA_signal_11174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6141 ( .C (clk), .D (new_AGEMA_signal_2544), .Q (new_AGEMA_signal_11178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6145 ( .C (clk), .D (new_AGEMA_signal_2545), .Q (new_AGEMA_signal_11182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6149 ( .C (clk), .D (RoundKey[47]), .Q (new_AGEMA_signal_11186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6153 ( .C (clk), .D (new_AGEMA_signal_2754), .Q (new_AGEMA_signal_11190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6157 ( .C (clk), .D (new_AGEMA_signal_2755), .Q (new_AGEMA_signal_11194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6161 ( .C (clk), .D (RoundKey[79]), .Q (new_AGEMA_signal_11198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6165 ( .C (clk), .D (new_AGEMA_signal_2964), .Q (new_AGEMA_signal_11202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6169 ( .C (clk), .D (new_AGEMA_signal_2965), .Q (new_AGEMA_signal_11206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6173 ( .C (clk), .D (KSSubBytesInput[14]), .Q (new_AGEMA_signal_11210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6177 ( .C (clk), .D (new_AGEMA_signal_2538), .Q (new_AGEMA_signal_11214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6181 ( .C (clk), .D (new_AGEMA_signal_2539), .Q (new_AGEMA_signal_11218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6185 ( .C (clk), .D (RoundKey[46]), .Q (new_AGEMA_signal_11222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6189 ( .C (clk), .D (new_AGEMA_signal_2748), .Q (new_AGEMA_signal_11226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6193 ( .C (clk), .D (new_AGEMA_signal_2749), .Q (new_AGEMA_signal_11230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6197 ( .C (clk), .D (RoundKey[78]), .Q (new_AGEMA_signal_11234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6201 ( .C (clk), .D (new_AGEMA_signal_2958), .Q (new_AGEMA_signal_11238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6205 ( .C (clk), .D (new_AGEMA_signal_2959), .Q (new_AGEMA_signal_11242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6209 ( .C (clk), .D (KSSubBytesInput[13]), .Q (new_AGEMA_signal_11246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6213 ( .C (clk), .D (new_AGEMA_signal_2532), .Q (new_AGEMA_signal_11250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6217 ( .C (clk), .D (new_AGEMA_signal_2533), .Q (new_AGEMA_signal_11254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6221 ( .C (clk), .D (RoundKey[45]), .Q (new_AGEMA_signal_11258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6225 ( .C (clk), .D (new_AGEMA_signal_2742), .Q (new_AGEMA_signal_11262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6229 ( .C (clk), .D (new_AGEMA_signal_2743), .Q (new_AGEMA_signal_11266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6233 ( .C (clk), .D (RoundKey[77]), .Q (new_AGEMA_signal_11270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6237 ( .C (clk), .D (new_AGEMA_signal_2952), .Q (new_AGEMA_signal_11274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6241 ( .C (clk), .D (new_AGEMA_signal_2953), .Q (new_AGEMA_signal_11278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6245 ( .C (clk), .D (KSSubBytesInput[12]), .Q (new_AGEMA_signal_11282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6249 ( .C (clk), .D (new_AGEMA_signal_2526), .Q (new_AGEMA_signal_11286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6253 ( .C (clk), .D (new_AGEMA_signal_2527), .Q (new_AGEMA_signal_11290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6257 ( .C (clk), .D (RoundKey[44]), .Q (new_AGEMA_signal_11294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6261 ( .C (clk), .D (new_AGEMA_signal_2736), .Q (new_AGEMA_signal_11298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6265 ( .C (clk), .D (new_AGEMA_signal_2737), .Q (new_AGEMA_signal_11302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6269 ( .C (clk), .D (RoundKey[76]), .Q (new_AGEMA_signal_11306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6273 ( .C (clk), .D (new_AGEMA_signal_2946), .Q (new_AGEMA_signal_11310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6277 ( .C (clk), .D (new_AGEMA_signal_2947), .Q (new_AGEMA_signal_11314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6281 ( .C (clk), .D (RoundKey[127]), .Q (new_AGEMA_signal_11318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6285 ( .C (clk), .D (new_AGEMA_signal_2520), .Q (new_AGEMA_signal_11322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6289 ( .C (clk), .D (new_AGEMA_signal_2521), .Q (new_AGEMA_signal_11326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6293 ( .C (clk), .D (RoundKey[126]), .Q (new_AGEMA_signal_11330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6297 ( .C (clk), .D (new_AGEMA_signal_2514), .Q (new_AGEMA_signal_11334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6301 ( .C (clk), .D (new_AGEMA_signal_2515), .Q (new_AGEMA_signal_11338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6305 ( .C (clk), .D (RoundKey[125]), .Q (new_AGEMA_signal_11342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6309 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_11346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6313 ( .C (clk), .D (new_AGEMA_signal_2509), .Q (new_AGEMA_signal_11350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6317 ( .C (clk), .D (RoundKey[124]), .Q (new_AGEMA_signal_11354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6321 ( .C (clk), .D (new_AGEMA_signal_2502), .Q (new_AGEMA_signal_11358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6325 ( .C (clk), .D (new_AGEMA_signal_2503), .Q (new_AGEMA_signal_11362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6329 ( .C (clk), .D (RoundKey[123]), .Q (new_AGEMA_signal_11366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6333 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_11370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6337 ( .C (clk), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_11374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6341 ( .C (clk), .D (RoundKey[122]), .Q (new_AGEMA_signal_11378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6345 ( .C (clk), .D (new_AGEMA_signal_2490), .Q (new_AGEMA_signal_11382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6349 ( .C (clk), .D (new_AGEMA_signal_2491), .Q (new_AGEMA_signal_11386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6353 ( .C (clk), .D (RoundKey[121]), .Q (new_AGEMA_signal_11390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6357 ( .C (clk), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_11394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6361 ( .C (clk), .D (new_AGEMA_signal_2485), .Q (new_AGEMA_signal_11398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6365 ( .C (clk), .D (RoundKey[120]), .Q (new_AGEMA_signal_11402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6369 ( .C (clk), .D (new_AGEMA_signal_2478), .Q (new_AGEMA_signal_11406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6373 ( .C (clk), .D (new_AGEMA_signal_2479), .Q (new_AGEMA_signal_11410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6377 ( .C (clk), .D (KSSubBytesInput[11]), .Q (new_AGEMA_signal_11414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6381 ( .C (clk), .D (new_AGEMA_signal_2472), .Q (new_AGEMA_signal_11418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6385 ( .C (clk), .D (new_AGEMA_signal_2473), .Q (new_AGEMA_signal_11422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6389 ( .C (clk), .D (RoundKey[43]), .Q (new_AGEMA_signal_11426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6393 ( .C (clk), .D (new_AGEMA_signal_2730), .Q (new_AGEMA_signal_11430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6397 ( .C (clk), .D (new_AGEMA_signal_2731), .Q (new_AGEMA_signal_11434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6401 ( .C (clk), .D (RoundKey[75]), .Q (new_AGEMA_signal_11438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6405 ( .C (clk), .D (new_AGEMA_signal_2940), .Q (new_AGEMA_signal_11442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6409 ( .C (clk), .D (new_AGEMA_signal_2941), .Q (new_AGEMA_signal_11446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6413 ( .C (clk), .D (RoundKey[119]), .Q (new_AGEMA_signal_11450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6417 ( .C (clk), .D (new_AGEMA_signal_2466), .Q (new_AGEMA_signal_11454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6421 ( .C (clk), .D (new_AGEMA_signal_2467), .Q (new_AGEMA_signal_11458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6425 ( .C (clk), .D (RoundKey[118]), .Q (new_AGEMA_signal_11462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6429 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_11466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6433 ( .C (clk), .D (new_AGEMA_signal_2461), .Q (new_AGEMA_signal_11470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6437 ( .C (clk), .D (RoundKey[117]), .Q (new_AGEMA_signal_11474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6441 ( .C (clk), .D (new_AGEMA_signal_2454), .Q (new_AGEMA_signal_11478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6445 ( .C (clk), .D (new_AGEMA_signal_2455), .Q (new_AGEMA_signal_11482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6449 ( .C (clk), .D (RoundKey[116]), .Q (new_AGEMA_signal_11486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6453 ( .C (clk), .D (new_AGEMA_signal_2448), .Q (new_AGEMA_signal_11490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6457 ( .C (clk), .D (new_AGEMA_signal_2449), .Q (new_AGEMA_signal_11494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6461 ( .C (clk), .D (RoundKey[115]), .Q (new_AGEMA_signal_11498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6465 ( .C (clk), .D (new_AGEMA_signal_2442), .Q (new_AGEMA_signal_11502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6469 ( .C (clk), .D (new_AGEMA_signal_2443), .Q (new_AGEMA_signal_11506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6473 ( .C (clk), .D (RoundKey[114]), .Q (new_AGEMA_signal_11510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6477 ( .C (clk), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_11514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6481 ( .C (clk), .D (new_AGEMA_signal_2437), .Q (new_AGEMA_signal_11518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6485 ( .C (clk), .D (RoundKey[113]), .Q (new_AGEMA_signal_11522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6489 ( .C (clk), .D (new_AGEMA_signal_2430), .Q (new_AGEMA_signal_11526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6493 ( .C (clk), .D (new_AGEMA_signal_2431), .Q (new_AGEMA_signal_11530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6497 ( .C (clk), .D (RoundKey[112]), .Q (new_AGEMA_signal_11534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6501 ( .C (clk), .D (new_AGEMA_signal_2424), .Q (new_AGEMA_signal_11538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6505 ( .C (clk), .D (new_AGEMA_signal_2425), .Q (new_AGEMA_signal_11542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6509 ( .C (clk), .D (RoundKey[111]), .Q (new_AGEMA_signal_11546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6513 ( .C (clk), .D (new_AGEMA_signal_2418), .Q (new_AGEMA_signal_11550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6517 ( .C (clk), .D (new_AGEMA_signal_2419), .Q (new_AGEMA_signal_11554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6521 ( .C (clk), .D (RoundKey[110]), .Q (new_AGEMA_signal_11558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6525 ( .C (clk), .D (new_AGEMA_signal_2412), .Q (new_AGEMA_signal_11562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6529 ( .C (clk), .D (new_AGEMA_signal_2413), .Q (new_AGEMA_signal_11566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6533 ( .C (clk), .D (KSSubBytesInput[10]), .Q (new_AGEMA_signal_11570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6537 ( .C (clk), .D (new_AGEMA_signal_2406), .Q (new_AGEMA_signal_11574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6541 ( .C (clk), .D (new_AGEMA_signal_2407), .Q (new_AGEMA_signal_11578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6545 ( .C (clk), .D (RoundKey[42]), .Q (new_AGEMA_signal_11582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6549 ( .C (clk), .D (new_AGEMA_signal_2724), .Q (new_AGEMA_signal_11586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6553 ( .C (clk), .D (new_AGEMA_signal_2725), .Q (new_AGEMA_signal_11590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6557 ( .C (clk), .D (RoundKey[74]), .Q (new_AGEMA_signal_11594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6561 ( .C (clk), .D (new_AGEMA_signal_2934), .Q (new_AGEMA_signal_11598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6565 ( .C (clk), .D (new_AGEMA_signal_2935), .Q (new_AGEMA_signal_11602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6569 ( .C (clk), .D (RoundKey[109]), .Q (new_AGEMA_signal_11606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6573 ( .C (clk), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_11610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6577 ( .C (clk), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_11614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6581 ( .C (clk), .D (RoundKey[108]), .Q (new_AGEMA_signal_11618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6585 ( .C (clk), .D (new_AGEMA_signal_2394), .Q (new_AGEMA_signal_11622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6589 ( .C (clk), .D (new_AGEMA_signal_2395), .Q (new_AGEMA_signal_11626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6593 ( .C (clk), .D (RoundKey[107]), .Q (new_AGEMA_signal_11630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6597 ( .C (clk), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_11634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6601 ( .C (clk), .D (new_AGEMA_signal_2389), .Q (new_AGEMA_signal_11638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6605 ( .C (clk), .D (RoundKey[106]), .Q (new_AGEMA_signal_11642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6609 ( .C (clk), .D (new_AGEMA_signal_2382), .Q (new_AGEMA_signal_11646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6613 ( .C (clk), .D (new_AGEMA_signal_2383), .Q (new_AGEMA_signal_11650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6617 ( .C (clk), .D (RoundKey[105]), .Q (new_AGEMA_signal_11654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6621 ( .C (clk), .D (new_AGEMA_signal_2376), .Q (new_AGEMA_signal_11658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6625 ( .C (clk), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_11662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6629 ( .C (clk), .D (RoundKey[104]), .Q (new_AGEMA_signal_11666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6633 ( .C (clk), .D (new_AGEMA_signal_2370), .Q (new_AGEMA_signal_11670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6637 ( .C (clk), .D (new_AGEMA_signal_2371), .Q (new_AGEMA_signal_11674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6641 ( .C (clk), .D (RoundKey[103]), .Q (new_AGEMA_signal_11678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6645 ( .C (clk), .D (new_AGEMA_signal_2364), .Q (new_AGEMA_signal_11682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6649 ( .C (clk), .D (new_AGEMA_signal_2365), .Q (new_AGEMA_signal_11686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6653 ( .C (clk), .D (RoundKey[102]), .Q (new_AGEMA_signal_11690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6657 ( .C (clk), .D (new_AGEMA_signal_2358), .Q (new_AGEMA_signal_11694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6661 ( .C (clk), .D (new_AGEMA_signal_2359), .Q (new_AGEMA_signal_11698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6665 ( .C (clk), .D (RoundKey[101]), .Q (new_AGEMA_signal_11702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6669 ( .C (clk), .D (new_AGEMA_signal_2352), .Q (new_AGEMA_signal_11706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6673 ( .C (clk), .D (new_AGEMA_signal_2353), .Q (new_AGEMA_signal_11710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6677 ( .C (clk), .D (RoundKey[100]), .Q (new_AGEMA_signal_11714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6681 ( .C (clk), .D (new_AGEMA_signal_2346), .Q (new_AGEMA_signal_11718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6685 ( .C (clk), .D (new_AGEMA_signal_2347), .Q (new_AGEMA_signal_11722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6689 ( .C (clk), .D (KSSubBytesInput[16]), .Q (new_AGEMA_signal_11726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6693 ( .C (clk), .D (new_AGEMA_signal_2340), .Q (new_AGEMA_signal_11730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6697 ( .C (clk), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_11734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6701 ( .C (clk), .D (RoundKey[32]), .Q (new_AGEMA_signal_11738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6705 ( .C (clk), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_11742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6709 ( .C (clk), .D (new_AGEMA_signal_2659), .Q (new_AGEMA_signal_11746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6713 ( .C (clk), .D (RoundKey[64]), .Q (new_AGEMA_signal_11750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6717 ( .C (clk), .D (new_AGEMA_signal_2868), .Q (new_AGEMA_signal_11754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6721 ( .C (clk), .D (new_AGEMA_signal_2869), .Q (new_AGEMA_signal_11758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6725 ( .C (clk), .D (RoundKey[96]), .Q (new_AGEMA_signal_11762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6729 ( .C (clk), .D (new_AGEMA_signal_3078), .Q (new_AGEMA_signal_11766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6733 ( .C (clk), .D (new_AGEMA_signal_3079), .Q (new_AGEMA_signal_11770) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C (clk), .D (Rcon[7]), .Q (new_AGEMA_signal_11774) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C (clk), .D (Rcon[6]), .Q (new_AGEMA_signal_11778) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C (clk), .D (Rcon[5]), .Q (new_AGEMA_signal_11782) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C (clk), .D (Rcon[4]), .Q (new_AGEMA_signal_11786) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C (clk), .D (Rcon[3]), .Q (new_AGEMA_signal_11790) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C (clk), .D (Rcon[2]), .Q (new_AGEMA_signal_11794) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C (clk), .D (Rcon[1]), .Q (new_AGEMA_signal_11798) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C (clk), .D (Rcon[0]), .Q (new_AGEMA_signal_11802) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C (clk), .D (MuxKeyExpansion_n15), .Q (new_AGEMA_signal_11806) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C (clk), .D (MuxKeyExpansion_n16), .Q (new_AGEMA_signal_11810) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C (clk), .D (MuxKeyExpansion_n17), .Q (new_AGEMA_signal_11814) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C (clk), .D (MuxKeyExpansion_n18), .Q (new_AGEMA_signal_11818) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C (clk), .D (MuxKeyExpansion_n19), .Q (new_AGEMA_signal_11822) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C (clk), .D (MuxKeyExpansion_n20), .Q (new_AGEMA_signal_11826) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C (clk), .D (MuxKeyExpansion_n14), .Q (new_AGEMA_signal_11830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6797 ( .C (clk), .D (RoundReg_Inst_ff_SDE_32_next_state), .Q (new_AGEMA_signal_11834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6801 ( .C (clk), .D (new_AGEMA_signal_3364), .Q (new_AGEMA_signal_11838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6805 ( .C (clk), .D (new_AGEMA_signal_3365), .Q (new_AGEMA_signal_11842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6809 ( .C (clk), .D (RoundReg_Inst_ff_SDE_33_next_state), .Q (new_AGEMA_signal_11846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6813 ( .C (clk), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_11850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6817 ( .C (clk), .D (new_AGEMA_signal_3369), .Q (new_AGEMA_signal_11854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6821 ( .C (clk), .D (RoundReg_Inst_ff_SDE_34_next_state), .Q (new_AGEMA_signal_11858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6825 ( .C (clk), .D (new_AGEMA_signal_3372), .Q (new_AGEMA_signal_11862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6829 ( .C (clk), .D (new_AGEMA_signal_3373), .Q (new_AGEMA_signal_11866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6833 ( .C (clk), .D (RoundReg_Inst_ff_SDE_35_next_state), .Q (new_AGEMA_signal_11870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6837 ( .C (clk), .D (new_AGEMA_signal_3376), .Q (new_AGEMA_signal_11874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6841 ( .C (clk), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_11878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6845 ( .C (clk), .D (RoundReg_Inst_ff_SDE_36_next_state), .Q (new_AGEMA_signal_11882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6849 ( .C (clk), .D (new_AGEMA_signal_3380), .Q (new_AGEMA_signal_11886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6853 ( .C (clk), .D (new_AGEMA_signal_3381), .Q (new_AGEMA_signal_11890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6857 ( .C (clk), .D (RoundReg_Inst_ff_SDE_37_next_state), .Q (new_AGEMA_signal_11894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6861 ( .C (clk), .D (new_AGEMA_signal_3384), .Q (new_AGEMA_signal_11898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6865 ( .C (clk), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_11902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6869 ( .C (clk), .D (RoundReg_Inst_ff_SDE_38_next_state), .Q (new_AGEMA_signal_11906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6873 ( .C (clk), .D (new_AGEMA_signal_3388), .Q (new_AGEMA_signal_11910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6877 ( .C (clk), .D (new_AGEMA_signal_3389), .Q (new_AGEMA_signal_11914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6881 ( .C (clk), .D (RoundReg_Inst_ff_SDE_39_next_state), .Q (new_AGEMA_signal_11918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6885 ( .C (clk), .D (new_AGEMA_signal_3392), .Q (new_AGEMA_signal_11922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6889 ( .C (clk), .D (new_AGEMA_signal_3393), .Q (new_AGEMA_signal_11926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6893 ( .C (clk), .D (RoundReg_Inst_ff_SDE_40_next_state), .Q (new_AGEMA_signal_11930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6897 ( .C (clk), .D (new_AGEMA_signal_3396), .Q (new_AGEMA_signal_11934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6901 ( .C (clk), .D (new_AGEMA_signal_3397), .Q (new_AGEMA_signal_11938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6905 ( .C (clk), .D (RoundReg_Inst_ff_SDE_41_next_state), .Q (new_AGEMA_signal_11942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6909 ( .C (clk), .D (new_AGEMA_signal_3400), .Q (new_AGEMA_signal_11946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6913 ( .C (clk), .D (new_AGEMA_signal_3401), .Q (new_AGEMA_signal_11950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6917 ( .C (clk), .D (RoundReg_Inst_ff_SDE_42_next_state), .Q (new_AGEMA_signal_11954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6921 ( .C (clk), .D (new_AGEMA_signal_3404), .Q (new_AGEMA_signal_11958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6925 ( .C (clk), .D (new_AGEMA_signal_3405), .Q (new_AGEMA_signal_11962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6929 ( .C (clk), .D (RoundReg_Inst_ff_SDE_43_next_state), .Q (new_AGEMA_signal_11966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6933 ( .C (clk), .D (new_AGEMA_signal_3408), .Q (new_AGEMA_signal_11970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6937 ( .C (clk), .D (new_AGEMA_signal_3409), .Q (new_AGEMA_signal_11974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6941 ( .C (clk), .D (RoundReg_Inst_ff_SDE_44_next_state), .Q (new_AGEMA_signal_11978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6945 ( .C (clk), .D (new_AGEMA_signal_3412), .Q (new_AGEMA_signal_11982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6949 ( .C (clk), .D (new_AGEMA_signal_3413), .Q (new_AGEMA_signal_11986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6953 ( .C (clk), .D (RoundReg_Inst_ff_SDE_45_next_state), .Q (new_AGEMA_signal_11990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6957 ( .C (clk), .D (new_AGEMA_signal_3416), .Q (new_AGEMA_signal_11994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6961 ( .C (clk), .D (new_AGEMA_signal_3417), .Q (new_AGEMA_signal_11998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6965 ( .C (clk), .D (RoundReg_Inst_ff_SDE_46_next_state), .Q (new_AGEMA_signal_12002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6969 ( .C (clk), .D (new_AGEMA_signal_3420), .Q (new_AGEMA_signal_12006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6973 ( .C (clk), .D (new_AGEMA_signal_3421), .Q (new_AGEMA_signal_12010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6977 ( .C (clk), .D (RoundReg_Inst_ff_SDE_47_next_state), .Q (new_AGEMA_signal_12014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6981 ( .C (clk), .D (new_AGEMA_signal_3424), .Q (new_AGEMA_signal_12018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6985 ( .C (clk), .D (new_AGEMA_signal_3425), .Q (new_AGEMA_signal_12022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6989 ( .C (clk), .D (RoundReg_Inst_ff_SDE_48_next_state), .Q (new_AGEMA_signal_12026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6993 ( .C (clk), .D (new_AGEMA_signal_3428), .Q (new_AGEMA_signal_12030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6997 ( .C (clk), .D (new_AGEMA_signal_3429), .Q (new_AGEMA_signal_12034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7001 ( .C (clk), .D (RoundReg_Inst_ff_SDE_49_next_state), .Q (new_AGEMA_signal_12038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7005 ( .C (clk), .D (new_AGEMA_signal_3432), .Q (new_AGEMA_signal_12042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7009 ( .C (clk), .D (new_AGEMA_signal_3433), .Q (new_AGEMA_signal_12046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7013 ( .C (clk), .D (RoundReg_Inst_ff_SDE_50_next_state), .Q (new_AGEMA_signal_12050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7017 ( .C (clk), .D (new_AGEMA_signal_3436), .Q (new_AGEMA_signal_12054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7021 ( .C (clk), .D (new_AGEMA_signal_3437), .Q (new_AGEMA_signal_12058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7025 ( .C (clk), .D (RoundReg_Inst_ff_SDE_51_next_state), .Q (new_AGEMA_signal_12062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7029 ( .C (clk), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_12066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7033 ( .C (clk), .D (new_AGEMA_signal_3441), .Q (new_AGEMA_signal_12070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7037 ( .C (clk), .D (RoundReg_Inst_ff_SDE_52_next_state), .Q (new_AGEMA_signal_12074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7041 ( .C (clk), .D (new_AGEMA_signal_3444), .Q (new_AGEMA_signal_12078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7045 ( .C (clk), .D (new_AGEMA_signal_3445), .Q (new_AGEMA_signal_12082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7049 ( .C (clk), .D (RoundReg_Inst_ff_SDE_53_next_state), .Q (new_AGEMA_signal_12086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7053 ( .C (clk), .D (new_AGEMA_signal_3448), .Q (new_AGEMA_signal_12090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7057 ( .C (clk), .D (new_AGEMA_signal_3449), .Q (new_AGEMA_signal_12094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7061 ( .C (clk), .D (RoundReg_Inst_ff_SDE_54_next_state), .Q (new_AGEMA_signal_12098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7065 ( .C (clk), .D (new_AGEMA_signal_3452), .Q (new_AGEMA_signal_12102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7069 ( .C (clk), .D (new_AGEMA_signal_3453), .Q (new_AGEMA_signal_12106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7073 ( .C (clk), .D (RoundReg_Inst_ff_SDE_55_next_state), .Q (new_AGEMA_signal_12110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7077 ( .C (clk), .D (new_AGEMA_signal_3456), .Q (new_AGEMA_signal_12114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7081 ( .C (clk), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_12118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7085 ( .C (clk), .D (RoundReg_Inst_ff_SDE_56_next_state), .Q (new_AGEMA_signal_12122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7089 ( .C (clk), .D (new_AGEMA_signal_3460), .Q (new_AGEMA_signal_12126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7093 ( .C (clk), .D (new_AGEMA_signal_3461), .Q (new_AGEMA_signal_12130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7097 ( .C (clk), .D (RoundReg_Inst_ff_SDE_57_next_state), .Q (new_AGEMA_signal_12134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7101 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_12138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7105 ( .C (clk), .D (new_AGEMA_signal_3465), .Q (new_AGEMA_signal_12142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7109 ( .C (clk), .D (RoundReg_Inst_ff_SDE_58_next_state), .Q (new_AGEMA_signal_12146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7113 ( .C (clk), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_12150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7117 ( .C (clk), .D (new_AGEMA_signal_3469), .Q (new_AGEMA_signal_12154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7121 ( .C (clk), .D (RoundReg_Inst_ff_SDE_59_next_state), .Q (new_AGEMA_signal_12158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7125 ( .C (clk), .D (new_AGEMA_signal_3472), .Q (new_AGEMA_signal_12162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7129 ( .C (clk), .D (new_AGEMA_signal_3473), .Q (new_AGEMA_signal_12166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7133 ( .C (clk), .D (RoundReg_Inst_ff_SDE_60_next_state), .Q (new_AGEMA_signal_12170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7137 ( .C (clk), .D (new_AGEMA_signal_3476), .Q (new_AGEMA_signal_12174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7141 ( .C (clk), .D (new_AGEMA_signal_3477), .Q (new_AGEMA_signal_12178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7145 ( .C (clk), .D (RoundReg_Inst_ff_SDE_61_next_state), .Q (new_AGEMA_signal_12182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7149 ( .C (clk), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_12186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7153 ( .C (clk), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_12190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7157 ( .C (clk), .D (RoundReg_Inst_ff_SDE_62_next_state), .Q (new_AGEMA_signal_12194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7161 ( .C (clk), .D (new_AGEMA_signal_3484), .Q (new_AGEMA_signal_12198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7165 ( .C (clk), .D (new_AGEMA_signal_3485), .Q (new_AGEMA_signal_12202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7169 ( .C (clk), .D (RoundReg_Inst_ff_SDE_63_next_state), .Q (new_AGEMA_signal_12206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7173 ( .C (clk), .D (new_AGEMA_signal_3488), .Q (new_AGEMA_signal_12210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7177 ( .C (clk), .D (new_AGEMA_signal_3489), .Q (new_AGEMA_signal_12214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7181 ( .C (clk), .D (RoundReg_Inst_ff_SDE_64_next_state), .Q (new_AGEMA_signal_12218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7185 ( .C (clk), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_12222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7189 ( .C (clk), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_12226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7193 ( .C (clk), .D (RoundReg_Inst_ff_SDE_65_next_state), .Q (new_AGEMA_signal_12230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7197 ( .C (clk), .D (new_AGEMA_signal_3496), .Q (new_AGEMA_signal_12234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7201 ( .C (clk), .D (new_AGEMA_signal_3497), .Q (new_AGEMA_signal_12238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7205 ( .C (clk), .D (RoundReg_Inst_ff_SDE_66_next_state), .Q (new_AGEMA_signal_12242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7209 ( .C (clk), .D (new_AGEMA_signal_3500), .Q (new_AGEMA_signal_12246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7213 ( .C (clk), .D (new_AGEMA_signal_3501), .Q (new_AGEMA_signal_12250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7217 ( .C (clk), .D (RoundReg_Inst_ff_SDE_67_next_state), .Q (new_AGEMA_signal_12254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7221 ( .C (clk), .D (new_AGEMA_signal_3504), .Q (new_AGEMA_signal_12258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7225 ( .C (clk), .D (new_AGEMA_signal_3505), .Q (new_AGEMA_signal_12262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7229 ( .C (clk), .D (RoundReg_Inst_ff_SDE_68_next_state), .Q (new_AGEMA_signal_12266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7233 ( .C (clk), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_12270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7237 ( .C (clk), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_12274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7241 ( .C (clk), .D (RoundReg_Inst_ff_SDE_69_next_state), .Q (new_AGEMA_signal_12278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7245 ( .C (clk), .D (new_AGEMA_signal_3512), .Q (new_AGEMA_signal_12282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7249 ( .C (clk), .D (new_AGEMA_signal_3513), .Q (new_AGEMA_signal_12286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7253 ( .C (clk), .D (RoundReg_Inst_ff_SDE_70_next_state), .Q (new_AGEMA_signal_12290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7257 ( .C (clk), .D (new_AGEMA_signal_3516), .Q (new_AGEMA_signal_12294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7261 ( .C (clk), .D (new_AGEMA_signal_3517), .Q (new_AGEMA_signal_12298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7265 ( .C (clk), .D (RoundReg_Inst_ff_SDE_71_next_state), .Q (new_AGEMA_signal_12302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7269 ( .C (clk), .D (new_AGEMA_signal_3520), .Q (new_AGEMA_signal_12306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7273 ( .C (clk), .D (new_AGEMA_signal_3521), .Q (new_AGEMA_signal_12310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7277 ( .C (clk), .D (RoundReg_Inst_ff_SDE_72_next_state), .Q (new_AGEMA_signal_12314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7281 ( .C (clk), .D (new_AGEMA_signal_3524), .Q (new_AGEMA_signal_12318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7285 ( .C (clk), .D (new_AGEMA_signal_3525), .Q (new_AGEMA_signal_12322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7289 ( .C (clk), .D (RoundReg_Inst_ff_SDE_73_next_state), .Q (new_AGEMA_signal_12326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7293 ( .C (clk), .D (new_AGEMA_signal_3528), .Q (new_AGEMA_signal_12330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7297 ( .C (clk), .D (new_AGEMA_signal_3529), .Q (new_AGEMA_signal_12334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7301 ( .C (clk), .D (RoundReg_Inst_ff_SDE_74_next_state), .Q (new_AGEMA_signal_12338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7305 ( .C (clk), .D (new_AGEMA_signal_3532), .Q (new_AGEMA_signal_12342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7309 ( .C (clk), .D (new_AGEMA_signal_3533), .Q (new_AGEMA_signal_12346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7313 ( .C (clk), .D (RoundReg_Inst_ff_SDE_75_next_state), .Q (new_AGEMA_signal_12350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7317 ( .C (clk), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_12354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7321 ( .C (clk), .D (new_AGEMA_signal_3537), .Q (new_AGEMA_signal_12358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7325 ( .C (clk), .D (RoundReg_Inst_ff_SDE_76_next_state), .Q (new_AGEMA_signal_12362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7329 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_12366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7333 ( .C (clk), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_12370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7337 ( .C (clk), .D (RoundReg_Inst_ff_SDE_77_next_state), .Q (new_AGEMA_signal_12374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7341 ( .C (clk), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_12378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7345 ( .C (clk), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_12382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7349 ( .C (clk), .D (RoundReg_Inst_ff_SDE_78_next_state), .Q (new_AGEMA_signal_12386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7353 ( .C (clk), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_12390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7357 ( .C (clk), .D (new_AGEMA_signal_3549), .Q (new_AGEMA_signal_12394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7361 ( .C (clk), .D (RoundReg_Inst_ff_SDE_79_next_state), .Q (new_AGEMA_signal_12398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7365 ( .C (clk), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_12402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7369 ( .C (clk), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_12406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7373 ( .C (clk), .D (RoundReg_Inst_ff_SDE_80_next_state), .Q (new_AGEMA_signal_12410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7377 ( .C (clk), .D (new_AGEMA_signal_3556), .Q (new_AGEMA_signal_12414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7381 ( .C (clk), .D (new_AGEMA_signal_3557), .Q (new_AGEMA_signal_12418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7385 ( .C (clk), .D (RoundReg_Inst_ff_SDE_81_next_state), .Q (new_AGEMA_signal_12422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7389 ( .C (clk), .D (new_AGEMA_signal_3560), .Q (new_AGEMA_signal_12426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7393 ( .C (clk), .D (new_AGEMA_signal_3561), .Q (new_AGEMA_signal_12430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7397 ( .C (clk), .D (RoundReg_Inst_ff_SDE_82_next_state), .Q (new_AGEMA_signal_12434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7401 ( .C (clk), .D (new_AGEMA_signal_3564), .Q (new_AGEMA_signal_12438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7405 ( .C (clk), .D (new_AGEMA_signal_3565), .Q (new_AGEMA_signal_12442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7409 ( .C (clk), .D (RoundReg_Inst_ff_SDE_83_next_state), .Q (new_AGEMA_signal_12446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7413 ( .C (clk), .D (new_AGEMA_signal_3568), .Q (new_AGEMA_signal_12450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7417 ( .C (clk), .D (new_AGEMA_signal_3569), .Q (new_AGEMA_signal_12454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7421 ( .C (clk), .D (RoundReg_Inst_ff_SDE_84_next_state), .Q (new_AGEMA_signal_12458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7425 ( .C (clk), .D (new_AGEMA_signal_3572), .Q (new_AGEMA_signal_12462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7429 ( .C (clk), .D (new_AGEMA_signal_3573), .Q (new_AGEMA_signal_12466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7433 ( .C (clk), .D (RoundReg_Inst_ff_SDE_85_next_state), .Q (new_AGEMA_signal_12470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7437 ( .C (clk), .D (new_AGEMA_signal_3576), .Q (new_AGEMA_signal_12474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7441 ( .C (clk), .D (new_AGEMA_signal_3577), .Q (new_AGEMA_signal_12478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7445 ( .C (clk), .D (RoundReg_Inst_ff_SDE_86_next_state), .Q (new_AGEMA_signal_12482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7449 ( .C (clk), .D (new_AGEMA_signal_3580), .Q (new_AGEMA_signal_12486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7453 ( .C (clk), .D (new_AGEMA_signal_3581), .Q (new_AGEMA_signal_12490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7457 ( .C (clk), .D (RoundReg_Inst_ff_SDE_87_next_state), .Q (new_AGEMA_signal_12494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7461 ( .C (clk), .D (new_AGEMA_signal_3584), .Q (new_AGEMA_signal_12498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7465 ( .C (clk), .D (new_AGEMA_signal_3585), .Q (new_AGEMA_signal_12502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7469 ( .C (clk), .D (RoundReg_Inst_ff_SDE_88_next_state), .Q (new_AGEMA_signal_12506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7473 ( .C (clk), .D (new_AGEMA_signal_3588), .Q (new_AGEMA_signal_12510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7477 ( .C (clk), .D (new_AGEMA_signal_3589), .Q (new_AGEMA_signal_12514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7481 ( .C (clk), .D (RoundReg_Inst_ff_SDE_89_next_state), .Q (new_AGEMA_signal_12518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7485 ( .C (clk), .D (new_AGEMA_signal_3592), .Q (new_AGEMA_signal_12522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7489 ( .C (clk), .D (new_AGEMA_signal_3593), .Q (new_AGEMA_signal_12526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7493 ( .C (clk), .D (RoundReg_Inst_ff_SDE_90_next_state), .Q (new_AGEMA_signal_12530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7497 ( .C (clk), .D (new_AGEMA_signal_3596), .Q (new_AGEMA_signal_12534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7501 ( .C (clk), .D (new_AGEMA_signal_3597), .Q (new_AGEMA_signal_12538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7505 ( .C (clk), .D (RoundReg_Inst_ff_SDE_91_next_state), .Q (new_AGEMA_signal_12542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7509 ( .C (clk), .D (new_AGEMA_signal_3600), .Q (new_AGEMA_signal_12546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7513 ( .C (clk), .D (new_AGEMA_signal_3601), .Q (new_AGEMA_signal_12550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7517 ( .C (clk), .D (RoundReg_Inst_ff_SDE_92_next_state), .Q (new_AGEMA_signal_12554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7521 ( .C (clk), .D (new_AGEMA_signal_3604), .Q (new_AGEMA_signal_12558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7525 ( .C (clk), .D (new_AGEMA_signal_3605), .Q (new_AGEMA_signal_12562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7529 ( .C (clk), .D (RoundReg_Inst_ff_SDE_93_next_state), .Q (new_AGEMA_signal_12566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7533 ( .C (clk), .D (new_AGEMA_signal_3608), .Q (new_AGEMA_signal_12570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7537 ( .C (clk), .D (new_AGEMA_signal_3609), .Q (new_AGEMA_signal_12574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7541 ( .C (clk), .D (RoundReg_Inst_ff_SDE_94_next_state), .Q (new_AGEMA_signal_12578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7545 ( .C (clk), .D (new_AGEMA_signal_3612), .Q (new_AGEMA_signal_12582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7549 ( .C (clk), .D (new_AGEMA_signal_3613), .Q (new_AGEMA_signal_12586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7553 ( .C (clk), .D (RoundReg_Inst_ff_SDE_95_next_state), .Q (new_AGEMA_signal_12590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7557 ( .C (clk), .D (new_AGEMA_signal_3616), .Q (new_AGEMA_signal_12594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7561 ( .C (clk), .D (new_AGEMA_signal_3617), .Q (new_AGEMA_signal_12598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7565 ( .C (clk), .D (RoundReg_Inst_ff_SDE_96_next_state), .Q (new_AGEMA_signal_12602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7569 ( .C (clk), .D (new_AGEMA_signal_3620), .Q (new_AGEMA_signal_12606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7573 ( .C (clk), .D (new_AGEMA_signal_3621), .Q (new_AGEMA_signal_12610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7577 ( .C (clk), .D (RoundReg_Inst_ff_SDE_97_next_state), .Q (new_AGEMA_signal_12614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7581 ( .C (clk), .D (new_AGEMA_signal_3624), .Q (new_AGEMA_signal_12618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7585 ( .C (clk), .D (new_AGEMA_signal_3625), .Q (new_AGEMA_signal_12622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7589 ( .C (clk), .D (RoundReg_Inst_ff_SDE_98_next_state), .Q (new_AGEMA_signal_12626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7593 ( .C (clk), .D (new_AGEMA_signal_3628), .Q (new_AGEMA_signal_12630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7597 ( .C (clk), .D (new_AGEMA_signal_3629), .Q (new_AGEMA_signal_12634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7601 ( .C (clk), .D (RoundReg_Inst_ff_SDE_99_next_state), .Q (new_AGEMA_signal_12638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7605 ( .C (clk), .D (new_AGEMA_signal_3632), .Q (new_AGEMA_signal_12642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7609 ( .C (clk), .D (new_AGEMA_signal_3633), .Q (new_AGEMA_signal_12646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7613 ( .C (clk), .D (RoundReg_Inst_ff_SDE_100_next_state), .Q (new_AGEMA_signal_12650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7617 ( .C (clk), .D (new_AGEMA_signal_3636), .Q (new_AGEMA_signal_12654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7621 ( .C (clk), .D (new_AGEMA_signal_3637), .Q (new_AGEMA_signal_12658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7625 ( .C (clk), .D (RoundReg_Inst_ff_SDE_101_next_state), .Q (new_AGEMA_signal_12662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7629 ( .C (clk), .D (new_AGEMA_signal_3640), .Q (new_AGEMA_signal_12666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7633 ( .C (clk), .D (new_AGEMA_signal_3641), .Q (new_AGEMA_signal_12670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7637 ( .C (clk), .D (RoundReg_Inst_ff_SDE_102_next_state), .Q (new_AGEMA_signal_12674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7641 ( .C (clk), .D (new_AGEMA_signal_3644), .Q (new_AGEMA_signal_12678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7645 ( .C (clk), .D (new_AGEMA_signal_3645), .Q (new_AGEMA_signal_12682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7649 ( .C (clk), .D (RoundReg_Inst_ff_SDE_103_next_state), .Q (new_AGEMA_signal_12686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7653 ( .C (clk), .D (new_AGEMA_signal_3648), .Q (new_AGEMA_signal_12690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7657 ( .C (clk), .D (new_AGEMA_signal_3649), .Q (new_AGEMA_signal_12694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7661 ( .C (clk), .D (RoundReg_Inst_ff_SDE_104_next_state), .Q (new_AGEMA_signal_12698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7665 ( .C (clk), .D (new_AGEMA_signal_3652), .Q (new_AGEMA_signal_12702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7669 ( .C (clk), .D (new_AGEMA_signal_3653), .Q (new_AGEMA_signal_12706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7673 ( .C (clk), .D (RoundReg_Inst_ff_SDE_105_next_state), .Q (new_AGEMA_signal_12710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7677 ( .C (clk), .D (new_AGEMA_signal_3656), .Q (new_AGEMA_signal_12714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7681 ( .C (clk), .D (new_AGEMA_signal_3657), .Q (new_AGEMA_signal_12718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7685 ( .C (clk), .D (RoundReg_Inst_ff_SDE_106_next_state), .Q (new_AGEMA_signal_12722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7689 ( .C (clk), .D (new_AGEMA_signal_3660), .Q (new_AGEMA_signal_12726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7693 ( .C (clk), .D (new_AGEMA_signal_3661), .Q (new_AGEMA_signal_12730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7697 ( .C (clk), .D (RoundReg_Inst_ff_SDE_107_next_state), .Q (new_AGEMA_signal_12734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7701 ( .C (clk), .D (new_AGEMA_signal_3664), .Q (new_AGEMA_signal_12738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7705 ( .C (clk), .D (new_AGEMA_signal_3665), .Q (new_AGEMA_signal_12742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7709 ( .C (clk), .D (RoundReg_Inst_ff_SDE_108_next_state), .Q (new_AGEMA_signal_12746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7713 ( .C (clk), .D (new_AGEMA_signal_3668), .Q (new_AGEMA_signal_12750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7717 ( .C (clk), .D (new_AGEMA_signal_3669), .Q (new_AGEMA_signal_12754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7721 ( .C (clk), .D (RoundReg_Inst_ff_SDE_109_next_state), .Q (new_AGEMA_signal_12758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7725 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_12762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7729 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_12766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7733 ( .C (clk), .D (RoundReg_Inst_ff_SDE_110_next_state), .Q (new_AGEMA_signal_12770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7737 ( .C (clk), .D (new_AGEMA_signal_3676), .Q (new_AGEMA_signal_12774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7741 ( .C (clk), .D (new_AGEMA_signal_3677), .Q (new_AGEMA_signal_12778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7745 ( .C (clk), .D (RoundReg_Inst_ff_SDE_111_next_state), .Q (new_AGEMA_signal_12782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7749 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_12786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7753 ( .C (clk), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_12790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7757 ( .C (clk), .D (RoundReg_Inst_ff_SDE_112_next_state), .Q (new_AGEMA_signal_12794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7761 ( .C (clk), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_12798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7765 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_12802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7769 ( .C (clk), .D (RoundReg_Inst_ff_SDE_113_next_state), .Q (new_AGEMA_signal_12806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7773 ( .C (clk), .D (new_AGEMA_signal_3688), .Q (new_AGEMA_signal_12810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7777 ( .C (clk), .D (new_AGEMA_signal_3689), .Q (new_AGEMA_signal_12814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7781 ( .C (clk), .D (RoundReg_Inst_ff_SDE_114_next_state), .Q (new_AGEMA_signal_12818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7785 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_12822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7789 ( .C (clk), .D (new_AGEMA_signal_3693), .Q (new_AGEMA_signal_12826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7793 ( .C (clk), .D (RoundReg_Inst_ff_SDE_115_next_state), .Q (new_AGEMA_signal_12830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7797 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_12834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7801 ( .C (clk), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_12838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7805 ( .C (clk), .D (RoundReg_Inst_ff_SDE_116_next_state), .Q (new_AGEMA_signal_12842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7809 ( .C (clk), .D (new_AGEMA_signal_3700), .Q (new_AGEMA_signal_12846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7813 ( .C (clk), .D (new_AGEMA_signal_3701), .Q (new_AGEMA_signal_12850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7817 ( .C (clk), .D (RoundReg_Inst_ff_SDE_117_next_state), .Q (new_AGEMA_signal_12854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7821 ( .C (clk), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_12858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7825 ( .C (clk), .D (new_AGEMA_signal_3705), .Q (new_AGEMA_signal_12862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7829 ( .C (clk), .D (RoundReg_Inst_ff_SDE_118_next_state), .Q (new_AGEMA_signal_12866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7833 ( .C (clk), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_12870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7837 ( .C (clk), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_12874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7841 ( .C (clk), .D (RoundReg_Inst_ff_SDE_119_next_state), .Q (new_AGEMA_signal_12878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7845 ( .C (clk), .D (new_AGEMA_signal_3712), .Q (new_AGEMA_signal_12882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7849 ( .C (clk), .D (new_AGEMA_signal_3713), .Q (new_AGEMA_signal_12886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7853 ( .C (clk), .D (RoundReg_Inst_ff_SDE_120_next_state), .Q (new_AGEMA_signal_12890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7857 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_12894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7861 ( .C (clk), .D (new_AGEMA_signal_3717), .Q (new_AGEMA_signal_12898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7865 ( .C (clk), .D (RoundReg_Inst_ff_SDE_121_next_state), .Q (new_AGEMA_signal_12902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7869 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_12906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7873 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_12910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7877 ( .C (clk), .D (RoundReg_Inst_ff_SDE_122_next_state), .Q (new_AGEMA_signal_12914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7881 ( .C (clk), .D (new_AGEMA_signal_3724), .Q (new_AGEMA_signal_12918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7885 ( .C (clk), .D (new_AGEMA_signal_3725), .Q (new_AGEMA_signal_12922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7889 ( .C (clk), .D (RoundReg_Inst_ff_SDE_123_next_state), .Q (new_AGEMA_signal_12926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7893 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_12930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7897 ( .C (clk), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_12934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7901 ( .C (clk), .D (RoundReg_Inst_ff_SDE_124_next_state), .Q (new_AGEMA_signal_12938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7905 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_12942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7909 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_12946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7913 ( .C (clk), .D (RoundReg_Inst_ff_SDE_125_next_state), .Q (new_AGEMA_signal_12950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7917 ( .C (clk), .D (new_AGEMA_signal_3736), .Q (new_AGEMA_signal_12954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7921 ( .C (clk), .D (new_AGEMA_signal_3737), .Q (new_AGEMA_signal_12958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7925 ( .C (clk), .D (RoundReg_Inst_ff_SDE_126_next_state), .Q (new_AGEMA_signal_12962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7929 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_12966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7933 ( .C (clk), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_12970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7937 ( .C (clk), .D (RoundReg_Inst_ff_SDE_127_next_state), .Q (new_AGEMA_signal_12974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7941 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_12978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7945 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_12982) ) ;
    buf_clk new_AGEMA_reg_buffer_7949 ( .C (clk), .D (RoundCounterIns_n45), .Q (new_AGEMA_signal_12986) ) ;
    buf_clk new_AGEMA_reg_buffer_7953 ( .C (clk), .D (RoundCounterIns_n44), .Q (new_AGEMA_signal_12990) ) ;
    buf_clk new_AGEMA_reg_buffer_7957 ( .C (clk), .D (RoundCounterIns_n1), .Q (new_AGEMA_signal_12994) ) ;
    buf_clk new_AGEMA_reg_buffer_7961 ( .C (clk), .D (RoundCounterIns_n42), .Q (new_AGEMA_signal_12998) ) ;
    buf_clk new_AGEMA_reg_buffer_7965 ( .C (clk), .D (InRoundCounterIns_n41), .Q (new_AGEMA_signal_13002) ) ;
    buf_clk new_AGEMA_reg_buffer_7969 ( .C (clk), .D (InRoundCounterIns_n40), .Q (new_AGEMA_signal_13006) ) ;
    buf_clk new_AGEMA_reg_buffer_7973 ( .C (clk), .D (InRoundCounterIns_n39), .Q (new_AGEMA_signal_13010) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_7148, new_AGEMA_signal_7147, new_AGEMA_signal_7146}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_7151, new_AGEMA_signal_7150, new_AGEMA_signal_7149}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4175, new_AGEMA_signal_4174, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, new_AGEMA_signal_7152}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_7157, new_AGEMA_signal_7156, new_AGEMA_signal_7155}), .b ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_4219, new_AGEMA_signal_4218, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_7160, new_AGEMA_signal_7159, new_AGEMA_signal_7158}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4183, new_AGEMA_signal_4182, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_7163, new_AGEMA_signal_7162, new_AGEMA_signal_7161}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, new_AGEMA_signal_7164}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_7169, new_AGEMA_signal_7168, new_AGEMA_signal_7167}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_4229, new_AGEMA_signal_4228, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_7172, new_AGEMA_signal_7171, new_AGEMA_signal_7170}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4193, new_AGEMA_signal_4192, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_7175, new_AGEMA_signal_7174, new_AGEMA_signal_7173}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, new_AGEMA_signal_7176}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4199, new_AGEMA_signal_4198, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_7181, new_AGEMA_signal_7180, new_AGEMA_signal_7179}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_7184, new_AGEMA_signal_7183, new_AGEMA_signal_7182}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_7187, new_AGEMA_signal_7186, new_AGEMA_signal_7185}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, new_AGEMA_signal_7188}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_7193, new_AGEMA_signal_7192, new_AGEMA_signal_7191}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2109 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_7146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_4110), .Q (new_AGEMA_signal_7147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_4111), .Q (new_AGEMA_signal_7148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2112 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_7149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_4138), .Q (new_AGEMA_signal_7150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_7151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2115 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_7152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_7153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_4143), .Q (new_AGEMA_signal_7154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2118 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_7155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_4170), .Q (new_AGEMA_signal_7156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_4171), .Q (new_AGEMA_signal_7157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2121 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_7158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_7159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_4119), .Q (new_AGEMA_signal_7160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2124 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_7161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_4146), .Q (new_AGEMA_signal_7162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_4147), .Q (new_AGEMA_signal_7163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2127 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_7164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_7165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_4151), .Q (new_AGEMA_signal_7166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2130 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_7167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_7168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_4181), .Q (new_AGEMA_signal_7169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2133 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_7170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_7171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_4127), .Q (new_AGEMA_signal_7172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2136 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_7173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_7174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_4155), .Q (new_AGEMA_signal_7175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2139 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_7176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_4158), .Q (new_AGEMA_signal_7177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_7178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2142 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_7179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_7180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_4191), .Q (new_AGEMA_signal_7181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2145 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_7182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_4134), .Q (new_AGEMA_signal_7183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_4135), .Q (new_AGEMA_signal_7184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2148 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_7185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_4162), .Q (new_AGEMA_signal_7186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_4163), .Q (new_AGEMA_signal_7187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2151 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_7188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_7189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_4167), .Q (new_AGEMA_signal_7190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2154 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_7191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_4200), .Q (new_AGEMA_signal_7192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_7193) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_7242), .Q (new_AGEMA_signal_7243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_7246), .Q (new_AGEMA_signal_7247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_7250), .Q (new_AGEMA_signal_7251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_7254), .Q (new_AGEMA_signal_7255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_7258), .Q (new_AGEMA_signal_7259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_7262), .Q (new_AGEMA_signal_7263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_7266), .Q (new_AGEMA_signal_7267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_7270), .Q (new_AGEMA_signal_7271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_7274), .Q (new_AGEMA_signal_7275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_7278), .Q (new_AGEMA_signal_7279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_7282), .Q (new_AGEMA_signal_7283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_7286), .Q (new_AGEMA_signal_7287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_7290), .Q (new_AGEMA_signal_7291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_7294), .Q (new_AGEMA_signal_7295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_7298), .Q (new_AGEMA_signal_7299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_7302), .Q (new_AGEMA_signal_7303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_7306), .Q (new_AGEMA_signal_7307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_7310), .Q (new_AGEMA_signal_7311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_7314), .Q (new_AGEMA_signal_7315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_7318), .Q (new_AGEMA_signal_7319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_7322), .Q (new_AGEMA_signal_7323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_7326), .Q (new_AGEMA_signal_7327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_7330), .Q (new_AGEMA_signal_7331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_7334), .Q (new_AGEMA_signal_7335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_7338), .Q (new_AGEMA_signal_7339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_7342), .Q (new_AGEMA_signal_7343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_7346), .Q (new_AGEMA_signal_7347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_7350), .Q (new_AGEMA_signal_7351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_7354), .Q (new_AGEMA_signal_7355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_7358), .Q (new_AGEMA_signal_7359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_7362), .Q (new_AGEMA_signal_7363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_7366), .Q (new_AGEMA_signal_7367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_7370), .Q (new_AGEMA_signal_7371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_7374), .Q (new_AGEMA_signal_7375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_7378), .Q (new_AGEMA_signal_7379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_7382), .Q (new_AGEMA_signal_7383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_7386), .Q (new_AGEMA_signal_7387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_7390), .Q (new_AGEMA_signal_7391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_7394), .Q (new_AGEMA_signal_7395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_7398), .Q (new_AGEMA_signal_7399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_7402), .Q (new_AGEMA_signal_7403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_7406), .Q (new_AGEMA_signal_7407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_7410), .Q (new_AGEMA_signal_7411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_7414), .Q (new_AGEMA_signal_7415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_7418), .Q (new_AGEMA_signal_7419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_7422), .Q (new_AGEMA_signal_7423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_7426), .Q (new_AGEMA_signal_7427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_7430), .Q (new_AGEMA_signal_7431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_7434), .Q (new_AGEMA_signal_7435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_7438), .Q (new_AGEMA_signal_7439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_7442), .Q (new_AGEMA_signal_7443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_7447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_7450), .Q (new_AGEMA_signal_7451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_7454), .Q (new_AGEMA_signal_7455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_7458), .Q (new_AGEMA_signal_7459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_7462), .Q (new_AGEMA_signal_7463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_7466), .Q (new_AGEMA_signal_7467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_7470), .Q (new_AGEMA_signal_7471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_7474), .Q (new_AGEMA_signal_7475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_7478), .Q (new_AGEMA_signal_7479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_7482), .Q (new_AGEMA_signal_7483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_7487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_7490), .Q (new_AGEMA_signal_7491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_7494), .Q (new_AGEMA_signal_7495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_7498), .Q (new_AGEMA_signal_7499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_7502), .Q (new_AGEMA_signal_7503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_7506), .Q (new_AGEMA_signal_7507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_7510), .Q (new_AGEMA_signal_7511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_7514), .Q (new_AGEMA_signal_7515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_7518), .Q (new_AGEMA_signal_7519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_7522), .Q (new_AGEMA_signal_7523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_7526), .Q (new_AGEMA_signal_7527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_7530), .Q (new_AGEMA_signal_7531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_7534), .Q (new_AGEMA_signal_7535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_7538), .Q (new_AGEMA_signal_7539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_7542), .Q (new_AGEMA_signal_7543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_7546), .Q (new_AGEMA_signal_7547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_7550), .Q (new_AGEMA_signal_7551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_7554), .Q (new_AGEMA_signal_7555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_7558), .Q (new_AGEMA_signal_7559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_7562), .Q (new_AGEMA_signal_7563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_7566), .Q (new_AGEMA_signal_7567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_7570), .Q (new_AGEMA_signal_7571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_7574), .Q (new_AGEMA_signal_7575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_7578), .Q (new_AGEMA_signal_7579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_7582), .Q (new_AGEMA_signal_7583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_7586), .Q (new_AGEMA_signal_7587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_7590), .Q (new_AGEMA_signal_7591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_7594), .Q (new_AGEMA_signal_7595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_7598), .Q (new_AGEMA_signal_7599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_7602), .Q (new_AGEMA_signal_7603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_7606), .Q (new_AGEMA_signal_7607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_7610), .Q (new_AGEMA_signal_7611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_7614), .Q (new_AGEMA_signal_7615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_7618), .Q (new_AGEMA_signal_7619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_7622), .Q (new_AGEMA_signal_7623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_7626), .Q (new_AGEMA_signal_7627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_7630), .Q (new_AGEMA_signal_7631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_7633), .Q (new_AGEMA_signal_7634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_7636), .Q (new_AGEMA_signal_7637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_7639), .Q (new_AGEMA_signal_7640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_7642), .Q (new_AGEMA_signal_7643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_7645), .Q (new_AGEMA_signal_7646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_7648), .Q (new_AGEMA_signal_7649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_7651), .Q (new_AGEMA_signal_7652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_7654), .Q (new_AGEMA_signal_7655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_7657), .Q (new_AGEMA_signal_7658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_7660), .Q (new_AGEMA_signal_7661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_7663), .Q (new_AGEMA_signal_7664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_7666), .Q (new_AGEMA_signal_7667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_7669), .Q (new_AGEMA_signal_7670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_7672), .Q (new_AGEMA_signal_7673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_7675), .Q (new_AGEMA_signal_7676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_7678), .Q (new_AGEMA_signal_7679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_7681), .Q (new_AGEMA_signal_7682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_7684), .Q (new_AGEMA_signal_7685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_7687), .Q (new_AGEMA_signal_7688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_7690), .Q (new_AGEMA_signal_7691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_7693), .Q (new_AGEMA_signal_7694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_7697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_7699), .Q (new_AGEMA_signal_7700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_7702), .Q (new_AGEMA_signal_7703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_7705), .Q (new_AGEMA_signal_7706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_7708), .Q (new_AGEMA_signal_7709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_7711), .Q (new_AGEMA_signal_7712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_7714), .Q (new_AGEMA_signal_7715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_7717), .Q (new_AGEMA_signal_7718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_7720), .Q (new_AGEMA_signal_7721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_7723), .Q (new_AGEMA_signal_7724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_7726), .Q (new_AGEMA_signal_7727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_7729), .Q (new_AGEMA_signal_7730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_7732), .Q (new_AGEMA_signal_7733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_7735), .Q (new_AGEMA_signal_7736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_7738), .Q (new_AGEMA_signal_7739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_7741), .Q (new_AGEMA_signal_7742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_7744), .Q (new_AGEMA_signal_7745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_7747), .Q (new_AGEMA_signal_7748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_7750), .Q (new_AGEMA_signal_7751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_7753), .Q (new_AGEMA_signal_7754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_7756), .Q (new_AGEMA_signal_7757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_7759), .Q (new_AGEMA_signal_7760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_7762), .Q (new_AGEMA_signal_7763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_7765), .Q (new_AGEMA_signal_7766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_7768), .Q (new_AGEMA_signal_7769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_7771), .Q (new_AGEMA_signal_7772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_7774), .Q (new_AGEMA_signal_7775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_7777), .Q (new_AGEMA_signal_7778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_7780), .Q (new_AGEMA_signal_7781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_7783), .Q (new_AGEMA_signal_7784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_7786), .Q (new_AGEMA_signal_7787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_7789), .Q (new_AGEMA_signal_7790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_7792), .Q (new_AGEMA_signal_7793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_7795), .Q (new_AGEMA_signal_7796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_7798), .Q (new_AGEMA_signal_7799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_7801), .Q (new_AGEMA_signal_7802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_7804), .Q (new_AGEMA_signal_7805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_7807), .Q (new_AGEMA_signal_7808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_7810), .Q (new_AGEMA_signal_7811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_7813), .Q (new_AGEMA_signal_7814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_7816), .Q (new_AGEMA_signal_7817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_7819), .Q (new_AGEMA_signal_7820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_7822), .Q (new_AGEMA_signal_7823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_7825), .Q (new_AGEMA_signal_7826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_7828), .Q (new_AGEMA_signal_7829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_7831), .Q (new_AGEMA_signal_7832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_7834), .Q (new_AGEMA_signal_7835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_7837), .Q (new_AGEMA_signal_7838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_7840), .Q (new_AGEMA_signal_7841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_7843), .Q (new_AGEMA_signal_7844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_7846), .Q (new_AGEMA_signal_7847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2813 ( .C (clk), .D (new_AGEMA_signal_7849), .Q (new_AGEMA_signal_7850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_7852), .Q (new_AGEMA_signal_7853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_7855), .Q (new_AGEMA_signal_7856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_7858), .Q (new_AGEMA_signal_7859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2825 ( .C (clk), .D (new_AGEMA_signal_7861), .Q (new_AGEMA_signal_7862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_7864), .Q (new_AGEMA_signal_7865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_7867), .Q (new_AGEMA_signal_7868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_7870), .Q (new_AGEMA_signal_7871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2837 ( .C (clk), .D (new_AGEMA_signal_7873), .Q (new_AGEMA_signal_7874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_7876), .Q (new_AGEMA_signal_7877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_7879), .Q (new_AGEMA_signal_7880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_7882), .Q (new_AGEMA_signal_7883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2849 ( .C (clk), .D (new_AGEMA_signal_7885), .Q (new_AGEMA_signal_7886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_7888), .Q (new_AGEMA_signal_7889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_7891), .Q (new_AGEMA_signal_7892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_7894), .Q (new_AGEMA_signal_7895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2861 ( .C (clk), .D (new_AGEMA_signal_7897), .Q (new_AGEMA_signal_7898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_7900), .Q (new_AGEMA_signal_7901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_7903), .Q (new_AGEMA_signal_7904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_7906), .Q (new_AGEMA_signal_7907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2873 ( .C (clk), .D (new_AGEMA_signal_7909), .Q (new_AGEMA_signal_7910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_7912), .Q (new_AGEMA_signal_7913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_7915), .Q (new_AGEMA_signal_7916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_7918), .Q (new_AGEMA_signal_7919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2885 ( .C (clk), .D (new_AGEMA_signal_7921), .Q (new_AGEMA_signal_7922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_7924), .Q (new_AGEMA_signal_7925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_7927), .Q (new_AGEMA_signal_7928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_7930), .Q (new_AGEMA_signal_7931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2897 ( .C (clk), .D (new_AGEMA_signal_7933), .Q (new_AGEMA_signal_7934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_7936), .Q (new_AGEMA_signal_7937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_7939), .Q (new_AGEMA_signal_7940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_7942), .Q (new_AGEMA_signal_7943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2909 ( .C (clk), .D (new_AGEMA_signal_7945), .Q (new_AGEMA_signal_7946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_7948), .Q (new_AGEMA_signal_7949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_7951), .Q (new_AGEMA_signal_7952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_7954), .Q (new_AGEMA_signal_7955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2921 ( .C (clk), .D (new_AGEMA_signal_7957), .Q (new_AGEMA_signal_7958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_7960), .Q (new_AGEMA_signal_7961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_7963), .Q (new_AGEMA_signal_7964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_7966), .Q (new_AGEMA_signal_7967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2933 ( .C (clk), .D (new_AGEMA_signal_7969), .Q (new_AGEMA_signal_7970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_7972), .Q (new_AGEMA_signal_7973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_7975), .Q (new_AGEMA_signal_7976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_7978), .Q (new_AGEMA_signal_7979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2945 ( .C (clk), .D (new_AGEMA_signal_7981), .Q (new_AGEMA_signal_7982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_7984), .Q (new_AGEMA_signal_7985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_7987), .Q (new_AGEMA_signal_7988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_7990), .Q (new_AGEMA_signal_7991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_7993), .Q (new_AGEMA_signal_7994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_7996), .Q (new_AGEMA_signal_7997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_7999), .Q (new_AGEMA_signal_8000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_8002), .Q (new_AGEMA_signal_8003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2969 ( .C (clk), .D (new_AGEMA_signal_8005), .Q (new_AGEMA_signal_8006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_8008), .Q (new_AGEMA_signal_8009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_8011), .Q (new_AGEMA_signal_8012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_8014), .Q (new_AGEMA_signal_8015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_8017), .Q (new_AGEMA_signal_8018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_8020), .Q (new_AGEMA_signal_8021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_8023), .Q (new_AGEMA_signal_8024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_8026), .Q (new_AGEMA_signal_8027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2993 ( .C (clk), .D (new_AGEMA_signal_8029), .Q (new_AGEMA_signal_8030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_8032), .Q (new_AGEMA_signal_8033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_8035), .Q (new_AGEMA_signal_8036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_8038), .Q (new_AGEMA_signal_8039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_8041), .Q (new_AGEMA_signal_8042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_8044), .Q (new_AGEMA_signal_8045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_8047), .Q (new_AGEMA_signal_8048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_8050), .Q (new_AGEMA_signal_8051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_8053), .Q (new_AGEMA_signal_8054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_8056), .Q (new_AGEMA_signal_8057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_8059), .Q (new_AGEMA_signal_8060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_8062), .Q (new_AGEMA_signal_8063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_8065), .Q (new_AGEMA_signal_8066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_8068), .Q (new_AGEMA_signal_8069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_8071), .Q (new_AGEMA_signal_8072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_8074), .Q (new_AGEMA_signal_8075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_8077), .Q (new_AGEMA_signal_8078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_8080), .Q (new_AGEMA_signal_8081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_8083), .Q (new_AGEMA_signal_8084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_8086), .Q (new_AGEMA_signal_8087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_8089), .Q (new_AGEMA_signal_8090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_8092), .Q (new_AGEMA_signal_8093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_8095), .Q (new_AGEMA_signal_8096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_8098), .Q (new_AGEMA_signal_8099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_8101), .Q (new_AGEMA_signal_8102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_8104), .Q (new_AGEMA_signal_8105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_8107), .Q (new_AGEMA_signal_8108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_8110), .Q (new_AGEMA_signal_8111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_8113), .Q (new_AGEMA_signal_8114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_8116), .Q (new_AGEMA_signal_8117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_8119), .Q (new_AGEMA_signal_8120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_8122), .Q (new_AGEMA_signal_8123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_8125), .Q (new_AGEMA_signal_8126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_8128), .Q (new_AGEMA_signal_8129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_8131), .Q (new_AGEMA_signal_8132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_8134), .Q (new_AGEMA_signal_8135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_8137), .Q (new_AGEMA_signal_8138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_8140), .Q (new_AGEMA_signal_8141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_8143), .Q (new_AGEMA_signal_8144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_8146), .Q (new_AGEMA_signal_8147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_8149), .Q (new_AGEMA_signal_8150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_8152), .Q (new_AGEMA_signal_8153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_8155), .Q (new_AGEMA_signal_8156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_8158), .Q (new_AGEMA_signal_8159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_8161), .Q (new_AGEMA_signal_8162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_8164), .Q (new_AGEMA_signal_8165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_8167), .Q (new_AGEMA_signal_8168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_8170), .Q (new_AGEMA_signal_8171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_8173), .Q (new_AGEMA_signal_8174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_8176), .Q (new_AGEMA_signal_8177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_8179), .Q (new_AGEMA_signal_8180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_8182), .Q (new_AGEMA_signal_8183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_8185), .Q (new_AGEMA_signal_8186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_8188), .Q (new_AGEMA_signal_8189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_8191), .Q (new_AGEMA_signal_8192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_8194), .Q (new_AGEMA_signal_8195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_8197), .Q (new_AGEMA_signal_8198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_8200), .Q (new_AGEMA_signal_8201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_8203), .Q (new_AGEMA_signal_8204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_8206), .Q (new_AGEMA_signal_8207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_8209), .Q (new_AGEMA_signal_8210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_8212), .Q (new_AGEMA_signal_8213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_8215), .Q (new_AGEMA_signal_8216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_8218), .Q (new_AGEMA_signal_8219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_8221), .Q (new_AGEMA_signal_8222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_8224), .Q (new_AGEMA_signal_8225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_8227), .Q (new_AGEMA_signal_8228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_8230), .Q (new_AGEMA_signal_8231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_8233), .Q (new_AGEMA_signal_8234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_8236), .Q (new_AGEMA_signal_8237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_8239), .Q (new_AGEMA_signal_8240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_8242), .Q (new_AGEMA_signal_8243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_8245), .Q (new_AGEMA_signal_8246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_8248), .Q (new_AGEMA_signal_8249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_8251), .Q (new_AGEMA_signal_8252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_8254), .Q (new_AGEMA_signal_8255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_8257), .Q (new_AGEMA_signal_8258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_8260), .Q (new_AGEMA_signal_8261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_8263), .Q (new_AGEMA_signal_8264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_8266), .Q (new_AGEMA_signal_8267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_8269), .Q (new_AGEMA_signal_8270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_8272), .Q (new_AGEMA_signal_8273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_8275), .Q (new_AGEMA_signal_8276) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_8278), .Q (new_AGEMA_signal_8279) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_8282), .Q (new_AGEMA_signal_8283) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_8286), .Q (new_AGEMA_signal_8287) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_8290), .Q (new_AGEMA_signal_8291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_8294), .Q (new_AGEMA_signal_8295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_8298), .Q (new_AGEMA_signal_8299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_8302), .Q (new_AGEMA_signal_8303) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_8306), .Q (new_AGEMA_signal_8307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_8310), .Q (new_AGEMA_signal_8311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_8314), .Q (new_AGEMA_signal_8315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_8318), .Q (new_AGEMA_signal_8319) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_8322), .Q (new_AGEMA_signal_8323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_8326), .Q (new_AGEMA_signal_8327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_8330), .Q (new_AGEMA_signal_8331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_8334), .Q (new_AGEMA_signal_8335) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_8338), .Q (new_AGEMA_signal_8339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_8342), .Q (new_AGEMA_signal_8343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_8346), .Q (new_AGEMA_signal_8347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_8350), .Q (new_AGEMA_signal_8351) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_8354), .Q (new_AGEMA_signal_8355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_8358), .Q (new_AGEMA_signal_8359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_8362), .Q (new_AGEMA_signal_8363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_8366), .Q (new_AGEMA_signal_8367) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_8370), .Q (new_AGEMA_signal_8371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_8374), .Q (new_AGEMA_signal_8375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_8378), .Q (new_AGEMA_signal_8379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_8382), .Q (new_AGEMA_signal_8383) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_8386), .Q (new_AGEMA_signal_8387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_8390), .Q (new_AGEMA_signal_8391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_8394), .Q (new_AGEMA_signal_8395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_8398), .Q (new_AGEMA_signal_8399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_8402), .Q (new_AGEMA_signal_8403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_8406), .Q (new_AGEMA_signal_8407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_8410), .Q (new_AGEMA_signal_8411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_8414), .Q (new_AGEMA_signal_8415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_8418), .Q (new_AGEMA_signal_8419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_8422), .Q (new_AGEMA_signal_8423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_8426), .Q (new_AGEMA_signal_8427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_8430), .Q (new_AGEMA_signal_8431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_8434), .Q (new_AGEMA_signal_8435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_8438), .Q (new_AGEMA_signal_8439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_8442), .Q (new_AGEMA_signal_8443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_8446), .Q (new_AGEMA_signal_8447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_8450), .Q (new_AGEMA_signal_8451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_8454), .Q (new_AGEMA_signal_8455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_8458), .Q (new_AGEMA_signal_8459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_8462), .Q (new_AGEMA_signal_8463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_8466), .Q (new_AGEMA_signal_8467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_8470), .Q (new_AGEMA_signal_8471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_8474), .Q (new_AGEMA_signal_8475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_8478), .Q (new_AGEMA_signal_8479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_8482), .Q (new_AGEMA_signal_8483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_8486), .Q (new_AGEMA_signal_8487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_8490), .Q (new_AGEMA_signal_8491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_8494), .Q (new_AGEMA_signal_8495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_8498), .Q (new_AGEMA_signal_8499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_8502), .Q (new_AGEMA_signal_8503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_8506), .Q (new_AGEMA_signal_8507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_8510), .Q (new_AGEMA_signal_8511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_8514), .Q (new_AGEMA_signal_8515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_8518), .Q (new_AGEMA_signal_8519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_8522), .Q (new_AGEMA_signal_8523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_8526), .Q (new_AGEMA_signal_8527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_8530), .Q (new_AGEMA_signal_8531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_8534), .Q (new_AGEMA_signal_8535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_8538), .Q (new_AGEMA_signal_8539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_8542), .Q (new_AGEMA_signal_8543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_8546), .Q (new_AGEMA_signal_8547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_8550), .Q (new_AGEMA_signal_8551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_8554), .Q (new_AGEMA_signal_8555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_8558), .Q (new_AGEMA_signal_8559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_8562), .Q (new_AGEMA_signal_8563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_8566), .Q (new_AGEMA_signal_8567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_8570), .Q (new_AGEMA_signal_8571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_8574), .Q (new_AGEMA_signal_8575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_8578), .Q (new_AGEMA_signal_8579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_8582), .Q (new_AGEMA_signal_8583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_8586), .Q (new_AGEMA_signal_8587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_8590), .Q (new_AGEMA_signal_8591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_8594), .Q (new_AGEMA_signal_8595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_8598), .Q (new_AGEMA_signal_8599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_8602), .Q (new_AGEMA_signal_8603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_8606), .Q (new_AGEMA_signal_8607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_8610), .Q (new_AGEMA_signal_8611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_8614), .Q (new_AGEMA_signal_8615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_8618), .Q (new_AGEMA_signal_8619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_8622), .Q (new_AGEMA_signal_8623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_8626), .Q (new_AGEMA_signal_8627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_8630), .Q (new_AGEMA_signal_8631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_8634), .Q (new_AGEMA_signal_8635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_8638), .Q (new_AGEMA_signal_8639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_8642), .Q (new_AGEMA_signal_8643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_8646), .Q (new_AGEMA_signal_8647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_8650), .Q (new_AGEMA_signal_8651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_8654), .Q (new_AGEMA_signal_8655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_8658), .Q (new_AGEMA_signal_8659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_8662), .Q (new_AGEMA_signal_8663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_8666), .Q (new_AGEMA_signal_8667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_8670), .Q (new_AGEMA_signal_8671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_8674), .Q (new_AGEMA_signal_8675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_8678), .Q (new_AGEMA_signal_8679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_8682), .Q (new_AGEMA_signal_8683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_8686), .Q (new_AGEMA_signal_8687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_8690), .Q (new_AGEMA_signal_8691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_8694), .Q (new_AGEMA_signal_8695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_8698), .Q (new_AGEMA_signal_8699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_8702), .Q (new_AGEMA_signal_8703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_8706), .Q (new_AGEMA_signal_8707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_8710), .Q (new_AGEMA_signal_8711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_8714), .Q (new_AGEMA_signal_8715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_8718), .Q (new_AGEMA_signal_8719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_8722), .Q (new_AGEMA_signal_8723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_8726), .Q (new_AGEMA_signal_8727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_8730), .Q (new_AGEMA_signal_8731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_8734), .Q (new_AGEMA_signal_8735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_8738), .Q (new_AGEMA_signal_8739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_8742), .Q (new_AGEMA_signal_8743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_8746), .Q (new_AGEMA_signal_8747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_8750), .Q (new_AGEMA_signal_8751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_8754), .Q (new_AGEMA_signal_8755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_8758), .Q (new_AGEMA_signal_8759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_8762), .Q (new_AGEMA_signal_8763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_8766), .Q (new_AGEMA_signal_8767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_8770), .Q (new_AGEMA_signal_8771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_8774), .Q (new_AGEMA_signal_8775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_8778), .Q (new_AGEMA_signal_8779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_8782), .Q (new_AGEMA_signal_8783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_8786), .Q (new_AGEMA_signal_8787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_8790), .Q (new_AGEMA_signal_8791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_8794), .Q (new_AGEMA_signal_8795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_8798), .Q (new_AGEMA_signal_8799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_8802), .Q (new_AGEMA_signal_8803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_8806), .Q (new_AGEMA_signal_8807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_8810), .Q (new_AGEMA_signal_8811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_8814), .Q (new_AGEMA_signal_8815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_8818), .Q (new_AGEMA_signal_8819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_8822), .Q (new_AGEMA_signal_8823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_8826), .Q (new_AGEMA_signal_8827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_8830), .Q (new_AGEMA_signal_8831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_8834), .Q (new_AGEMA_signal_8835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_8838), .Q (new_AGEMA_signal_8839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_8842), .Q (new_AGEMA_signal_8843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_8846), .Q (new_AGEMA_signal_8847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_8850), .Q (new_AGEMA_signal_8851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_8854), .Q (new_AGEMA_signal_8855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_8858), .Q (new_AGEMA_signal_8859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_8862), .Q (new_AGEMA_signal_8863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_8866), .Q (new_AGEMA_signal_8867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_8870), .Q (new_AGEMA_signal_8871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_8874), .Q (new_AGEMA_signal_8875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_8878), .Q (new_AGEMA_signal_8879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_8882), .Q (new_AGEMA_signal_8883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_8886), .Q (new_AGEMA_signal_8887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_8890), .Q (new_AGEMA_signal_8891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_8894), .Q (new_AGEMA_signal_8895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_8898), .Q (new_AGEMA_signal_8899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_8902), .Q (new_AGEMA_signal_8903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_8906), .Q (new_AGEMA_signal_8907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_8910), .Q (new_AGEMA_signal_8911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_8914), .Q (new_AGEMA_signal_8915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_8918), .Q (new_AGEMA_signal_8919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_8922), .Q (new_AGEMA_signal_8923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_8926), .Q (new_AGEMA_signal_8927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_8930), .Q (new_AGEMA_signal_8931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_8934), .Q (new_AGEMA_signal_8935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_8938), .Q (new_AGEMA_signal_8939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_8942), .Q (new_AGEMA_signal_8943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_8946), .Q (new_AGEMA_signal_8947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_8950), .Q (new_AGEMA_signal_8951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_8954), .Q (new_AGEMA_signal_8955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_8958), .Q (new_AGEMA_signal_8959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_8962), .Q (new_AGEMA_signal_8963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_8966), .Q (new_AGEMA_signal_8967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_8970), .Q (new_AGEMA_signal_8971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_8974), .Q (new_AGEMA_signal_8975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_8978), .Q (new_AGEMA_signal_8979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_8982), .Q (new_AGEMA_signal_8983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_8986), .Q (new_AGEMA_signal_8987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_8990), .Q (new_AGEMA_signal_8991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_8994), .Q (new_AGEMA_signal_8995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_8998), .Q (new_AGEMA_signal_8999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_9002), .Q (new_AGEMA_signal_9003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_9006), .Q (new_AGEMA_signal_9007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_9010), .Q (new_AGEMA_signal_9011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_9014), .Q (new_AGEMA_signal_9015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_9018), .Q (new_AGEMA_signal_9019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_9022), .Q (new_AGEMA_signal_9023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_9026), .Q (new_AGEMA_signal_9027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_9030), .Q (new_AGEMA_signal_9031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_9034), .Q (new_AGEMA_signal_9035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_9038), .Q (new_AGEMA_signal_9039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_9042), .Q (new_AGEMA_signal_9043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_9046), .Q (new_AGEMA_signal_9047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_9050), .Q (new_AGEMA_signal_9051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_9054), .Q (new_AGEMA_signal_9055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_9058), .Q (new_AGEMA_signal_9059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_9062), .Q (new_AGEMA_signal_9063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_9066), .Q (new_AGEMA_signal_9067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_9070), .Q (new_AGEMA_signal_9071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_9074), .Q (new_AGEMA_signal_9075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_9078), .Q (new_AGEMA_signal_9079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_9082), .Q (new_AGEMA_signal_9083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_9086), .Q (new_AGEMA_signal_9087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_9090), .Q (new_AGEMA_signal_9091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_9094), .Q (new_AGEMA_signal_9095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_9098), .Q (new_AGEMA_signal_9099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_9102), .Q (new_AGEMA_signal_9103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_9106), .Q (new_AGEMA_signal_9107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_9110), .Q (new_AGEMA_signal_9111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_9114), .Q (new_AGEMA_signal_9115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_9118), .Q (new_AGEMA_signal_9119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_9122), .Q (new_AGEMA_signal_9123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_9126), .Q (new_AGEMA_signal_9127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_9130), .Q (new_AGEMA_signal_9131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_9134), .Q (new_AGEMA_signal_9135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_9138), .Q (new_AGEMA_signal_9139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_9142), .Q (new_AGEMA_signal_9143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_9146), .Q (new_AGEMA_signal_9147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_9150), .Q (new_AGEMA_signal_9151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_9154), .Q (new_AGEMA_signal_9155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_9158), .Q (new_AGEMA_signal_9159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_9162), .Q (new_AGEMA_signal_9163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_9166), .Q (new_AGEMA_signal_9167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_9170), .Q (new_AGEMA_signal_9171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_9174), .Q (new_AGEMA_signal_9175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_9178), .Q (new_AGEMA_signal_9179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_9182), .Q (new_AGEMA_signal_9183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_9186), .Q (new_AGEMA_signal_9187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_9190), .Q (new_AGEMA_signal_9191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_9194), .Q (new_AGEMA_signal_9195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_9198), .Q (new_AGEMA_signal_9199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_9202), .Q (new_AGEMA_signal_9203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_9206), .Q (new_AGEMA_signal_9207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_9210), .Q (new_AGEMA_signal_9211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_9214), .Q (new_AGEMA_signal_9215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_9218), .Q (new_AGEMA_signal_9219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_9222), .Q (new_AGEMA_signal_9223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_9226), .Q (new_AGEMA_signal_9227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_9230), .Q (new_AGEMA_signal_9231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_9234), .Q (new_AGEMA_signal_9235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_9238), .Q (new_AGEMA_signal_9239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_9242), .Q (new_AGEMA_signal_9243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_9246), .Q (new_AGEMA_signal_9247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_9250), .Q (new_AGEMA_signal_9251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_9254), .Q (new_AGEMA_signal_9255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_9258), .Q (new_AGEMA_signal_9259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_9262), .Q (new_AGEMA_signal_9263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_9266), .Q (new_AGEMA_signal_9267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_9270), .Q (new_AGEMA_signal_9271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_9274), .Q (new_AGEMA_signal_9275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_9278), .Q (new_AGEMA_signal_9279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_9282), .Q (new_AGEMA_signal_9283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_9286), .Q (new_AGEMA_signal_9287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_9290), .Q (new_AGEMA_signal_9291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_9294), .Q (new_AGEMA_signal_9295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_9298), .Q (new_AGEMA_signal_9299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_9302), .Q (new_AGEMA_signal_9303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_9306), .Q (new_AGEMA_signal_9307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_9310), .Q (new_AGEMA_signal_9311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_9314), .Q (new_AGEMA_signal_9315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_9318), .Q (new_AGEMA_signal_9319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_9322), .Q (new_AGEMA_signal_9323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_9326), .Q (new_AGEMA_signal_9327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_9330), .Q (new_AGEMA_signal_9331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_9334), .Q (new_AGEMA_signal_9335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_9338), .Q (new_AGEMA_signal_9339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_9342), .Q (new_AGEMA_signal_9343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_9346), .Q (new_AGEMA_signal_9347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_9350), .Q (new_AGEMA_signal_9351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_9354), .Q (new_AGEMA_signal_9355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_9358), .Q (new_AGEMA_signal_9359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_9362), .Q (new_AGEMA_signal_9363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_9366), .Q (new_AGEMA_signal_9367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_9370), .Q (new_AGEMA_signal_9371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_9374), .Q (new_AGEMA_signal_9375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_9378), .Q (new_AGEMA_signal_9379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_9382), .Q (new_AGEMA_signal_9383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_9386), .Q (new_AGEMA_signal_9387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_9390), .Q (new_AGEMA_signal_9391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_9394), .Q (new_AGEMA_signal_9395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_9398), .Q (new_AGEMA_signal_9399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_9402), .Q (new_AGEMA_signal_9403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_9406), .Q (new_AGEMA_signal_9407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_9410), .Q (new_AGEMA_signal_9411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_9414), .Q (new_AGEMA_signal_9415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_9418), .Q (new_AGEMA_signal_9419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_9422), .Q (new_AGEMA_signal_9423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_9426), .Q (new_AGEMA_signal_9427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_9430), .Q (new_AGEMA_signal_9431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_9434), .Q (new_AGEMA_signal_9435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_9438), .Q (new_AGEMA_signal_9439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_9442), .Q (new_AGEMA_signal_9443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_9446), .Q (new_AGEMA_signal_9447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_9450), .Q (new_AGEMA_signal_9451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_9454), .Q (new_AGEMA_signal_9455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_9458), .Q (new_AGEMA_signal_9459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_9462), .Q (new_AGEMA_signal_9463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_9466), .Q (new_AGEMA_signal_9467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_9470), .Q (new_AGEMA_signal_9471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_9474), .Q (new_AGEMA_signal_9475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_9478), .Q (new_AGEMA_signal_9479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_9482), .Q (new_AGEMA_signal_9483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_9486), .Q (new_AGEMA_signal_9487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_9490), .Q (new_AGEMA_signal_9491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_9494), .Q (new_AGEMA_signal_9495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_9498), .Q (new_AGEMA_signal_9499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_9502), .Q (new_AGEMA_signal_9503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_9506), .Q (new_AGEMA_signal_9507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_9510), .Q (new_AGEMA_signal_9511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_9514), .Q (new_AGEMA_signal_9515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_9518), .Q (new_AGEMA_signal_9519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_9522), .Q (new_AGEMA_signal_9523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_9526), .Q (new_AGEMA_signal_9527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_9530), .Q (new_AGEMA_signal_9531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_9534), .Q (new_AGEMA_signal_9535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_9538), .Q (new_AGEMA_signal_9539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_9542), .Q (new_AGEMA_signal_9543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_9546), .Q (new_AGEMA_signal_9547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_9550), .Q (new_AGEMA_signal_9551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_9554), .Q (new_AGEMA_signal_9555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_9558), .Q (new_AGEMA_signal_9559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_9562), .Q (new_AGEMA_signal_9563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_9566), .Q (new_AGEMA_signal_9567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_9570), .Q (new_AGEMA_signal_9571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_9574), .Q (new_AGEMA_signal_9575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_9578), .Q (new_AGEMA_signal_9579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_9582), .Q (new_AGEMA_signal_9583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_9586), .Q (new_AGEMA_signal_9587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_9590), .Q (new_AGEMA_signal_9591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_9594), .Q (new_AGEMA_signal_9595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_9598), .Q (new_AGEMA_signal_9599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_9602), .Q (new_AGEMA_signal_9603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_9606), .Q (new_AGEMA_signal_9607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_9610), .Q (new_AGEMA_signal_9611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_9614), .Q (new_AGEMA_signal_9615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_9618), .Q (new_AGEMA_signal_9619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_9622), .Q (new_AGEMA_signal_9623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_9626), .Q (new_AGEMA_signal_9627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_9630), .Q (new_AGEMA_signal_9631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_9634), .Q (new_AGEMA_signal_9635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_9638), .Q (new_AGEMA_signal_9639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_9642), .Q (new_AGEMA_signal_9643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_9646), .Q (new_AGEMA_signal_9647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_9650), .Q (new_AGEMA_signal_9651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_9654), .Q (new_AGEMA_signal_9655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_9658), .Q (new_AGEMA_signal_9659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_9662), .Q (new_AGEMA_signal_9663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_9666), .Q (new_AGEMA_signal_9667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_9670), .Q (new_AGEMA_signal_9671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_9674), .Q (new_AGEMA_signal_9675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_9678), .Q (new_AGEMA_signal_9679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_9682), .Q (new_AGEMA_signal_9683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_9686), .Q (new_AGEMA_signal_9687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_9690), .Q (new_AGEMA_signal_9691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_9694), .Q (new_AGEMA_signal_9695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_9698), .Q (new_AGEMA_signal_9699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_9702), .Q (new_AGEMA_signal_9703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_9706), .Q (new_AGEMA_signal_9707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_9710), .Q (new_AGEMA_signal_9711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_9714), .Q (new_AGEMA_signal_9715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_9718), .Q (new_AGEMA_signal_9719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_9722), .Q (new_AGEMA_signal_9723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_9726), .Q (new_AGEMA_signal_9727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_9730), .Q (new_AGEMA_signal_9731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_9734), .Q (new_AGEMA_signal_9735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_9738), .Q (new_AGEMA_signal_9739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_9742), .Q (new_AGEMA_signal_9743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_9746), .Q (new_AGEMA_signal_9747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_9750), .Q (new_AGEMA_signal_9751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_9754), .Q (new_AGEMA_signal_9755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_9758), .Q (new_AGEMA_signal_9759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_9762), .Q (new_AGEMA_signal_9763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_9766), .Q (new_AGEMA_signal_9767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_9770), .Q (new_AGEMA_signal_9771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_9774), .Q (new_AGEMA_signal_9775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_9778), .Q (new_AGEMA_signal_9779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_9782), .Q (new_AGEMA_signal_9783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_9786), .Q (new_AGEMA_signal_9787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_9790), .Q (new_AGEMA_signal_9791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_9794), .Q (new_AGEMA_signal_9795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_9798), .Q (new_AGEMA_signal_9799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_9802), .Q (new_AGEMA_signal_9803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_9806), .Q (new_AGEMA_signal_9807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_9810), .Q (new_AGEMA_signal_9811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_9814), .Q (new_AGEMA_signal_9815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_9818), .Q (new_AGEMA_signal_9819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_9822), .Q (new_AGEMA_signal_9823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_9826), .Q (new_AGEMA_signal_9827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_9830), .Q (new_AGEMA_signal_9831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_9834), .Q (new_AGEMA_signal_9835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_9838), .Q (new_AGEMA_signal_9839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_9842), .Q (new_AGEMA_signal_9843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_9846), .Q (new_AGEMA_signal_9847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_9850), .Q (new_AGEMA_signal_9851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_9854), .Q (new_AGEMA_signal_9855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_9858), .Q (new_AGEMA_signal_9859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_9862), .Q (new_AGEMA_signal_9863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_9866), .Q (new_AGEMA_signal_9867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_9870), .Q (new_AGEMA_signal_9871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_9874), .Q (new_AGEMA_signal_9875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_9878), .Q (new_AGEMA_signal_9879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_9882), .Q (new_AGEMA_signal_9883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_9886), .Q (new_AGEMA_signal_9887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_9890), .Q (new_AGEMA_signal_9891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_9894), .Q (new_AGEMA_signal_9895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_9898), .Q (new_AGEMA_signal_9899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_9902), .Q (new_AGEMA_signal_9903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_9906), .Q (new_AGEMA_signal_9907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_9910), .Q (new_AGEMA_signal_9911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_9914), .Q (new_AGEMA_signal_9915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_9918), .Q (new_AGEMA_signal_9919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_9922), .Q (new_AGEMA_signal_9923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_9926), .Q (new_AGEMA_signal_9927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_9930), .Q (new_AGEMA_signal_9931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_9934), .Q (new_AGEMA_signal_9935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4902 ( .C (clk), .D (new_AGEMA_signal_9938), .Q (new_AGEMA_signal_9939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_9942), .Q (new_AGEMA_signal_9943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_9946), .Q (new_AGEMA_signal_9947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4914 ( .C (clk), .D (new_AGEMA_signal_9950), .Q (new_AGEMA_signal_9951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_9954), .Q (new_AGEMA_signal_9955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_9958), .Q (new_AGEMA_signal_9959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4926 ( .C (clk), .D (new_AGEMA_signal_9962), .Q (new_AGEMA_signal_9963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_9966), .Q (new_AGEMA_signal_9967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_9970), .Q (new_AGEMA_signal_9971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_9974), .Q (new_AGEMA_signal_9975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_9978), .Q (new_AGEMA_signal_9979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_9982), .Q (new_AGEMA_signal_9983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_9986), .Q (new_AGEMA_signal_9987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_9990), .Q (new_AGEMA_signal_9991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_9994), .Q (new_AGEMA_signal_9995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_9998), .Q (new_AGEMA_signal_9999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_10002), .Q (new_AGEMA_signal_10003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_10006), .Q (new_AGEMA_signal_10007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_10010), .Q (new_AGEMA_signal_10011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_10014), .Q (new_AGEMA_signal_10015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_10018), .Q (new_AGEMA_signal_10019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_10022), .Q (new_AGEMA_signal_10023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_10026), .Q (new_AGEMA_signal_10027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_10030), .Q (new_AGEMA_signal_10031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_10034), .Q (new_AGEMA_signal_10035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_10038), .Q (new_AGEMA_signal_10039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_10042), .Q (new_AGEMA_signal_10043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_10046), .Q (new_AGEMA_signal_10047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_10050), .Q (new_AGEMA_signal_10051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_10054), .Q (new_AGEMA_signal_10055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_10058), .Q (new_AGEMA_signal_10059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_10062), .Q (new_AGEMA_signal_10063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_10066), .Q (new_AGEMA_signal_10067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_10070), .Q (new_AGEMA_signal_10071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_10074), .Q (new_AGEMA_signal_10075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_10078), .Q (new_AGEMA_signal_10079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_10082), .Q (new_AGEMA_signal_10083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_10086), .Q (new_AGEMA_signal_10087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_10090), .Q (new_AGEMA_signal_10091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_10094), .Q (new_AGEMA_signal_10095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_10098), .Q (new_AGEMA_signal_10099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_10102), .Q (new_AGEMA_signal_10103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_10106), .Q (new_AGEMA_signal_10107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_10110), .Q (new_AGEMA_signal_10111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_10114), .Q (new_AGEMA_signal_10115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_10118), .Q (new_AGEMA_signal_10119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_10122), .Q (new_AGEMA_signal_10123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_10126), .Q (new_AGEMA_signal_10127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_10130), .Q (new_AGEMA_signal_10131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_10134), .Q (new_AGEMA_signal_10135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_10138), .Q (new_AGEMA_signal_10139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_10142), .Q (new_AGEMA_signal_10143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_10146), .Q (new_AGEMA_signal_10147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_10150), .Q (new_AGEMA_signal_10151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_10154), .Q (new_AGEMA_signal_10155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_10158), .Q (new_AGEMA_signal_10159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_10162), .Q (new_AGEMA_signal_10163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_10166), .Q (new_AGEMA_signal_10167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_10170), .Q (new_AGEMA_signal_10171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_10174), .Q (new_AGEMA_signal_10175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_10178), .Q (new_AGEMA_signal_10179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_10182), .Q (new_AGEMA_signal_10183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_10186), .Q (new_AGEMA_signal_10187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_10190), .Q (new_AGEMA_signal_10191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_10194), .Q (new_AGEMA_signal_10195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_10198), .Q (new_AGEMA_signal_10199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_10202), .Q (new_AGEMA_signal_10203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_10206), .Q (new_AGEMA_signal_10207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_10210), .Q (new_AGEMA_signal_10211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_10214), .Q (new_AGEMA_signal_10215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_10218), .Q (new_AGEMA_signal_10219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_10222), .Q (new_AGEMA_signal_10223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_10226), .Q (new_AGEMA_signal_10227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_10230), .Q (new_AGEMA_signal_10231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_10234), .Q (new_AGEMA_signal_10235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_10238), .Q (new_AGEMA_signal_10239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_10242), .Q (new_AGEMA_signal_10243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_10246), .Q (new_AGEMA_signal_10247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_10250), .Q (new_AGEMA_signal_10251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_10254), .Q (new_AGEMA_signal_10255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_10258), .Q (new_AGEMA_signal_10259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_10262), .Q (new_AGEMA_signal_10263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_10266), .Q (new_AGEMA_signal_10267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_10270), .Q (new_AGEMA_signal_10271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_10274), .Q (new_AGEMA_signal_10275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_10278), .Q (new_AGEMA_signal_10279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_10282), .Q (new_AGEMA_signal_10283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_10286), .Q (new_AGEMA_signal_10287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_10290), .Q (new_AGEMA_signal_10291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_10294), .Q (new_AGEMA_signal_10295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_10298), .Q (new_AGEMA_signal_10299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_10302), .Q (new_AGEMA_signal_10303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_10306), .Q (new_AGEMA_signal_10307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_10310), .Q (new_AGEMA_signal_10311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_10314), .Q (new_AGEMA_signal_10315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_10318), .Q (new_AGEMA_signal_10319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_10322), .Q (new_AGEMA_signal_10323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_10326), .Q (new_AGEMA_signal_10327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_10330), .Q (new_AGEMA_signal_10331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_10334), .Q (new_AGEMA_signal_10335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_10338), .Q (new_AGEMA_signal_10339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_10342), .Q (new_AGEMA_signal_10343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_10346), .Q (new_AGEMA_signal_10347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_10350), .Q (new_AGEMA_signal_10351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_10354), .Q (new_AGEMA_signal_10355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_10358), .Q (new_AGEMA_signal_10359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_10362), .Q (new_AGEMA_signal_10363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_10366), .Q (new_AGEMA_signal_10367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_10370), .Q (new_AGEMA_signal_10371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_10374), .Q (new_AGEMA_signal_10375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_10378), .Q (new_AGEMA_signal_10379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_10382), .Q (new_AGEMA_signal_10383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_10386), .Q (new_AGEMA_signal_10387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_10390), .Q (new_AGEMA_signal_10391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_10394), .Q (new_AGEMA_signal_10395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_10398), .Q (new_AGEMA_signal_10399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_10402), .Q (new_AGEMA_signal_10403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_10406), .Q (new_AGEMA_signal_10407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_10410), .Q (new_AGEMA_signal_10411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_10414), .Q (new_AGEMA_signal_10415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_10418), .Q (new_AGEMA_signal_10419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_10422), .Q (new_AGEMA_signal_10423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_10426), .Q (new_AGEMA_signal_10427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_10430), .Q (new_AGEMA_signal_10431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_10434), .Q (new_AGEMA_signal_10435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_10438), .Q (new_AGEMA_signal_10439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_10442), .Q (new_AGEMA_signal_10443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_10446), .Q (new_AGEMA_signal_10447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_10450), .Q (new_AGEMA_signal_10451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_10454), .Q (new_AGEMA_signal_10455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_10458), .Q (new_AGEMA_signal_10459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_10462), .Q (new_AGEMA_signal_10463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_10466), .Q (new_AGEMA_signal_10467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_10470), .Q (new_AGEMA_signal_10471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_10474), .Q (new_AGEMA_signal_10475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_10478), .Q (new_AGEMA_signal_10479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_10482), .Q (new_AGEMA_signal_10483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_10486), .Q (new_AGEMA_signal_10487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_10490), .Q (new_AGEMA_signal_10491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_10494), .Q (new_AGEMA_signal_10495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_10498), .Q (new_AGEMA_signal_10499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_10502), .Q (new_AGEMA_signal_10503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_10506), .Q (new_AGEMA_signal_10507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_10510), .Q (new_AGEMA_signal_10511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_10514), .Q (new_AGEMA_signal_10515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_10518), .Q (new_AGEMA_signal_10519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_10522), .Q (new_AGEMA_signal_10523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_10526), .Q (new_AGEMA_signal_10527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_10530), .Q (new_AGEMA_signal_10531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_10534), .Q (new_AGEMA_signal_10535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_10538), .Q (new_AGEMA_signal_10539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_10542), .Q (new_AGEMA_signal_10543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_10546), .Q (new_AGEMA_signal_10547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_10550), .Q (new_AGEMA_signal_10551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_10554), .Q (new_AGEMA_signal_10555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_10558), .Q (new_AGEMA_signal_10559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_10562), .Q (new_AGEMA_signal_10563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_10566), .Q (new_AGEMA_signal_10567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_10570), .Q (new_AGEMA_signal_10571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_10574), .Q (new_AGEMA_signal_10575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_10578), .Q (new_AGEMA_signal_10579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_10582), .Q (new_AGEMA_signal_10583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_10586), .Q (new_AGEMA_signal_10587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_10590), .Q (new_AGEMA_signal_10591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_10594), .Q (new_AGEMA_signal_10595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_10598), .Q (new_AGEMA_signal_10599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_10602), .Q (new_AGEMA_signal_10603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_10606), .Q (new_AGEMA_signal_10607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_10610), .Q (new_AGEMA_signal_10611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_10614), .Q (new_AGEMA_signal_10615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_10618), .Q (new_AGEMA_signal_10619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_10622), .Q (new_AGEMA_signal_10623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_10626), .Q (new_AGEMA_signal_10627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_10630), .Q (new_AGEMA_signal_10631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_10634), .Q (new_AGEMA_signal_10635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_10638), .Q (new_AGEMA_signal_10639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_10642), .Q (new_AGEMA_signal_10643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_10646), .Q (new_AGEMA_signal_10647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_10650), .Q (new_AGEMA_signal_10651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_10654), .Q (new_AGEMA_signal_10655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_10658), .Q (new_AGEMA_signal_10659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_10662), .Q (new_AGEMA_signal_10663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_10666), .Q (new_AGEMA_signal_10667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_10670), .Q (new_AGEMA_signal_10671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_10674), .Q (new_AGEMA_signal_10675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_10678), .Q (new_AGEMA_signal_10679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_10682), .Q (new_AGEMA_signal_10683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_10686), .Q (new_AGEMA_signal_10687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_10690), .Q (new_AGEMA_signal_10691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_10694), .Q (new_AGEMA_signal_10695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_10698), .Q (new_AGEMA_signal_10699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_10702), .Q (new_AGEMA_signal_10703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_10706), .Q (new_AGEMA_signal_10707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_10710), .Q (new_AGEMA_signal_10711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_10714), .Q (new_AGEMA_signal_10715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_10718), .Q (new_AGEMA_signal_10719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_10722), .Q (new_AGEMA_signal_10723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_10726), .Q (new_AGEMA_signal_10727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_10730), .Q (new_AGEMA_signal_10731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_10734), .Q (new_AGEMA_signal_10735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_10738), .Q (new_AGEMA_signal_10739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_10742), .Q (new_AGEMA_signal_10743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_10746), .Q (new_AGEMA_signal_10747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_10750), .Q (new_AGEMA_signal_10751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_10754), .Q (new_AGEMA_signal_10755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_10758), .Q (new_AGEMA_signal_10759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_10762), .Q (new_AGEMA_signal_10763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_10766), .Q (new_AGEMA_signal_10767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_10770), .Q (new_AGEMA_signal_10771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_10774), .Q (new_AGEMA_signal_10775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_10778), .Q (new_AGEMA_signal_10779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_10782), .Q (new_AGEMA_signal_10783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_10786), .Q (new_AGEMA_signal_10787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_10790), .Q (new_AGEMA_signal_10791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_10794), .Q (new_AGEMA_signal_10795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_10798), .Q (new_AGEMA_signal_10799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_10802), .Q (new_AGEMA_signal_10803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_10806), .Q (new_AGEMA_signal_10807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_10810), .Q (new_AGEMA_signal_10811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_10814), .Q (new_AGEMA_signal_10815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_10818), .Q (new_AGEMA_signal_10819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_10822), .Q (new_AGEMA_signal_10823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_10826), .Q (new_AGEMA_signal_10827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_10830), .Q (new_AGEMA_signal_10831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_10834), .Q (new_AGEMA_signal_10835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_10838), .Q (new_AGEMA_signal_10839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_10842), .Q (new_AGEMA_signal_10843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_10846), .Q (new_AGEMA_signal_10847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_10850), .Q (new_AGEMA_signal_10851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_10854), .Q (new_AGEMA_signal_10855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_10858), .Q (new_AGEMA_signal_10859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_10862), .Q (new_AGEMA_signal_10863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_10866), .Q (new_AGEMA_signal_10867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_10870), .Q (new_AGEMA_signal_10871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_10874), .Q (new_AGEMA_signal_10875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_10878), .Q (new_AGEMA_signal_10879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_10882), .Q (new_AGEMA_signal_10883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_10886), .Q (new_AGEMA_signal_10887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_10890), .Q (new_AGEMA_signal_10891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_10894), .Q (new_AGEMA_signal_10895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_10898), .Q (new_AGEMA_signal_10899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_10902), .Q (new_AGEMA_signal_10903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_10906), .Q (new_AGEMA_signal_10907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_10910), .Q (new_AGEMA_signal_10911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_10914), .Q (new_AGEMA_signal_10915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_10918), .Q (new_AGEMA_signal_10919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_10922), .Q (new_AGEMA_signal_10923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_10926), .Q (new_AGEMA_signal_10927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_10930), .Q (new_AGEMA_signal_10931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_10934), .Q (new_AGEMA_signal_10935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_10938), .Q (new_AGEMA_signal_10939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_10942), .Q (new_AGEMA_signal_10943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_10946), .Q (new_AGEMA_signal_10947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_10950), .Q (new_AGEMA_signal_10951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_10954), .Q (new_AGEMA_signal_10955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_10958), .Q (new_AGEMA_signal_10959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_10962), .Q (new_AGEMA_signal_10963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_10966), .Q (new_AGEMA_signal_10967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_10970), .Q (new_AGEMA_signal_10971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_10974), .Q (new_AGEMA_signal_10975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_10978), .Q (new_AGEMA_signal_10979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_10982), .Q (new_AGEMA_signal_10983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_10986), .Q (new_AGEMA_signal_10987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_10990), .Q (new_AGEMA_signal_10991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_10994), .Q (new_AGEMA_signal_10995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_10998), .Q (new_AGEMA_signal_10999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_11002), .Q (new_AGEMA_signal_11003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_11006), .Q (new_AGEMA_signal_11007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_11010), .Q (new_AGEMA_signal_11011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_11014), .Q (new_AGEMA_signal_11015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_11018), .Q (new_AGEMA_signal_11019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_11022), .Q (new_AGEMA_signal_11023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_11026), .Q (new_AGEMA_signal_11027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_11030), .Q (new_AGEMA_signal_11031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_11034), .Q (new_AGEMA_signal_11035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_11038), .Q (new_AGEMA_signal_11039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_11042), .Q (new_AGEMA_signal_11043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_11046), .Q (new_AGEMA_signal_11047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_11050), .Q (new_AGEMA_signal_11051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_11054), .Q (new_AGEMA_signal_11055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_11058), .Q (new_AGEMA_signal_11059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_11062), .Q (new_AGEMA_signal_11063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_11066), .Q (new_AGEMA_signal_11067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_11070), .Q (new_AGEMA_signal_11071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_11074), .Q (new_AGEMA_signal_11075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_11078), .Q (new_AGEMA_signal_11079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_11082), .Q (new_AGEMA_signal_11083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6050 ( .C (clk), .D (new_AGEMA_signal_11086), .Q (new_AGEMA_signal_11087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6054 ( .C (clk), .D (new_AGEMA_signal_11090), .Q (new_AGEMA_signal_11091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6058 ( .C (clk), .D (new_AGEMA_signal_11094), .Q (new_AGEMA_signal_11095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6062 ( .C (clk), .D (new_AGEMA_signal_11098), .Q (new_AGEMA_signal_11099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6066 ( .C (clk), .D (new_AGEMA_signal_11102), .Q (new_AGEMA_signal_11103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6070 ( .C (clk), .D (new_AGEMA_signal_11106), .Q (new_AGEMA_signal_11107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6074 ( .C (clk), .D (new_AGEMA_signal_11110), .Q (new_AGEMA_signal_11111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6078 ( .C (clk), .D (new_AGEMA_signal_11114), .Q (new_AGEMA_signal_11115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6082 ( .C (clk), .D (new_AGEMA_signal_11118), .Q (new_AGEMA_signal_11119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6086 ( .C (clk), .D (new_AGEMA_signal_11122), .Q (new_AGEMA_signal_11123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6090 ( .C (clk), .D (new_AGEMA_signal_11126), .Q (new_AGEMA_signal_11127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6094 ( .C (clk), .D (new_AGEMA_signal_11130), .Q (new_AGEMA_signal_11131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6098 ( .C (clk), .D (new_AGEMA_signal_11134), .Q (new_AGEMA_signal_11135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6102 ( .C (clk), .D (new_AGEMA_signal_11138), .Q (new_AGEMA_signal_11139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6106 ( .C (clk), .D (new_AGEMA_signal_11142), .Q (new_AGEMA_signal_11143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6110 ( .C (clk), .D (new_AGEMA_signal_11146), .Q (new_AGEMA_signal_11147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6114 ( .C (clk), .D (new_AGEMA_signal_11150), .Q (new_AGEMA_signal_11151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6118 ( .C (clk), .D (new_AGEMA_signal_11154), .Q (new_AGEMA_signal_11155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6122 ( .C (clk), .D (new_AGEMA_signal_11158), .Q (new_AGEMA_signal_11159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6126 ( .C (clk), .D (new_AGEMA_signal_11162), .Q (new_AGEMA_signal_11163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6130 ( .C (clk), .D (new_AGEMA_signal_11166), .Q (new_AGEMA_signal_11167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6134 ( .C (clk), .D (new_AGEMA_signal_11170), .Q (new_AGEMA_signal_11171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6138 ( .C (clk), .D (new_AGEMA_signal_11174), .Q (new_AGEMA_signal_11175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6142 ( .C (clk), .D (new_AGEMA_signal_11178), .Q (new_AGEMA_signal_11179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6146 ( .C (clk), .D (new_AGEMA_signal_11182), .Q (new_AGEMA_signal_11183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6150 ( .C (clk), .D (new_AGEMA_signal_11186), .Q (new_AGEMA_signal_11187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6154 ( .C (clk), .D (new_AGEMA_signal_11190), .Q (new_AGEMA_signal_11191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6158 ( .C (clk), .D (new_AGEMA_signal_11194), .Q (new_AGEMA_signal_11195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6162 ( .C (clk), .D (new_AGEMA_signal_11198), .Q (new_AGEMA_signal_11199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6166 ( .C (clk), .D (new_AGEMA_signal_11202), .Q (new_AGEMA_signal_11203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6170 ( .C (clk), .D (new_AGEMA_signal_11206), .Q (new_AGEMA_signal_11207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6174 ( .C (clk), .D (new_AGEMA_signal_11210), .Q (new_AGEMA_signal_11211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6178 ( .C (clk), .D (new_AGEMA_signal_11214), .Q (new_AGEMA_signal_11215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6182 ( .C (clk), .D (new_AGEMA_signal_11218), .Q (new_AGEMA_signal_11219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6186 ( .C (clk), .D (new_AGEMA_signal_11222), .Q (new_AGEMA_signal_11223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6190 ( .C (clk), .D (new_AGEMA_signal_11226), .Q (new_AGEMA_signal_11227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6194 ( .C (clk), .D (new_AGEMA_signal_11230), .Q (new_AGEMA_signal_11231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6198 ( .C (clk), .D (new_AGEMA_signal_11234), .Q (new_AGEMA_signal_11235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6202 ( .C (clk), .D (new_AGEMA_signal_11238), .Q (new_AGEMA_signal_11239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6206 ( .C (clk), .D (new_AGEMA_signal_11242), .Q (new_AGEMA_signal_11243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6210 ( .C (clk), .D (new_AGEMA_signal_11246), .Q (new_AGEMA_signal_11247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6214 ( .C (clk), .D (new_AGEMA_signal_11250), .Q (new_AGEMA_signal_11251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6218 ( .C (clk), .D (new_AGEMA_signal_11254), .Q (new_AGEMA_signal_11255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6222 ( .C (clk), .D (new_AGEMA_signal_11258), .Q (new_AGEMA_signal_11259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6226 ( .C (clk), .D (new_AGEMA_signal_11262), .Q (new_AGEMA_signal_11263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6230 ( .C (clk), .D (new_AGEMA_signal_11266), .Q (new_AGEMA_signal_11267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6234 ( .C (clk), .D (new_AGEMA_signal_11270), .Q (new_AGEMA_signal_11271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6238 ( .C (clk), .D (new_AGEMA_signal_11274), .Q (new_AGEMA_signal_11275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6242 ( .C (clk), .D (new_AGEMA_signal_11278), .Q (new_AGEMA_signal_11279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6246 ( .C (clk), .D (new_AGEMA_signal_11282), .Q (new_AGEMA_signal_11283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6250 ( .C (clk), .D (new_AGEMA_signal_11286), .Q (new_AGEMA_signal_11287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6254 ( .C (clk), .D (new_AGEMA_signal_11290), .Q (new_AGEMA_signal_11291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6258 ( .C (clk), .D (new_AGEMA_signal_11294), .Q (new_AGEMA_signal_11295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6262 ( .C (clk), .D (new_AGEMA_signal_11298), .Q (new_AGEMA_signal_11299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6266 ( .C (clk), .D (new_AGEMA_signal_11302), .Q (new_AGEMA_signal_11303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6270 ( .C (clk), .D (new_AGEMA_signal_11306), .Q (new_AGEMA_signal_11307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6274 ( .C (clk), .D (new_AGEMA_signal_11310), .Q (new_AGEMA_signal_11311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6278 ( .C (clk), .D (new_AGEMA_signal_11314), .Q (new_AGEMA_signal_11315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6282 ( .C (clk), .D (new_AGEMA_signal_11318), .Q (new_AGEMA_signal_11319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6286 ( .C (clk), .D (new_AGEMA_signal_11322), .Q (new_AGEMA_signal_11323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6290 ( .C (clk), .D (new_AGEMA_signal_11326), .Q (new_AGEMA_signal_11327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6294 ( .C (clk), .D (new_AGEMA_signal_11330), .Q (new_AGEMA_signal_11331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6298 ( .C (clk), .D (new_AGEMA_signal_11334), .Q (new_AGEMA_signal_11335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6302 ( .C (clk), .D (new_AGEMA_signal_11338), .Q (new_AGEMA_signal_11339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6306 ( .C (clk), .D (new_AGEMA_signal_11342), .Q (new_AGEMA_signal_11343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6310 ( .C (clk), .D (new_AGEMA_signal_11346), .Q (new_AGEMA_signal_11347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6314 ( .C (clk), .D (new_AGEMA_signal_11350), .Q (new_AGEMA_signal_11351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6318 ( .C (clk), .D (new_AGEMA_signal_11354), .Q (new_AGEMA_signal_11355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6322 ( .C (clk), .D (new_AGEMA_signal_11358), .Q (new_AGEMA_signal_11359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6326 ( .C (clk), .D (new_AGEMA_signal_11362), .Q (new_AGEMA_signal_11363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6330 ( .C (clk), .D (new_AGEMA_signal_11366), .Q (new_AGEMA_signal_11367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6334 ( .C (clk), .D (new_AGEMA_signal_11370), .Q (new_AGEMA_signal_11371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6338 ( .C (clk), .D (new_AGEMA_signal_11374), .Q (new_AGEMA_signal_11375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6342 ( .C (clk), .D (new_AGEMA_signal_11378), .Q (new_AGEMA_signal_11379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6346 ( .C (clk), .D (new_AGEMA_signal_11382), .Q (new_AGEMA_signal_11383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6350 ( .C (clk), .D (new_AGEMA_signal_11386), .Q (new_AGEMA_signal_11387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6354 ( .C (clk), .D (new_AGEMA_signal_11390), .Q (new_AGEMA_signal_11391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6358 ( .C (clk), .D (new_AGEMA_signal_11394), .Q (new_AGEMA_signal_11395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6362 ( .C (clk), .D (new_AGEMA_signal_11398), .Q (new_AGEMA_signal_11399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6366 ( .C (clk), .D (new_AGEMA_signal_11402), .Q (new_AGEMA_signal_11403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6370 ( .C (clk), .D (new_AGEMA_signal_11406), .Q (new_AGEMA_signal_11407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6374 ( .C (clk), .D (new_AGEMA_signal_11410), .Q (new_AGEMA_signal_11411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6378 ( .C (clk), .D (new_AGEMA_signal_11414), .Q (new_AGEMA_signal_11415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6382 ( .C (clk), .D (new_AGEMA_signal_11418), .Q (new_AGEMA_signal_11419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6386 ( .C (clk), .D (new_AGEMA_signal_11422), .Q (new_AGEMA_signal_11423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6390 ( .C (clk), .D (new_AGEMA_signal_11426), .Q (new_AGEMA_signal_11427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6394 ( .C (clk), .D (new_AGEMA_signal_11430), .Q (new_AGEMA_signal_11431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6398 ( .C (clk), .D (new_AGEMA_signal_11434), .Q (new_AGEMA_signal_11435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6402 ( .C (clk), .D (new_AGEMA_signal_11438), .Q (new_AGEMA_signal_11439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6406 ( .C (clk), .D (new_AGEMA_signal_11442), .Q (new_AGEMA_signal_11443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6410 ( .C (clk), .D (new_AGEMA_signal_11446), .Q (new_AGEMA_signal_11447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6414 ( .C (clk), .D (new_AGEMA_signal_11450), .Q (new_AGEMA_signal_11451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6418 ( .C (clk), .D (new_AGEMA_signal_11454), .Q (new_AGEMA_signal_11455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6422 ( .C (clk), .D (new_AGEMA_signal_11458), .Q (new_AGEMA_signal_11459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6426 ( .C (clk), .D (new_AGEMA_signal_11462), .Q (new_AGEMA_signal_11463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6430 ( .C (clk), .D (new_AGEMA_signal_11466), .Q (new_AGEMA_signal_11467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6434 ( .C (clk), .D (new_AGEMA_signal_11470), .Q (new_AGEMA_signal_11471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6438 ( .C (clk), .D (new_AGEMA_signal_11474), .Q (new_AGEMA_signal_11475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6442 ( .C (clk), .D (new_AGEMA_signal_11478), .Q (new_AGEMA_signal_11479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6446 ( .C (clk), .D (new_AGEMA_signal_11482), .Q (new_AGEMA_signal_11483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6450 ( .C (clk), .D (new_AGEMA_signal_11486), .Q (new_AGEMA_signal_11487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6454 ( .C (clk), .D (new_AGEMA_signal_11490), .Q (new_AGEMA_signal_11491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6458 ( .C (clk), .D (new_AGEMA_signal_11494), .Q (new_AGEMA_signal_11495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6462 ( .C (clk), .D (new_AGEMA_signal_11498), .Q (new_AGEMA_signal_11499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6466 ( .C (clk), .D (new_AGEMA_signal_11502), .Q (new_AGEMA_signal_11503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6470 ( .C (clk), .D (new_AGEMA_signal_11506), .Q (new_AGEMA_signal_11507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6474 ( .C (clk), .D (new_AGEMA_signal_11510), .Q (new_AGEMA_signal_11511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6478 ( .C (clk), .D (new_AGEMA_signal_11514), .Q (new_AGEMA_signal_11515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6482 ( .C (clk), .D (new_AGEMA_signal_11518), .Q (new_AGEMA_signal_11519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6486 ( .C (clk), .D (new_AGEMA_signal_11522), .Q (new_AGEMA_signal_11523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6490 ( .C (clk), .D (new_AGEMA_signal_11526), .Q (new_AGEMA_signal_11527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6494 ( .C (clk), .D (new_AGEMA_signal_11530), .Q (new_AGEMA_signal_11531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6498 ( .C (clk), .D (new_AGEMA_signal_11534), .Q (new_AGEMA_signal_11535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6502 ( .C (clk), .D (new_AGEMA_signal_11538), .Q (new_AGEMA_signal_11539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6506 ( .C (clk), .D (new_AGEMA_signal_11542), .Q (new_AGEMA_signal_11543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6510 ( .C (clk), .D (new_AGEMA_signal_11546), .Q (new_AGEMA_signal_11547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6514 ( .C (clk), .D (new_AGEMA_signal_11550), .Q (new_AGEMA_signal_11551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6518 ( .C (clk), .D (new_AGEMA_signal_11554), .Q (new_AGEMA_signal_11555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6522 ( .C (clk), .D (new_AGEMA_signal_11558), .Q (new_AGEMA_signal_11559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6526 ( .C (clk), .D (new_AGEMA_signal_11562), .Q (new_AGEMA_signal_11563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6530 ( .C (clk), .D (new_AGEMA_signal_11566), .Q (new_AGEMA_signal_11567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6534 ( .C (clk), .D (new_AGEMA_signal_11570), .Q (new_AGEMA_signal_11571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6538 ( .C (clk), .D (new_AGEMA_signal_11574), .Q (new_AGEMA_signal_11575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6542 ( .C (clk), .D (new_AGEMA_signal_11578), .Q (new_AGEMA_signal_11579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6546 ( .C (clk), .D (new_AGEMA_signal_11582), .Q (new_AGEMA_signal_11583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6550 ( .C (clk), .D (new_AGEMA_signal_11586), .Q (new_AGEMA_signal_11587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6554 ( .C (clk), .D (new_AGEMA_signal_11590), .Q (new_AGEMA_signal_11591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6558 ( .C (clk), .D (new_AGEMA_signal_11594), .Q (new_AGEMA_signal_11595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6562 ( .C (clk), .D (new_AGEMA_signal_11598), .Q (new_AGEMA_signal_11599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6566 ( .C (clk), .D (new_AGEMA_signal_11602), .Q (new_AGEMA_signal_11603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6570 ( .C (clk), .D (new_AGEMA_signal_11606), .Q (new_AGEMA_signal_11607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6574 ( .C (clk), .D (new_AGEMA_signal_11610), .Q (new_AGEMA_signal_11611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6578 ( .C (clk), .D (new_AGEMA_signal_11614), .Q (new_AGEMA_signal_11615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6582 ( .C (clk), .D (new_AGEMA_signal_11618), .Q (new_AGEMA_signal_11619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6586 ( .C (clk), .D (new_AGEMA_signal_11622), .Q (new_AGEMA_signal_11623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6590 ( .C (clk), .D (new_AGEMA_signal_11626), .Q (new_AGEMA_signal_11627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6594 ( .C (clk), .D (new_AGEMA_signal_11630), .Q (new_AGEMA_signal_11631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6598 ( .C (clk), .D (new_AGEMA_signal_11634), .Q (new_AGEMA_signal_11635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6602 ( .C (clk), .D (new_AGEMA_signal_11638), .Q (new_AGEMA_signal_11639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6606 ( .C (clk), .D (new_AGEMA_signal_11642), .Q (new_AGEMA_signal_11643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6610 ( .C (clk), .D (new_AGEMA_signal_11646), .Q (new_AGEMA_signal_11647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6614 ( .C (clk), .D (new_AGEMA_signal_11650), .Q (new_AGEMA_signal_11651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6618 ( .C (clk), .D (new_AGEMA_signal_11654), .Q (new_AGEMA_signal_11655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6622 ( .C (clk), .D (new_AGEMA_signal_11658), .Q (new_AGEMA_signal_11659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6626 ( .C (clk), .D (new_AGEMA_signal_11662), .Q (new_AGEMA_signal_11663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6630 ( .C (clk), .D (new_AGEMA_signal_11666), .Q (new_AGEMA_signal_11667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6634 ( .C (clk), .D (new_AGEMA_signal_11670), .Q (new_AGEMA_signal_11671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6638 ( .C (clk), .D (new_AGEMA_signal_11674), .Q (new_AGEMA_signal_11675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6642 ( .C (clk), .D (new_AGEMA_signal_11678), .Q (new_AGEMA_signal_11679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6646 ( .C (clk), .D (new_AGEMA_signal_11682), .Q (new_AGEMA_signal_11683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6650 ( .C (clk), .D (new_AGEMA_signal_11686), .Q (new_AGEMA_signal_11687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6654 ( .C (clk), .D (new_AGEMA_signal_11690), .Q (new_AGEMA_signal_11691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6658 ( .C (clk), .D (new_AGEMA_signal_11694), .Q (new_AGEMA_signal_11695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6662 ( .C (clk), .D (new_AGEMA_signal_11698), .Q (new_AGEMA_signal_11699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6666 ( .C (clk), .D (new_AGEMA_signal_11702), .Q (new_AGEMA_signal_11703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6670 ( .C (clk), .D (new_AGEMA_signal_11706), .Q (new_AGEMA_signal_11707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6674 ( .C (clk), .D (new_AGEMA_signal_11710), .Q (new_AGEMA_signal_11711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6678 ( .C (clk), .D (new_AGEMA_signal_11714), .Q (new_AGEMA_signal_11715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6682 ( .C (clk), .D (new_AGEMA_signal_11718), .Q (new_AGEMA_signal_11719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6686 ( .C (clk), .D (new_AGEMA_signal_11722), .Q (new_AGEMA_signal_11723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6690 ( .C (clk), .D (new_AGEMA_signal_11726), .Q (new_AGEMA_signal_11727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6694 ( .C (clk), .D (new_AGEMA_signal_11730), .Q (new_AGEMA_signal_11731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6698 ( .C (clk), .D (new_AGEMA_signal_11734), .Q (new_AGEMA_signal_11735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6702 ( .C (clk), .D (new_AGEMA_signal_11738), .Q (new_AGEMA_signal_11739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6706 ( .C (clk), .D (new_AGEMA_signal_11742), .Q (new_AGEMA_signal_11743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6710 ( .C (clk), .D (new_AGEMA_signal_11746), .Q (new_AGEMA_signal_11747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6714 ( .C (clk), .D (new_AGEMA_signal_11750), .Q (new_AGEMA_signal_11751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6718 ( .C (clk), .D (new_AGEMA_signal_11754), .Q (new_AGEMA_signal_11755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6722 ( .C (clk), .D (new_AGEMA_signal_11758), .Q (new_AGEMA_signal_11759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6726 ( .C (clk), .D (new_AGEMA_signal_11762), .Q (new_AGEMA_signal_11763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6730 ( .C (clk), .D (new_AGEMA_signal_11766), .Q (new_AGEMA_signal_11767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6734 ( .C (clk), .D (new_AGEMA_signal_11770), .Q (new_AGEMA_signal_11771) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C (clk), .D (new_AGEMA_signal_11774), .Q (new_AGEMA_signal_11775) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C (clk), .D (new_AGEMA_signal_11778), .Q (new_AGEMA_signal_11779) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C (clk), .D (new_AGEMA_signal_11782), .Q (new_AGEMA_signal_11783) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C (clk), .D (new_AGEMA_signal_11786), .Q (new_AGEMA_signal_11787) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C (clk), .D (new_AGEMA_signal_11790), .Q (new_AGEMA_signal_11791) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C (clk), .D (new_AGEMA_signal_11794), .Q (new_AGEMA_signal_11795) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C (clk), .D (new_AGEMA_signal_11798), .Q (new_AGEMA_signal_11799) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C (clk), .D (new_AGEMA_signal_11802), .Q (new_AGEMA_signal_11803) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C (clk), .D (new_AGEMA_signal_11806), .Q (new_AGEMA_signal_11807) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C (clk), .D (new_AGEMA_signal_11810), .Q (new_AGEMA_signal_11811) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C (clk), .D (new_AGEMA_signal_11814), .Q (new_AGEMA_signal_11815) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C (clk), .D (new_AGEMA_signal_11818), .Q (new_AGEMA_signal_11819) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C (clk), .D (new_AGEMA_signal_11822), .Q (new_AGEMA_signal_11823) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C (clk), .D (new_AGEMA_signal_11826), .Q (new_AGEMA_signal_11827) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C (clk), .D (new_AGEMA_signal_11830), .Q (new_AGEMA_signal_11831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6798 ( .C (clk), .D (new_AGEMA_signal_11834), .Q (new_AGEMA_signal_11835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6802 ( .C (clk), .D (new_AGEMA_signal_11838), .Q (new_AGEMA_signal_11839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6806 ( .C (clk), .D (new_AGEMA_signal_11842), .Q (new_AGEMA_signal_11843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6810 ( .C (clk), .D (new_AGEMA_signal_11846), .Q (new_AGEMA_signal_11847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6814 ( .C (clk), .D (new_AGEMA_signal_11850), .Q (new_AGEMA_signal_11851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6818 ( .C (clk), .D (new_AGEMA_signal_11854), .Q (new_AGEMA_signal_11855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6822 ( .C (clk), .D (new_AGEMA_signal_11858), .Q (new_AGEMA_signal_11859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6826 ( .C (clk), .D (new_AGEMA_signal_11862), .Q (new_AGEMA_signal_11863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6830 ( .C (clk), .D (new_AGEMA_signal_11866), .Q (new_AGEMA_signal_11867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6834 ( .C (clk), .D (new_AGEMA_signal_11870), .Q (new_AGEMA_signal_11871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6838 ( .C (clk), .D (new_AGEMA_signal_11874), .Q (new_AGEMA_signal_11875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6842 ( .C (clk), .D (new_AGEMA_signal_11878), .Q (new_AGEMA_signal_11879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6846 ( .C (clk), .D (new_AGEMA_signal_11882), .Q (new_AGEMA_signal_11883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6850 ( .C (clk), .D (new_AGEMA_signal_11886), .Q (new_AGEMA_signal_11887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6854 ( .C (clk), .D (new_AGEMA_signal_11890), .Q (new_AGEMA_signal_11891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6858 ( .C (clk), .D (new_AGEMA_signal_11894), .Q (new_AGEMA_signal_11895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6862 ( .C (clk), .D (new_AGEMA_signal_11898), .Q (new_AGEMA_signal_11899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6866 ( .C (clk), .D (new_AGEMA_signal_11902), .Q (new_AGEMA_signal_11903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6870 ( .C (clk), .D (new_AGEMA_signal_11906), .Q (new_AGEMA_signal_11907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6874 ( .C (clk), .D (new_AGEMA_signal_11910), .Q (new_AGEMA_signal_11911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6878 ( .C (clk), .D (new_AGEMA_signal_11914), .Q (new_AGEMA_signal_11915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6882 ( .C (clk), .D (new_AGEMA_signal_11918), .Q (new_AGEMA_signal_11919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6886 ( .C (clk), .D (new_AGEMA_signal_11922), .Q (new_AGEMA_signal_11923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6890 ( .C (clk), .D (new_AGEMA_signal_11926), .Q (new_AGEMA_signal_11927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6894 ( .C (clk), .D (new_AGEMA_signal_11930), .Q (new_AGEMA_signal_11931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6898 ( .C (clk), .D (new_AGEMA_signal_11934), .Q (new_AGEMA_signal_11935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6902 ( .C (clk), .D (new_AGEMA_signal_11938), .Q (new_AGEMA_signal_11939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6906 ( .C (clk), .D (new_AGEMA_signal_11942), .Q (new_AGEMA_signal_11943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6910 ( .C (clk), .D (new_AGEMA_signal_11946), .Q (new_AGEMA_signal_11947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6914 ( .C (clk), .D (new_AGEMA_signal_11950), .Q (new_AGEMA_signal_11951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6918 ( .C (clk), .D (new_AGEMA_signal_11954), .Q (new_AGEMA_signal_11955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6922 ( .C (clk), .D (new_AGEMA_signal_11958), .Q (new_AGEMA_signal_11959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6926 ( .C (clk), .D (new_AGEMA_signal_11962), .Q (new_AGEMA_signal_11963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6930 ( .C (clk), .D (new_AGEMA_signal_11966), .Q (new_AGEMA_signal_11967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6934 ( .C (clk), .D (new_AGEMA_signal_11970), .Q (new_AGEMA_signal_11971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6938 ( .C (clk), .D (new_AGEMA_signal_11974), .Q (new_AGEMA_signal_11975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6942 ( .C (clk), .D (new_AGEMA_signal_11978), .Q (new_AGEMA_signal_11979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6946 ( .C (clk), .D (new_AGEMA_signal_11982), .Q (new_AGEMA_signal_11983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6950 ( .C (clk), .D (new_AGEMA_signal_11986), .Q (new_AGEMA_signal_11987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6954 ( .C (clk), .D (new_AGEMA_signal_11990), .Q (new_AGEMA_signal_11991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6958 ( .C (clk), .D (new_AGEMA_signal_11994), .Q (new_AGEMA_signal_11995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6962 ( .C (clk), .D (new_AGEMA_signal_11998), .Q (new_AGEMA_signal_11999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6966 ( .C (clk), .D (new_AGEMA_signal_12002), .Q (new_AGEMA_signal_12003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6970 ( .C (clk), .D (new_AGEMA_signal_12006), .Q (new_AGEMA_signal_12007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6974 ( .C (clk), .D (new_AGEMA_signal_12010), .Q (new_AGEMA_signal_12011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6978 ( .C (clk), .D (new_AGEMA_signal_12014), .Q (new_AGEMA_signal_12015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6982 ( .C (clk), .D (new_AGEMA_signal_12018), .Q (new_AGEMA_signal_12019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6986 ( .C (clk), .D (new_AGEMA_signal_12022), .Q (new_AGEMA_signal_12023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6990 ( .C (clk), .D (new_AGEMA_signal_12026), .Q (new_AGEMA_signal_12027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6994 ( .C (clk), .D (new_AGEMA_signal_12030), .Q (new_AGEMA_signal_12031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6998 ( .C (clk), .D (new_AGEMA_signal_12034), .Q (new_AGEMA_signal_12035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7002 ( .C (clk), .D (new_AGEMA_signal_12038), .Q (new_AGEMA_signal_12039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7006 ( .C (clk), .D (new_AGEMA_signal_12042), .Q (new_AGEMA_signal_12043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7010 ( .C (clk), .D (new_AGEMA_signal_12046), .Q (new_AGEMA_signal_12047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7014 ( .C (clk), .D (new_AGEMA_signal_12050), .Q (new_AGEMA_signal_12051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7018 ( .C (clk), .D (new_AGEMA_signal_12054), .Q (new_AGEMA_signal_12055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7022 ( .C (clk), .D (new_AGEMA_signal_12058), .Q (new_AGEMA_signal_12059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7026 ( .C (clk), .D (new_AGEMA_signal_12062), .Q (new_AGEMA_signal_12063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7030 ( .C (clk), .D (new_AGEMA_signal_12066), .Q (new_AGEMA_signal_12067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7034 ( .C (clk), .D (new_AGEMA_signal_12070), .Q (new_AGEMA_signal_12071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7038 ( .C (clk), .D (new_AGEMA_signal_12074), .Q (new_AGEMA_signal_12075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7042 ( .C (clk), .D (new_AGEMA_signal_12078), .Q (new_AGEMA_signal_12079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7046 ( .C (clk), .D (new_AGEMA_signal_12082), .Q (new_AGEMA_signal_12083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7050 ( .C (clk), .D (new_AGEMA_signal_12086), .Q (new_AGEMA_signal_12087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7054 ( .C (clk), .D (new_AGEMA_signal_12090), .Q (new_AGEMA_signal_12091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7058 ( .C (clk), .D (new_AGEMA_signal_12094), .Q (new_AGEMA_signal_12095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7062 ( .C (clk), .D (new_AGEMA_signal_12098), .Q (new_AGEMA_signal_12099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7066 ( .C (clk), .D (new_AGEMA_signal_12102), .Q (new_AGEMA_signal_12103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7070 ( .C (clk), .D (new_AGEMA_signal_12106), .Q (new_AGEMA_signal_12107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7074 ( .C (clk), .D (new_AGEMA_signal_12110), .Q (new_AGEMA_signal_12111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7078 ( .C (clk), .D (new_AGEMA_signal_12114), .Q (new_AGEMA_signal_12115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7082 ( .C (clk), .D (new_AGEMA_signal_12118), .Q (new_AGEMA_signal_12119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7086 ( .C (clk), .D (new_AGEMA_signal_12122), .Q (new_AGEMA_signal_12123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7090 ( .C (clk), .D (new_AGEMA_signal_12126), .Q (new_AGEMA_signal_12127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7094 ( .C (clk), .D (new_AGEMA_signal_12130), .Q (new_AGEMA_signal_12131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7098 ( .C (clk), .D (new_AGEMA_signal_12134), .Q (new_AGEMA_signal_12135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7102 ( .C (clk), .D (new_AGEMA_signal_12138), .Q (new_AGEMA_signal_12139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7106 ( .C (clk), .D (new_AGEMA_signal_12142), .Q (new_AGEMA_signal_12143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7110 ( .C (clk), .D (new_AGEMA_signal_12146), .Q (new_AGEMA_signal_12147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7114 ( .C (clk), .D (new_AGEMA_signal_12150), .Q (new_AGEMA_signal_12151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7118 ( .C (clk), .D (new_AGEMA_signal_12154), .Q (new_AGEMA_signal_12155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7122 ( .C (clk), .D (new_AGEMA_signal_12158), .Q (new_AGEMA_signal_12159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7126 ( .C (clk), .D (new_AGEMA_signal_12162), .Q (new_AGEMA_signal_12163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7130 ( .C (clk), .D (new_AGEMA_signal_12166), .Q (new_AGEMA_signal_12167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7134 ( .C (clk), .D (new_AGEMA_signal_12170), .Q (new_AGEMA_signal_12171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7138 ( .C (clk), .D (new_AGEMA_signal_12174), .Q (new_AGEMA_signal_12175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7142 ( .C (clk), .D (new_AGEMA_signal_12178), .Q (new_AGEMA_signal_12179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7146 ( .C (clk), .D (new_AGEMA_signal_12182), .Q (new_AGEMA_signal_12183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7150 ( .C (clk), .D (new_AGEMA_signal_12186), .Q (new_AGEMA_signal_12187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7154 ( .C (clk), .D (new_AGEMA_signal_12190), .Q (new_AGEMA_signal_12191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7158 ( .C (clk), .D (new_AGEMA_signal_12194), .Q (new_AGEMA_signal_12195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7162 ( .C (clk), .D (new_AGEMA_signal_12198), .Q (new_AGEMA_signal_12199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7166 ( .C (clk), .D (new_AGEMA_signal_12202), .Q (new_AGEMA_signal_12203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7170 ( .C (clk), .D (new_AGEMA_signal_12206), .Q (new_AGEMA_signal_12207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7174 ( .C (clk), .D (new_AGEMA_signal_12210), .Q (new_AGEMA_signal_12211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7178 ( .C (clk), .D (new_AGEMA_signal_12214), .Q (new_AGEMA_signal_12215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7182 ( .C (clk), .D (new_AGEMA_signal_12218), .Q (new_AGEMA_signal_12219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7186 ( .C (clk), .D (new_AGEMA_signal_12222), .Q (new_AGEMA_signal_12223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7190 ( .C (clk), .D (new_AGEMA_signal_12226), .Q (new_AGEMA_signal_12227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7194 ( .C (clk), .D (new_AGEMA_signal_12230), .Q (new_AGEMA_signal_12231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7198 ( .C (clk), .D (new_AGEMA_signal_12234), .Q (new_AGEMA_signal_12235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7202 ( .C (clk), .D (new_AGEMA_signal_12238), .Q (new_AGEMA_signal_12239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7206 ( .C (clk), .D (new_AGEMA_signal_12242), .Q (new_AGEMA_signal_12243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7210 ( .C (clk), .D (new_AGEMA_signal_12246), .Q (new_AGEMA_signal_12247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7214 ( .C (clk), .D (new_AGEMA_signal_12250), .Q (new_AGEMA_signal_12251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7218 ( .C (clk), .D (new_AGEMA_signal_12254), .Q (new_AGEMA_signal_12255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7222 ( .C (clk), .D (new_AGEMA_signal_12258), .Q (new_AGEMA_signal_12259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7226 ( .C (clk), .D (new_AGEMA_signal_12262), .Q (new_AGEMA_signal_12263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7230 ( .C (clk), .D (new_AGEMA_signal_12266), .Q (new_AGEMA_signal_12267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7234 ( .C (clk), .D (new_AGEMA_signal_12270), .Q (new_AGEMA_signal_12271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7238 ( .C (clk), .D (new_AGEMA_signal_12274), .Q (new_AGEMA_signal_12275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7242 ( .C (clk), .D (new_AGEMA_signal_12278), .Q (new_AGEMA_signal_12279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7246 ( .C (clk), .D (new_AGEMA_signal_12282), .Q (new_AGEMA_signal_12283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7250 ( .C (clk), .D (new_AGEMA_signal_12286), .Q (new_AGEMA_signal_12287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7254 ( .C (clk), .D (new_AGEMA_signal_12290), .Q (new_AGEMA_signal_12291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7258 ( .C (clk), .D (new_AGEMA_signal_12294), .Q (new_AGEMA_signal_12295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7262 ( .C (clk), .D (new_AGEMA_signal_12298), .Q (new_AGEMA_signal_12299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7266 ( .C (clk), .D (new_AGEMA_signal_12302), .Q (new_AGEMA_signal_12303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7270 ( .C (clk), .D (new_AGEMA_signal_12306), .Q (new_AGEMA_signal_12307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7274 ( .C (clk), .D (new_AGEMA_signal_12310), .Q (new_AGEMA_signal_12311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7278 ( .C (clk), .D (new_AGEMA_signal_12314), .Q (new_AGEMA_signal_12315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7282 ( .C (clk), .D (new_AGEMA_signal_12318), .Q (new_AGEMA_signal_12319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7286 ( .C (clk), .D (new_AGEMA_signal_12322), .Q (new_AGEMA_signal_12323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7290 ( .C (clk), .D (new_AGEMA_signal_12326), .Q (new_AGEMA_signal_12327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7294 ( .C (clk), .D (new_AGEMA_signal_12330), .Q (new_AGEMA_signal_12331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7298 ( .C (clk), .D (new_AGEMA_signal_12334), .Q (new_AGEMA_signal_12335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7302 ( .C (clk), .D (new_AGEMA_signal_12338), .Q (new_AGEMA_signal_12339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7306 ( .C (clk), .D (new_AGEMA_signal_12342), .Q (new_AGEMA_signal_12343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7310 ( .C (clk), .D (new_AGEMA_signal_12346), .Q (new_AGEMA_signal_12347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7314 ( .C (clk), .D (new_AGEMA_signal_12350), .Q (new_AGEMA_signal_12351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7318 ( .C (clk), .D (new_AGEMA_signal_12354), .Q (new_AGEMA_signal_12355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7322 ( .C (clk), .D (new_AGEMA_signal_12358), .Q (new_AGEMA_signal_12359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7326 ( .C (clk), .D (new_AGEMA_signal_12362), .Q (new_AGEMA_signal_12363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7330 ( .C (clk), .D (new_AGEMA_signal_12366), .Q (new_AGEMA_signal_12367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7334 ( .C (clk), .D (new_AGEMA_signal_12370), .Q (new_AGEMA_signal_12371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7338 ( .C (clk), .D (new_AGEMA_signal_12374), .Q (new_AGEMA_signal_12375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7342 ( .C (clk), .D (new_AGEMA_signal_12378), .Q (new_AGEMA_signal_12379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7346 ( .C (clk), .D (new_AGEMA_signal_12382), .Q (new_AGEMA_signal_12383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7350 ( .C (clk), .D (new_AGEMA_signal_12386), .Q (new_AGEMA_signal_12387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7354 ( .C (clk), .D (new_AGEMA_signal_12390), .Q (new_AGEMA_signal_12391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7358 ( .C (clk), .D (new_AGEMA_signal_12394), .Q (new_AGEMA_signal_12395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7362 ( .C (clk), .D (new_AGEMA_signal_12398), .Q (new_AGEMA_signal_12399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7366 ( .C (clk), .D (new_AGEMA_signal_12402), .Q (new_AGEMA_signal_12403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7370 ( .C (clk), .D (new_AGEMA_signal_12406), .Q (new_AGEMA_signal_12407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7374 ( .C (clk), .D (new_AGEMA_signal_12410), .Q (new_AGEMA_signal_12411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7378 ( .C (clk), .D (new_AGEMA_signal_12414), .Q (new_AGEMA_signal_12415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7382 ( .C (clk), .D (new_AGEMA_signal_12418), .Q (new_AGEMA_signal_12419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7386 ( .C (clk), .D (new_AGEMA_signal_12422), .Q (new_AGEMA_signal_12423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7390 ( .C (clk), .D (new_AGEMA_signal_12426), .Q (new_AGEMA_signal_12427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7394 ( .C (clk), .D (new_AGEMA_signal_12430), .Q (new_AGEMA_signal_12431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7398 ( .C (clk), .D (new_AGEMA_signal_12434), .Q (new_AGEMA_signal_12435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7402 ( .C (clk), .D (new_AGEMA_signal_12438), .Q (new_AGEMA_signal_12439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7406 ( .C (clk), .D (new_AGEMA_signal_12442), .Q (new_AGEMA_signal_12443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7410 ( .C (clk), .D (new_AGEMA_signal_12446), .Q (new_AGEMA_signal_12447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7414 ( .C (clk), .D (new_AGEMA_signal_12450), .Q (new_AGEMA_signal_12451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7418 ( .C (clk), .D (new_AGEMA_signal_12454), .Q (new_AGEMA_signal_12455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7422 ( .C (clk), .D (new_AGEMA_signal_12458), .Q (new_AGEMA_signal_12459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7426 ( .C (clk), .D (new_AGEMA_signal_12462), .Q (new_AGEMA_signal_12463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7430 ( .C (clk), .D (new_AGEMA_signal_12466), .Q (new_AGEMA_signal_12467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7434 ( .C (clk), .D (new_AGEMA_signal_12470), .Q (new_AGEMA_signal_12471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7438 ( .C (clk), .D (new_AGEMA_signal_12474), .Q (new_AGEMA_signal_12475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7442 ( .C (clk), .D (new_AGEMA_signal_12478), .Q (new_AGEMA_signal_12479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7446 ( .C (clk), .D (new_AGEMA_signal_12482), .Q (new_AGEMA_signal_12483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7450 ( .C (clk), .D (new_AGEMA_signal_12486), .Q (new_AGEMA_signal_12487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7454 ( .C (clk), .D (new_AGEMA_signal_12490), .Q (new_AGEMA_signal_12491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7458 ( .C (clk), .D (new_AGEMA_signal_12494), .Q (new_AGEMA_signal_12495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7462 ( .C (clk), .D (new_AGEMA_signal_12498), .Q (new_AGEMA_signal_12499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7466 ( .C (clk), .D (new_AGEMA_signal_12502), .Q (new_AGEMA_signal_12503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7470 ( .C (clk), .D (new_AGEMA_signal_12506), .Q (new_AGEMA_signal_12507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7474 ( .C (clk), .D (new_AGEMA_signal_12510), .Q (new_AGEMA_signal_12511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7478 ( .C (clk), .D (new_AGEMA_signal_12514), .Q (new_AGEMA_signal_12515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7482 ( .C (clk), .D (new_AGEMA_signal_12518), .Q (new_AGEMA_signal_12519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7486 ( .C (clk), .D (new_AGEMA_signal_12522), .Q (new_AGEMA_signal_12523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7490 ( .C (clk), .D (new_AGEMA_signal_12526), .Q (new_AGEMA_signal_12527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7494 ( .C (clk), .D (new_AGEMA_signal_12530), .Q (new_AGEMA_signal_12531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7498 ( .C (clk), .D (new_AGEMA_signal_12534), .Q (new_AGEMA_signal_12535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7502 ( .C (clk), .D (new_AGEMA_signal_12538), .Q (new_AGEMA_signal_12539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7506 ( .C (clk), .D (new_AGEMA_signal_12542), .Q (new_AGEMA_signal_12543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7510 ( .C (clk), .D (new_AGEMA_signal_12546), .Q (new_AGEMA_signal_12547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7514 ( .C (clk), .D (new_AGEMA_signal_12550), .Q (new_AGEMA_signal_12551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7518 ( .C (clk), .D (new_AGEMA_signal_12554), .Q (new_AGEMA_signal_12555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7522 ( .C (clk), .D (new_AGEMA_signal_12558), .Q (new_AGEMA_signal_12559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7526 ( .C (clk), .D (new_AGEMA_signal_12562), .Q (new_AGEMA_signal_12563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7530 ( .C (clk), .D (new_AGEMA_signal_12566), .Q (new_AGEMA_signal_12567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7534 ( .C (clk), .D (new_AGEMA_signal_12570), .Q (new_AGEMA_signal_12571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7538 ( .C (clk), .D (new_AGEMA_signal_12574), .Q (new_AGEMA_signal_12575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7542 ( .C (clk), .D (new_AGEMA_signal_12578), .Q (new_AGEMA_signal_12579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7546 ( .C (clk), .D (new_AGEMA_signal_12582), .Q (new_AGEMA_signal_12583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7550 ( .C (clk), .D (new_AGEMA_signal_12586), .Q (new_AGEMA_signal_12587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7554 ( .C (clk), .D (new_AGEMA_signal_12590), .Q (new_AGEMA_signal_12591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7558 ( .C (clk), .D (new_AGEMA_signal_12594), .Q (new_AGEMA_signal_12595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7562 ( .C (clk), .D (new_AGEMA_signal_12598), .Q (new_AGEMA_signal_12599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7566 ( .C (clk), .D (new_AGEMA_signal_12602), .Q (new_AGEMA_signal_12603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7570 ( .C (clk), .D (new_AGEMA_signal_12606), .Q (new_AGEMA_signal_12607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7574 ( .C (clk), .D (new_AGEMA_signal_12610), .Q (new_AGEMA_signal_12611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7578 ( .C (clk), .D (new_AGEMA_signal_12614), .Q (new_AGEMA_signal_12615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7582 ( .C (clk), .D (new_AGEMA_signal_12618), .Q (new_AGEMA_signal_12619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7586 ( .C (clk), .D (new_AGEMA_signal_12622), .Q (new_AGEMA_signal_12623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7590 ( .C (clk), .D (new_AGEMA_signal_12626), .Q (new_AGEMA_signal_12627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7594 ( .C (clk), .D (new_AGEMA_signal_12630), .Q (new_AGEMA_signal_12631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7598 ( .C (clk), .D (new_AGEMA_signal_12634), .Q (new_AGEMA_signal_12635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7602 ( .C (clk), .D (new_AGEMA_signal_12638), .Q (new_AGEMA_signal_12639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7606 ( .C (clk), .D (new_AGEMA_signal_12642), .Q (new_AGEMA_signal_12643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7610 ( .C (clk), .D (new_AGEMA_signal_12646), .Q (new_AGEMA_signal_12647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7614 ( .C (clk), .D (new_AGEMA_signal_12650), .Q (new_AGEMA_signal_12651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7618 ( .C (clk), .D (new_AGEMA_signal_12654), .Q (new_AGEMA_signal_12655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7622 ( .C (clk), .D (new_AGEMA_signal_12658), .Q (new_AGEMA_signal_12659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7626 ( .C (clk), .D (new_AGEMA_signal_12662), .Q (new_AGEMA_signal_12663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7630 ( .C (clk), .D (new_AGEMA_signal_12666), .Q (new_AGEMA_signal_12667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7634 ( .C (clk), .D (new_AGEMA_signal_12670), .Q (new_AGEMA_signal_12671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7638 ( .C (clk), .D (new_AGEMA_signal_12674), .Q (new_AGEMA_signal_12675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7642 ( .C (clk), .D (new_AGEMA_signal_12678), .Q (new_AGEMA_signal_12679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7646 ( .C (clk), .D (new_AGEMA_signal_12682), .Q (new_AGEMA_signal_12683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7650 ( .C (clk), .D (new_AGEMA_signal_12686), .Q (new_AGEMA_signal_12687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7654 ( .C (clk), .D (new_AGEMA_signal_12690), .Q (new_AGEMA_signal_12691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7658 ( .C (clk), .D (new_AGEMA_signal_12694), .Q (new_AGEMA_signal_12695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7662 ( .C (clk), .D (new_AGEMA_signal_12698), .Q (new_AGEMA_signal_12699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7666 ( .C (clk), .D (new_AGEMA_signal_12702), .Q (new_AGEMA_signal_12703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7670 ( .C (clk), .D (new_AGEMA_signal_12706), .Q (new_AGEMA_signal_12707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7674 ( .C (clk), .D (new_AGEMA_signal_12710), .Q (new_AGEMA_signal_12711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7678 ( .C (clk), .D (new_AGEMA_signal_12714), .Q (new_AGEMA_signal_12715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7682 ( .C (clk), .D (new_AGEMA_signal_12718), .Q (new_AGEMA_signal_12719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7686 ( .C (clk), .D (new_AGEMA_signal_12722), .Q (new_AGEMA_signal_12723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7690 ( .C (clk), .D (new_AGEMA_signal_12726), .Q (new_AGEMA_signal_12727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7694 ( .C (clk), .D (new_AGEMA_signal_12730), .Q (new_AGEMA_signal_12731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7698 ( .C (clk), .D (new_AGEMA_signal_12734), .Q (new_AGEMA_signal_12735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7702 ( .C (clk), .D (new_AGEMA_signal_12738), .Q (new_AGEMA_signal_12739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7706 ( .C (clk), .D (new_AGEMA_signal_12742), .Q (new_AGEMA_signal_12743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7710 ( .C (clk), .D (new_AGEMA_signal_12746), .Q (new_AGEMA_signal_12747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7714 ( .C (clk), .D (new_AGEMA_signal_12750), .Q (new_AGEMA_signal_12751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7718 ( .C (clk), .D (new_AGEMA_signal_12754), .Q (new_AGEMA_signal_12755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7722 ( .C (clk), .D (new_AGEMA_signal_12758), .Q (new_AGEMA_signal_12759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7726 ( .C (clk), .D (new_AGEMA_signal_12762), .Q (new_AGEMA_signal_12763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7730 ( .C (clk), .D (new_AGEMA_signal_12766), .Q (new_AGEMA_signal_12767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7734 ( .C (clk), .D (new_AGEMA_signal_12770), .Q (new_AGEMA_signal_12771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7738 ( .C (clk), .D (new_AGEMA_signal_12774), .Q (new_AGEMA_signal_12775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7742 ( .C (clk), .D (new_AGEMA_signal_12778), .Q (new_AGEMA_signal_12779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7746 ( .C (clk), .D (new_AGEMA_signal_12782), .Q (new_AGEMA_signal_12783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7750 ( .C (clk), .D (new_AGEMA_signal_12786), .Q (new_AGEMA_signal_12787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7754 ( .C (clk), .D (new_AGEMA_signal_12790), .Q (new_AGEMA_signal_12791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7758 ( .C (clk), .D (new_AGEMA_signal_12794), .Q (new_AGEMA_signal_12795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7762 ( .C (clk), .D (new_AGEMA_signal_12798), .Q (new_AGEMA_signal_12799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7766 ( .C (clk), .D (new_AGEMA_signal_12802), .Q (new_AGEMA_signal_12803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7770 ( .C (clk), .D (new_AGEMA_signal_12806), .Q (new_AGEMA_signal_12807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7774 ( .C (clk), .D (new_AGEMA_signal_12810), .Q (new_AGEMA_signal_12811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7778 ( .C (clk), .D (new_AGEMA_signal_12814), .Q (new_AGEMA_signal_12815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7782 ( .C (clk), .D (new_AGEMA_signal_12818), .Q (new_AGEMA_signal_12819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7786 ( .C (clk), .D (new_AGEMA_signal_12822), .Q (new_AGEMA_signal_12823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7790 ( .C (clk), .D (new_AGEMA_signal_12826), .Q (new_AGEMA_signal_12827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7794 ( .C (clk), .D (new_AGEMA_signal_12830), .Q (new_AGEMA_signal_12831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7798 ( .C (clk), .D (new_AGEMA_signal_12834), .Q (new_AGEMA_signal_12835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7802 ( .C (clk), .D (new_AGEMA_signal_12838), .Q (new_AGEMA_signal_12839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7806 ( .C (clk), .D (new_AGEMA_signal_12842), .Q (new_AGEMA_signal_12843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7810 ( .C (clk), .D (new_AGEMA_signal_12846), .Q (new_AGEMA_signal_12847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7814 ( .C (clk), .D (new_AGEMA_signal_12850), .Q (new_AGEMA_signal_12851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7818 ( .C (clk), .D (new_AGEMA_signal_12854), .Q (new_AGEMA_signal_12855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7822 ( .C (clk), .D (new_AGEMA_signal_12858), .Q (new_AGEMA_signal_12859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7826 ( .C (clk), .D (new_AGEMA_signal_12862), .Q (new_AGEMA_signal_12863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7830 ( .C (clk), .D (new_AGEMA_signal_12866), .Q (new_AGEMA_signal_12867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7834 ( .C (clk), .D (new_AGEMA_signal_12870), .Q (new_AGEMA_signal_12871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7838 ( .C (clk), .D (new_AGEMA_signal_12874), .Q (new_AGEMA_signal_12875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7842 ( .C (clk), .D (new_AGEMA_signal_12878), .Q (new_AGEMA_signal_12879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7846 ( .C (clk), .D (new_AGEMA_signal_12882), .Q (new_AGEMA_signal_12883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7850 ( .C (clk), .D (new_AGEMA_signal_12886), .Q (new_AGEMA_signal_12887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7854 ( .C (clk), .D (new_AGEMA_signal_12890), .Q (new_AGEMA_signal_12891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7858 ( .C (clk), .D (new_AGEMA_signal_12894), .Q (new_AGEMA_signal_12895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7862 ( .C (clk), .D (new_AGEMA_signal_12898), .Q (new_AGEMA_signal_12899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7866 ( .C (clk), .D (new_AGEMA_signal_12902), .Q (new_AGEMA_signal_12903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7870 ( .C (clk), .D (new_AGEMA_signal_12906), .Q (new_AGEMA_signal_12907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7874 ( .C (clk), .D (new_AGEMA_signal_12910), .Q (new_AGEMA_signal_12911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7878 ( .C (clk), .D (new_AGEMA_signal_12914), .Q (new_AGEMA_signal_12915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7882 ( .C (clk), .D (new_AGEMA_signal_12918), .Q (new_AGEMA_signal_12919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7886 ( .C (clk), .D (new_AGEMA_signal_12922), .Q (new_AGEMA_signal_12923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7890 ( .C (clk), .D (new_AGEMA_signal_12926), .Q (new_AGEMA_signal_12927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7894 ( .C (clk), .D (new_AGEMA_signal_12930), .Q (new_AGEMA_signal_12931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7898 ( .C (clk), .D (new_AGEMA_signal_12934), .Q (new_AGEMA_signal_12935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7902 ( .C (clk), .D (new_AGEMA_signal_12938), .Q (new_AGEMA_signal_12939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7906 ( .C (clk), .D (new_AGEMA_signal_12942), .Q (new_AGEMA_signal_12943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7910 ( .C (clk), .D (new_AGEMA_signal_12946), .Q (new_AGEMA_signal_12947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7914 ( .C (clk), .D (new_AGEMA_signal_12950), .Q (new_AGEMA_signal_12951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7918 ( .C (clk), .D (new_AGEMA_signal_12954), .Q (new_AGEMA_signal_12955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7922 ( .C (clk), .D (new_AGEMA_signal_12958), .Q (new_AGEMA_signal_12959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7926 ( .C (clk), .D (new_AGEMA_signal_12962), .Q (new_AGEMA_signal_12963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7930 ( .C (clk), .D (new_AGEMA_signal_12966), .Q (new_AGEMA_signal_12967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7934 ( .C (clk), .D (new_AGEMA_signal_12970), .Q (new_AGEMA_signal_12971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7938 ( .C (clk), .D (new_AGEMA_signal_12974), .Q (new_AGEMA_signal_12975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7942 ( .C (clk), .D (new_AGEMA_signal_12978), .Q (new_AGEMA_signal_12979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7946 ( .C (clk), .D (new_AGEMA_signal_12982), .Q (new_AGEMA_signal_12983) ) ;
    buf_clk new_AGEMA_reg_buffer_7950 ( .C (clk), .D (new_AGEMA_signal_12986), .Q (new_AGEMA_signal_12987) ) ;
    buf_clk new_AGEMA_reg_buffer_7954 ( .C (clk), .D (new_AGEMA_signal_12990), .Q (new_AGEMA_signal_12991) ) ;
    buf_clk new_AGEMA_reg_buffer_7958 ( .C (clk), .D (new_AGEMA_signal_12994), .Q (new_AGEMA_signal_12995) ) ;
    buf_clk new_AGEMA_reg_buffer_7962 ( .C (clk), .D (new_AGEMA_signal_12998), .Q (new_AGEMA_signal_12999) ) ;
    buf_clk new_AGEMA_reg_buffer_7966 ( .C (clk), .D (new_AGEMA_signal_13002), .Q (new_AGEMA_signal_13003) ) ;
    buf_clk new_AGEMA_reg_buffer_7970 ( .C (clk), .D (new_AGEMA_signal_13006), .Q (new_AGEMA_signal_13007) ) ;
    buf_clk new_AGEMA_reg_buffer_7974 ( .C (clk), .D (new_AGEMA_signal_13010), .Q (new_AGEMA_signal_13011) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_4175, new_AGEMA_signal_4174, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, new_AGEMA_signal_7152}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_4211, new_AGEMA_signal_4210, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_7157, new_AGEMA_signal_7156, new_AGEMA_signal_7155}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_7154, new_AGEMA_signal_7153, new_AGEMA_signal_7152}), .b ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_7157, new_AGEMA_signal_7156, new_AGEMA_signal_7155}), .b ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_7196, new_AGEMA_signal_7195, new_AGEMA_signal_7194}), .b ({new_AGEMA_signal_4211, new_AGEMA_signal_4210, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_7199, new_AGEMA_signal_7198, new_AGEMA_signal_7197}), .c ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_7202, new_AGEMA_signal_7201, new_AGEMA_signal_7200}), .b ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_7205, new_AGEMA_signal_7204, new_AGEMA_signal_7203}), .c ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, new_AGEMA_signal_7164}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_4183, new_AGEMA_signal_4182, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_7169, new_AGEMA_signal_7168, new_AGEMA_signal_7167}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_7166, new_AGEMA_signal_7165, new_AGEMA_signal_7164}), .b ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_7169, new_AGEMA_signal_7168, new_AGEMA_signal_7167}), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_7208, new_AGEMA_signal_7207, new_AGEMA_signal_7206}), .b ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_7211, new_AGEMA_signal_7210, new_AGEMA_signal_7209}), .c ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_7214, new_AGEMA_signal_7213, new_AGEMA_signal_7212}), .b ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_7217, new_AGEMA_signal_7216, new_AGEMA_signal_7215}), .c ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, new_AGEMA_signal_7176}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_4193, new_AGEMA_signal_4192, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_7181, new_AGEMA_signal_7180, new_AGEMA_signal_7179}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_7178, new_AGEMA_signal_7177, new_AGEMA_signal_7176}), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_7181, new_AGEMA_signal_7180, new_AGEMA_signal_7179}), .b ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_7220, new_AGEMA_signal_7219, new_AGEMA_signal_7218}), .b ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_7223, new_AGEMA_signal_7222, new_AGEMA_signal_7221}), .c ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_7226, new_AGEMA_signal_7225, new_AGEMA_signal_7224}), .b ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_7229, new_AGEMA_signal_7228, new_AGEMA_signal_7227}), .c ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, new_AGEMA_signal_7188}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_7193, new_AGEMA_signal_7192, new_AGEMA_signal_7191}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_7190, new_AGEMA_signal_7189, new_AGEMA_signal_7188}), .b ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_7193, new_AGEMA_signal_7192, new_AGEMA_signal_7191}), .b ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_4247, new_AGEMA_signal_4246, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_7232, new_AGEMA_signal_7231, new_AGEMA_signal_7230}), .b ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_7235, new_AGEMA_signal_7234, new_AGEMA_signal_7233}), .c ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_7238, new_AGEMA_signal_7237, new_AGEMA_signal_7236}), .b ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_4247, new_AGEMA_signal_4246, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_7241, new_AGEMA_signal_7240, new_AGEMA_signal_7239}), .c ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_7146), .Q (new_AGEMA_signal_7194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_7195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_7148), .Q (new_AGEMA_signal_7196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2160 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_7197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_7198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_4179), .Q (new_AGEMA_signal_7199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_7149), .Q (new_AGEMA_signal_7200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_7150), .Q (new_AGEMA_signal_7201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_7202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2166 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_7203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_4218), .Q (new_AGEMA_signal_7204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_4219), .Q (new_AGEMA_signal_7205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_7158), .Q (new_AGEMA_signal_7206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_7159), .Q (new_AGEMA_signal_7207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_7160), .Q (new_AGEMA_signal_7208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2172 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_7209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_4188), .Q (new_AGEMA_signal_7210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_4189), .Q (new_AGEMA_signal_7211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_7161), .Q (new_AGEMA_signal_7212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_7162), .Q (new_AGEMA_signal_7213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_7163), .Q (new_AGEMA_signal_7214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2178 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_7215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_7216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_7217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_7170), .Q (new_AGEMA_signal_7218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_7171), .Q (new_AGEMA_signal_7219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_7220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2184 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_7221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_7222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_4199), .Q (new_AGEMA_signal_7223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_7173), .Q (new_AGEMA_signal_7224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_7174), .Q (new_AGEMA_signal_7225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_7175), .Q (new_AGEMA_signal_7226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2190 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_7227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_7228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_4239), .Q (new_AGEMA_signal_7229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_7182), .Q (new_AGEMA_signal_7230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_7231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_7184), .Q (new_AGEMA_signal_7232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2196 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_7233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_7234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_7235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_7185), .Q (new_AGEMA_signal_7236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_7237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_7238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2202 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_7239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_4248), .Q (new_AGEMA_signal_7240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_7241) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_7243), .Q (new_AGEMA_signal_7244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_7247), .Q (new_AGEMA_signal_7248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_7251), .Q (new_AGEMA_signal_7252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_7256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_7260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_7263), .Q (new_AGEMA_signal_7264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_7267), .Q (new_AGEMA_signal_7268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_7271), .Q (new_AGEMA_signal_7272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_7275), .Q (new_AGEMA_signal_7276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_7279), .Q (new_AGEMA_signal_7280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_7283), .Q (new_AGEMA_signal_7284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_7287), .Q (new_AGEMA_signal_7288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_7292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_7296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_7299), .Q (new_AGEMA_signal_7300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_7303), .Q (new_AGEMA_signal_7304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_7307), .Q (new_AGEMA_signal_7308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_7311), .Q (new_AGEMA_signal_7312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_7315), .Q (new_AGEMA_signal_7316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_7319), .Q (new_AGEMA_signal_7320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_7323), .Q (new_AGEMA_signal_7324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_7328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_7332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_7336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_7339), .Q (new_AGEMA_signal_7340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_7344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_7347), .Q (new_AGEMA_signal_7348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_7351), .Q (new_AGEMA_signal_7352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_7355), .Q (new_AGEMA_signal_7356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_7359), .Q (new_AGEMA_signal_7360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_7363), .Q (new_AGEMA_signal_7364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_7368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_7371), .Q (new_AGEMA_signal_7372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_7376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_7379), .Q (new_AGEMA_signal_7380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_7384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_7387), .Q (new_AGEMA_signal_7388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_7391), .Q (new_AGEMA_signal_7392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_7395), .Q (new_AGEMA_signal_7396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_7399), .Q (new_AGEMA_signal_7400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_7403), .Q (new_AGEMA_signal_7404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_7408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_7411), .Q (new_AGEMA_signal_7412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_7416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_7419), .Q (new_AGEMA_signal_7420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_7424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_7427), .Q (new_AGEMA_signal_7428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_7431), .Q (new_AGEMA_signal_7432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_7435), .Q (new_AGEMA_signal_7436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_7439), .Q (new_AGEMA_signal_7440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_7443), .Q (new_AGEMA_signal_7444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_7448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_7451), .Q (new_AGEMA_signal_7452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_7456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_7459), .Q (new_AGEMA_signal_7460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_7464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_7467), .Q (new_AGEMA_signal_7468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_7471), .Q (new_AGEMA_signal_7472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_7475), .Q (new_AGEMA_signal_7476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_7479), .Q (new_AGEMA_signal_7480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_7483), .Q (new_AGEMA_signal_7484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_7488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_7491), .Q (new_AGEMA_signal_7492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_7496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_7499), .Q (new_AGEMA_signal_7500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_7504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_7507), .Q (new_AGEMA_signal_7508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_7511), .Q (new_AGEMA_signal_7512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_7515), .Q (new_AGEMA_signal_7516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_7519), .Q (new_AGEMA_signal_7520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_7523), .Q (new_AGEMA_signal_7524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_7528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_7531), .Q (new_AGEMA_signal_7532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_7536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_7539), .Q (new_AGEMA_signal_7540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_7543), .Q (new_AGEMA_signal_7544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_7547), .Q (new_AGEMA_signal_7548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_7551), .Q (new_AGEMA_signal_7552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_7555), .Q (new_AGEMA_signal_7556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_7559), .Q (new_AGEMA_signal_7560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_7563), .Q (new_AGEMA_signal_7564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_7567), .Q (new_AGEMA_signal_7568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_7571), .Q (new_AGEMA_signal_7572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_7575), .Q (new_AGEMA_signal_7576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_7579), .Q (new_AGEMA_signal_7580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_7583), .Q (new_AGEMA_signal_7584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_7587), .Q (new_AGEMA_signal_7588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_7591), .Q (new_AGEMA_signal_7592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_7595), .Q (new_AGEMA_signal_7596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_7599), .Q (new_AGEMA_signal_7600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_7603), .Q (new_AGEMA_signal_7604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_7607), .Q (new_AGEMA_signal_7608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_7611), .Q (new_AGEMA_signal_7612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_7616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_7619), .Q (new_AGEMA_signal_7620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_7623), .Q (new_AGEMA_signal_7624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_7627), .Q (new_AGEMA_signal_7628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_7631), .Q (new_AGEMA_signal_7632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_7634), .Q (new_AGEMA_signal_7635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_7637), .Q (new_AGEMA_signal_7638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_7640), .Q (new_AGEMA_signal_7641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_7643), .Q (new_AGEMA_signal_7644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_7646), .Q (new_AGEMA_signal_7647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2613 ( .C (clk), .D (new_AGEMA_signal_7649), .Q (new_AGEMA_signal_7650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_7652), .Q (new_AGEMA_signal_7653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_7655), .Q (new_AGEMA_signal_7656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_7658), .Q (new_AGEMA_signal_7659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_7661), .Q (new_AGEMA_signal_7662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_7664), .Q (new_AGEMA_signal_7665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_7667), .Q (new_AGEMA_signal_7668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_7670), .Q (new_AGEMA_signal_7671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_7673), .Q (new_AGEMA_signal_7674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_7676), .Q (new_AGEMA_signal_7677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_7679), .Q (new_AGEMA_signal_7680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_7682), .Q (new_AGEMA_signal_7683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_7685), .Q (new_AGEMA_signal_7686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_7688), .Q (new_AGEMA_signal_7689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_7691), .Q (new_AGEMA_signal_7692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_7694), .Q (new_AGEMA_signal_7695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_7697), .Q (new_AGEMA_signal_7698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_7700), .Q (new_AGEMA_signal_7701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_7703), .Q (new_AGEMA_signal_7704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_7706), .Q (new_AGEMA_signal_7707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_7709), .Q (new_AGEMA_signal_7710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_7712), .Q (new_AGEMA_signal_7713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_7715), .Q (new_AGEMA_signal_7716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_7718), .Q (new_AGEMA_signal_7719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_7721), .Q (new_AGEMA_signal_7722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_7724), .Q (new_AGEMA_signal_7725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_7727), .Q (new_AGEMA_signal_7728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_7730), .Q (new_AGEMA_signal_7731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_7733), .Q (new_AGEMA_signal_7734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_7736), .Q (new_AGEMA_signal_7737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_7739), .Q (new_AGEMA_signal_7740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_7742), .Q (new_AGEMA_signal_7743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_7745), .Q (new_AGEMA_signal_7746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_7748), .Q (new_AGEMA_signal_7749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_7751), .Q (new_AGEMA_signal_7752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_7754), .Q (new_AGEMA_signal_7755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_7757), .Q (new_AGEMA_signal_7758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_7760), .Q (new_AGEMA_signal_7761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_7763), .Q (new_AGEMA_signal_7764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_7766), .Q (new_AGEMA_signal_7767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_7769), .Q (new_AGEMA_signal_7770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_7772), .Q (new_AGEMA_signal_7773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_7775), .Q (new_AGEMA_signal_7776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_7778), .Q (new_AGEMA_signal_7779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_7781), .Q (new_AGEMA_signal_7782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_7784), .Q (new_AGEMA_signal_7785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_7787), .Q (new_AGEMA_signal_7788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_7790), .Q (new_AGEMA_signal_7791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_7793), .Q (new_AGEMA_signal_7794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_7796), .Q (new_AGEMA_signal_7797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_7799), .Q (new_AGEMA_signal_7800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_7802), .Q (new_AGEMA_signal_7803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_7805), .Q (new_AGEMA_signal_7806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_7808), .Q (new_AGEMA_signal_7809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_7811), .Q (new_AGEMA_signal_7812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_7814), .Q (new_AGEMA_signal_7815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_7817), .Q (new_AGEMA_signal_7818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_7820), .Q (new_AGEMA_signal_7821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_7823), .Q (new_AGEMA_signal_7824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_7826), .Q (new_AGEMA_signal_7827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_7829), .Q (new_AGEMA_signal_7830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_7832), .Q (new_AGEMA_signal_7833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_7835), .Q (new_AGEMA_signal_7836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_7838), .Q (new_AGEMA_signal_7839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_7841), .Q (new_AGEMA_signal_7842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_7844), .Q (new_AGEMA_signal_7845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_7847), .Q (new_AGEMA_signal_7848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_7850), .Q (new_AGEMA_signal_7851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_7853), .Q (new_AGEMA_signal_7854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_7856), .Q (new_AGEMA_signal_7857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_7859), .Q (new_AGEMA_signal_7860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_7862), .Q (new_AGEMA_signal_7863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_7865), .Q (new_AGEMA_signal_7866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_7868), .Q (new_AGEMA_signal_7869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_7871), .Q (new_AGEMA_signal_7872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_7874), .Q (new_AGEMA_signal_7875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_7877), .Q (new_AGEMA_signal_7878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_7880), .Q (new_AGEMA_signal_7881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_7883), .Q (new_AGEMA_signal_7884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_7886), .Q (new_AGEMA_signal_7887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_7889), .Q (new_AGEMA_signal_7890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_7892), .Q (new_AGEMA_signal_7893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_7895), .Q (new_AGEMA_signal_7896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_7898), .Q (new_AGEMA_signal_7899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2865 ( .C (clk), .D (new_AGEMA_signal_7901), .Q (new_AGEMA_signal_7902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_7904), .Q (new_AGEMA_signal_7905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_7907), .Q (new_AGEMA_signal_7908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_7910), .Q (new_AGEMA_signal_7911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_7913), .Q (new_AGEMA_signal_7914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_7916), .Q (new_AGEMA_signal_7917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_7919), .Q (new_AGEMA_signal_7920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_7922), .Q (new_AGEMA_signal_7923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_7925), .Q (new_AGEMA_signal_7926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_7928), .Q (new_AGEMA_signal_7929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_7931), .Q (new_AGEMA_signal_7932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_7934), .Q (new_AGEMA_signal_7935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2901 ( .C (clk), .D (new_AGEMA_signal_7937), .Q (new_AGEMA_signal_7938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_7940), .Q (new_AGEMA_signal_7941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_7943), .Q (new_AGEMA_signal_7944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_7946), .Q (new_AGEMA_signal_7947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_7949), .Q (new_AGEMA_signal_7950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_7952), .Q (new_AGEMA_signal_7953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_7955), .Q (new_AGEMA_signal_7956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_7958), .Q (new_AGEMA_signal_7959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_7961), .Q (new_AGEMA_signal_7962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_7964), .Q (new_AGEMA_signal_7965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_7967), .Q (new_AGEMA_signal_7968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_7970), .Q (new_AGEMA_signal_7971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2937 ( .C (clk), .D (new_AGEMA_signal_7973), .Q (new_AGEMA_signal_7974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_7976), .Q (new_AGEMA_signal_7977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_7979), .Q (new_AGEMA_signal_7980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_7982), .Q (new_AGEMA_signal_7983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_7985), .Q (new_AGEMA_signal_7986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_7988), .Q (new_AGEMA_signal_7989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_7991), .Q (new_AGEMA_signal_7992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_7994), .Q (new_AGEMA_signal_7995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_7997), .Q (new_AGEMA_signal_7998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_8000), .Q (new_AGEMA_signal_8001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_8003), .Q (new_AGEMA_signal_8004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_8006), .Q (new_AGEMA_signal_8007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_8009), .Q (new_AGEMA_signal_8010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_8012), .Q (new_AGEMA_signal_8013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_8015), .Q (new_AGEMA_signal_8016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_8018), .Q (new_AGEMA_signal_8019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_8021), .Q (new_AGEMA_signal_8022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_8024), .Q (new_AGEMA_signal_8025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_8027), .Q (new_AGEMA_signal_8028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_8030), .Q (new_AGEMA_signal_8031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_8033), .Q (new_AGEMA_signal_8034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_8036), .Q (new_AGEMA_signal_8037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_8039), .Q (new_AGEMA_signal_8040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_8042), .Q (new_AGEMA_signal_8043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_8045), .Q (new_AGEMA_signal_8046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_8048), .Q (new_AGEMA_signal_8049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_8051), .Q (new_AGEMA_signal_8052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_8054), .Q (new_AGEMA_signal_8055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_8057), .Q (new_AGEMA_signal_8058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_8060), .Q (new_AGEMA_signal_8061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_8063), .Q (new_AGEMA_signal_8064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_8066), .Q (new_AGEMA_signal_8067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_8069), .Q (new_AGEMA_signal_8070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_8072), .Q (new_AGEMA_signal_8073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_8075), .Q (new_AGEMA_signal_8076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_8078), .Q (new_AGEMA_signal_8079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_8081), .Q (new_AGEMA_signal_8082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_8084), .Q (new_AGEMA_signal_8085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3051 ( .C (clk), .D (new_AGEMA_signal_8087), .Q (new_AGEMA_signal_8088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_8090), .Q (new_AGEMA_signal_8091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_8093), .Q (new_AGEMA_signal_8094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_8096), .Q (new_AGEMA_signal_8097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_8099), .Q (new_AGEMA_signal_8100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_8102), .Q (new_AGEMA_signal_8103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_8105), .Q (new_AGEMA_signal_8106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_8108), .Q (new_AGEMA_signal_8109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_8111), .Q (new_AGEMA_signal_8112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_8114), .Q (new_AGEMA_signal_8115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_8117), .Q (new_AGEMA_signal_8118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_8120), .Q (new_AGEMA_signal_8121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_8123), .Q (new_AGEMA_signal_8124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_8126), .Q (new_AGEMA_signal_8127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_8129), .Q (new_AGEMA_signal_8130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_8132), .Q (new_AGEMA_signal_8133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_8135), .Q (new_AGEMA_signal_8136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_8138), .Q (new_AGEMA_signal_8139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_8141), .Q (new_AGEMA_signal_8142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_8144), .Q (new_AGEMA_signal_8145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_8147), .Q (new_AGEMA_signal_8148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_8150), .Q (new_AGEMA_signal_8151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_8153), .Q (new_AGEMA_signal_8154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_8156), .Q (new_AGEMA_signal_8157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_8159), .Q (new_AGEMA_signal_8160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_8162), .Q (new_AGEMA_signal_8163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_8165), .Q (new_AGEMA_signal_8166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_8168), .Q (new_AGEMA_signal_8169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_8171), .Q (new_AGEMA_signal_8172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_8174), .Q (new_AGEMA_signal_8175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_8177), .Q (new_AGEMA_signal_8178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_8180), .Q (new_AGEMA_signal_8181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_8183), .Q (new_AGEMA_signal_8184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_8186), .Q (new_AGEMA_signal_8187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_8189), .Q (new_AGEMA_signal_8190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_8192), .Q (new_AGEMA_signal_8193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_8195), .Q (new_AGEMA_signal_8196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_8198), .Q (new_AGEMA_signal_8199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_8201), .Q (new_AGEMA_signal_8202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_8204), .Q (new_AGEMA_signal_8205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_8207), .Q (new_AGEMA_signal_8208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_8210), .Q (new_AGEMA_signal_8211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_8213), .Q (new_AGEMA_signal_8214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_8216), .Q (new_AGEMA_signal_8217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_8219), .Q (new_AGEMA_signal_8220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_8222), .Q (new_AGEMA_signal_8223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_8225), .Q (new_AGEMA_signal_8226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_8228), .Q (new_AGEMA_signal_8229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_8231), .Q (new_AGEMA_signal_8232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_8234), .Q (new_AGEMA_signal_8235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_8237), .Q (new_AGEMA_signal_8238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_8240), .Q (new_AGEMA_signal_8241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_8243), .Q (new_AGEMA_signal_8244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_8246), .Q (new_AGEMA_signal_8247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_8249), .Q (new_AGEMA_signal_8250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_8252), .Q (new_AGEMA_signal_8253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_8255), .Q (new_AGEMA_signal_8256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_8258), .Q (new_AGEMA_signal_8259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_8261), .Q (new_AGEMA_signal_8262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_8264), .Q (new_AGEMA_signal_8265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_8267), .Q (new_AGEMA_signal_8268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_8270), .Q (new_AGEMA_signal_8271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_8273), .Q (new_AGEMA_signal_8274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_8276), .Q (new_AGEMA_signal_8277) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_8279), .Q (new_AGEMA_signal_8280) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_8283), .Q (new_AGEMA_signal_8284) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_8287), .Q (new_AGEMA_signal_8288) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_8291), .Q (new_AGEMA_signal_8292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_8295), .Q (new_AGEMA_signal_8296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_8299), .Q (new_AGEMA_signal_8300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_8303), .Q (new_AGEMA_signal_8304) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_8307), .Q (new_AGEMA_signal_8308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_8311), .Q (new_AGEMA_signal_8312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_8315), .Q (new_AGEMA_signal_8316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_8319), .Q (new_AGEMA_signal_8320) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_8323), .Q (new_AGEMA_signal_8324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_8327), .Q (new_AGEMA_signal_8328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_8331), .Q (new_AGEMA_signal_8332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_8335), .Q (new_AGEMA_signal_8336) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_8339), .Q (new_AGEMA_signal_8340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_8343), .Q (new_AGEMA_signal_8344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_8347), .Q (new_AGEMA_signal_8348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_8351), .Q (new_AGEMA_signal_8352) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_8355), .Q (new_AGEMA_signal_8356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_8359), .Q (new_AGEMA_signal_8360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_8363), .Q (new_AGEMA_signal_8364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_8367), .Q (new_AGEMA_signal_8368) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_8371), .Q (new_AGEMA_signal_8372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3339 ( .C (clk), .D (new_AGEMA_signal_8375), .Q (new_AGEMA_signal_8376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_8379), .Q (new_AGEMA_signal_8380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_8383), .Q (new_AGEMA_signal_8384) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_8387), .Q (new_AGEMA_signal_8388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_8391), .Q (new_AGEMA_signal_8392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_8395), .Q (new_AGEMA_signal_8396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_8399), .Q (new_AGEMA_signal_8400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_8403), .Q (new_AGEMA_signal_8404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_8407), .Q (new_AGEMA_signal_8408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_8411), .Q (new_AGEMA_signal_8412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_8415), .Q (new_AGEMA_signal_8416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_8419), .Q (new_AGEMA_signal_8420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_8423), .Q (new_AGEMA_signal_8424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_8427), .Q (new_AGEMA_signal_8428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_8431), .Q (new_AGEMA_signal_8432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_8435), .Q (new_AGEMA_signal_8436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_8439), .Q (new_AGEMA_signal_8440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_8443), .Q (new_AGEMA_signal_8444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_8447), .Q (new_AGEMA_signal_8448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_8451), .Q (new_AGEMA_signal_8452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_8455), .Q (new_AGEMA_signal_8456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_8459), .Q (new_AGEMA_signal_8460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_8463), .Q (new_AGEMA_signal_8464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_8467), .Q (new_AGEMA_signal_8468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_8471), .Q (new_AGEMA_signal_8472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_8475), .Q (new_AGEMA_signal_8476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_8479), .Q (new_AGEMA_signal_8480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_8483), .Q (new_AGEMA_signal_8484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_8487), .Q (new_AGEMA_signal_8488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_8491), .Q (new_AGEMA_signal_8492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_8495), .Q (new_AGEMA_signal_8496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_8499), .Q (new_AGEMA_signal_8500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_8503), .Q (new_AGEMA_signal_8504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_8507), .Q (new_AGEMA_signal_8508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_8511), .Q (new_AGEMA_signal_8512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_8515), .Q (new_AGEMA_signal_8516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_8519), .Q (new_AGEMA_signal_8520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_8523), .Q (new_AGEMA_signal_8524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_8527), .Q (new_AGEMA_signal_8528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_8531), .Q (new_AGEMA_signal_8532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_8535), .Q (new_AGEMA_signal_8536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_8539), .Q (new_AGEMA_signal_8540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_8543), .Q (new_AGEMA_signal_8544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_8547), .Q (new_AGEMA_signal_8548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_8551), .Q (new_AGEMA_signal_8552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_8555), .Q (new_AGEMA_signal_8556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_8559), .Q (new_AGEMA_signal_8560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_8563), .Q (new_AGEMA_signal_8564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_8567), .Q (new_AGEMA_signal_8568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_8571), .Q (new_AGEMA_signal_8572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_8575), .Q (new_AGEMA_signal_8576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_8579), .Q (new_AGEMA_signal_8580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_8583), .Q (new_AGEMA_signal_8584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_8587), .Q (new_AGEMA_signal_8588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_8591), .Q (new_AGEMA_signal_8592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_8595), .Q (new_AGEMA_signal_8596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_8599), .Q (new_AGEMA_signal_8600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_8603), .Q (new_AGEMA_signal_8604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_8607), .Q (new_AGEMA_signal_8608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_8611), .Q (new_AGEMA_signal_8612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_8615), .Q (new_AGEMA_signal_8616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_8619), .Q (new_AGEMA_signal_8620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_8623), .Q (new_AGEMA_signal_8624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_8627), .Q (new_AGEMA_signal_8628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_8631), .Q (new_AGEMA_signal_8632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_8635), .Q (new_AGEMA_signal_8636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_8639), .Q (new_AGEMA_signal_8640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_8643), .Q (new_AGEMA_signal_8644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_8647), .Q (new_AGEMA_signal_8648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_8651), .Q (new_AGEMA_signal_8652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_8655), .Q (new_AGEMA_signal_8656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_8659), .Q (new_AGEMA_signal_8660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_8663), .Q (new_AGEMA_signal_8664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_8667), .Q (new_AGEMA_signal_8668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_8671), .Q (new_AGEMA_signal_8672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_8675), .Q (new_AGEMA_signal_8676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_8679), .Q (new_AGEMA_signal_8680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_8683), .Q (new_AGEMA_signal_8684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_8687), .Q (new_AGEMA_signal_8688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_8691), .Q (new_AGEMA_signal_8692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_8695), .Q (new_AGEMA_signal_8696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_8699), .Q (new_AGEMA_signal_8700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_8703), .Q (new_AGEMA_signal_8704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_8707), .Q (new_AGEMA_signal_8708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_8711), .Q (new_AGEMA_signal_8712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_8715), .Q (new_AGEMA_signal_8716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_8719), .Q (new_AGEMA_signal_8720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_8723), .Q (new_AGEMA_signal_8724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_8727), .Q (new_AGEMA_signal_8728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_8731), .Q (new_AGEMA_signal_8732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_8735), .Q (new_AGEMA_signal_8736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_8739), .Q (new_AGEMA_signal_8740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_8743), .Q (new_AGEMA_signal_8744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_8747), .Q (new_AGEMA_signal_8748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_8751), .Q (new_AGEMA_signal_8752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_8755), .Q (new_AGEMA_signal_8756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_8759), .Q (new_AGEMA_signal_8760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_8763), .Q (new_AGEMA_signal_8764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_8767), .Q (new_AGEMA_signal_8768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_8771), .Q (new_AGEMA_signal_8772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_8775), .Q (new_AGEMA_signal_8776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_8779), .Q (new_AGEMA_signal_8780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_8783), .Q (new_AGEMA_signal_8784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_8787), .Q (new_AGEMA_signal_8788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_8791), .Q (new_AGEMA_signal_8792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_8795), .Q (new_AGEMA_signal_8796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_8799), .Q (new_AGEMA_signal_8800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_8803), .Q (new_AGEMA_signal_8804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3771 ( .C (clk), .D (new_AGEMA_signal_8807), .Q (new_AGEMA_signal_8808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_8811), .Q (new_AGEMA_signal_8812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_8815), .Q (new_AGEMA_signal_8816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_8819), .Q (new_AGEMA_signal_8820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_8823), .Q (new_AGEMA_signal_8824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_8827), .Q (new_AGEMA_signal_8828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_8831), .Q (new_AGEMA_signal_8832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_8835), .Q (new_AGEMA_signal_8836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_8839), .Q (new_AGEMA_signal_8840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_8843), .Q (new_AGEMA_signal_8844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_8847), .Q (new_AGEMA_signal_8848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_8851), .Q (new_AGEMA_signal_8852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_8855), .Q (new_AGEMA_signal_8856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_8859), .Q (new_AGEMA_signal_8860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_8863), .Q (new_AGEMA_signal_8864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_8867), .Q (new_AGEMA_signal_8868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_8871), .Q (new_AGEMA_signal_8872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_8875), .Q (new_AGEMA_signal_8876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_8879), .Q (new_AGEMA_signal_8880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_8883), .Q (new_AGEMA_signal_8884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_8887), .Q (new_AGEMA_signal_8888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_8891), .Q (new_AGEMA_signal_8892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_8895), .Q (new_AGEMA_signal_8896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_8899), .Q (new_AGEMA_signal_8900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3867 ( .C (clk), .D (new_AGEMA_signal_8903), .Q (new_AGEMA_signal_8904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_8907), .Q (new_AGEMA_signal_8908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_8911), .Q (new_AGEMA_signal_8912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_8915), .Q (new_AGEMA_signal_8916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_8919), .Q (new_AGEMA_signal_8920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_8923), .Q (new_AGEMA_signal_8924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_8927), .Q (new_AGEMA_signal_8928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_8931), .Q (new_AGEMA_signal_8932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3899 ( .C (clk), .D (new_AGEMA_signal_8935), .Q (new_AGEMA_signal_8936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_8939), .Q (new_AGEMA_signal_8940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_8943), .Q (new_AGEMA_signal_8944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_8947), .Q (new_AGEMA_signal_8948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_8951), .Q (new_AGEMA_signal_8952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_8955), .Q (new_AGEMA_signal_8956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_8959), .Q (new_AGEMA_signal_8960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_8963), .Q (new_AGEMA_signal_8964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_8967), .Q (new_AGEMA_signal_8968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_8971), .Q (new_AGEMA_signal_8972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_8975), .Q (new_AGEMA_signal_8976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_8979), .Q (new_AGEMA_signal_8980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3947 ( .C (clk), .D (new_AGEMA_signal_8983), .Q (new_AGEMA_signal_8984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_8987), .Q (new_AGEMA_signal_8988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_8991), .Q (new_AGEMA_signal_8992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_8995), .Q (new_AGEMA_signal_8996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_8999), .Q (new_AGEMA_signal_9000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_9003), .Q (new_AGEMA_signal_9004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_9007), .Q (new_AGEMA_signal_9008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_9011), .Q (new_AGEMA_signal_9012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_9015), .Q (new_AGEMA_signal_9016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_9019), .Q (new_AGEMA_signal_9020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_9023), .Q (new_AGEMA_signal_9024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_9027), .Q (new_AGEMA_signal_9028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3995 ( .C (clk), .D (new_AGEMA_signal_9031), .Q (new_AGEMA_signal_9032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_9035), .Q (new_AGEMA_signal_9036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_9039), .Q (new_AGEMA_signal_9040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_9043), .Q (new_AGEMA_signal_9044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4011 ( .C (clk), .D (new_AGEMA_signal_9047), .Q (new_AGEMA_signal_9048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_9051), .Q (new_AGEMA_signal_9052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_9055), .Q (new_AGEMA_signal_9056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_9059), .Q (new_AGEMA_signal_9060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_9063), .Q (new_AGEMA_signal_9064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_9067), .Q (new_AGEMA_signal_9068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_9071), .Q (new_AGEMA_signal_9072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_9075), .Q (new_AGEMA_signal_9076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_9079), .Q (new_AGEMA_signal_9080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_9083), .Q (new_AGEMA_signal_9084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_9087), .Q (new_AGEMA_signal_9088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_9091), .Q (new_AGEMA_signal_9092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_9095), .Q (new_AGEMA_signal_9096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_9099), .Q (new_AGEMA_signal_9100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_9103), .Q (new_AGEMA_signal_9104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_9107), .Q (new_AGEMA_signal_9108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_9111), .Q (new_AGEMA_signal_9112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_9115), .Q (new_AGEMA_signal_9116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_9119), .Q (new_AGEMA_signal_9120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_9123), .Q (new_AGEMA_signal_9124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_9127), .Q (new_AGEMA_signal_9128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_9131), .Q (new_AGEMA_signal_9132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_9135), .Q (new_AGEMA_signal_9136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_9139), .Q (new_AGEMA_signal_9140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_9143), .Q (new_AGEMA_signal_9144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_9147), .Q (new_AGEMA_signal_9148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_9151), .Q (new_AGEMA_signal_9152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_9155), .Q (new_AGEMA_signal_9156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_9159), .Q (new_AGEMA_signal_9160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_9163), .Q (new_AGEMA_signal_9164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_9167), .Q (new_AGEMA_signal_9168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_9171), .Q (new_AGEMA_signal_9172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_9175), .Q (new_AGEMA_signal_9176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_9179), .Q (new_AGEMA_signal_9180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_9183), .Q (new_AGEMA_signal_9184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_9187), .Q (new_AGEMA_signal_9188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_9191), .Q (new_AGEMA_signal_9192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_9195), .Q (new_AGEMA_signal_9196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_9199), .Q (new_AGEMA_signal_9200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_9203), .Q (new_AGEMA_signal_9204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_9207), .Q (new_AGEMA_signal_9208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_9211), .Q (new_AGEMA_signal_9212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_9215), .Q (new_AGEMA_signal_9216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_9219), .Q (new_AGEMA_signal_9220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_9223), .Q (new_AGEMA_signal_9224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_9227), .Q (new_AGEMA_signal_9228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_9231), .Q (new_AGEMA_signal_9232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_9235), .Q (new_AGEMA_signal_9236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_9239), .Q (new_AGEMA_signal_9240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_9243), .Q (new_AGEMA_signal_9244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_9247), .Q (new_AGEMA_signal_9248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_9251), .Q (new_AGEMA_signal_9252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_9255), .Q (new_AGEMA_signal_9256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_9259), .Q (new_AGEMA_signal_9260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_9263), .Q (new_AGEMA_signal_9264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_9267), .Q (new_AGEMA_signal_9268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_9271), .Q (new_AGEMA_signal_9272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_9275), .Q (new_AGEMA_signal_9276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_9279), .Q (new_AGEMA_signal_9280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_9283), .Q (new_AGEMA_signal_9284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_9287), .Q (new_AGEMA_signal_9288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_9291), .Q (new_AGEMA_signal_9292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_9295), .Q (new_AGEMA_signal_9296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_9299), .Q (new_AGEMA_signal_9300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_9303), .Q (new_AGEMA_signal_9304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_9307), .Q (new_AGEMA_signal_9308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_9311), .Q (new_AGEMA_signal_9312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_9315), .Q (new_AGEMA_signal_9316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_9319), .Q (new_AGEMA_signal_9320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_9323), .Q (new_AGEMA_signal_9324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_9327), .Q (new_AGEMA_signal_9328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_9331), .Q (new_AGEMA_signal_9332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_9335), .Q (new_AGEMA_signal_9336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_9339), .Q (new_AGEMA_signal_9340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_9343), .Q (new_AGEMA_signal_9344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_9347), .Q (new_AGEMA_signal_9348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_9351), .Q (new_AGEMA_signal_9352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_9355), .Q (new_AGEMA_signal_9356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_9359), .Q (new_AGEMA_signal_9360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_9363), .Q (new_AGEMA_signal_9364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_9367), .Q (new_AGEMA_signal_9368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_9371), .Q (new_AGEMA_signal_9372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_9375), .Q (new_AGEMA_signal_9376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_9379), .Q (new_AGEMA_signal_9380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_9383), .Q (new_AGEMA_signal_9384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_9387), .Q (new_AGEMA_signal_9388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_9391), .Q (new_AGEMA_signal_9392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_9395), .Q (new_AGEMA_signal_9396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_9399), .Q (new_AGEMA_signal_9400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_9403), .Q (new_AGEMA_signal_9404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_9407), .Q (new_AGEMA_signal_9408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_9411), .Q (new_AGEMA_signal_9412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_9415), .Q (new_AGEMA_signal_9416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_9419), .Q (new_AGEMA_signal_9420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_9423), .Q (new_AGEMA_signal_9424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_9427), .Q (new_AGEMA_signal_9428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_9431), .Q (new_AGEMA_signal_9432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_9435), .Q (new_AGEMA_signal_9436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_9439), .Q (new_AGEMA_signal_9440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_9443), .Q (new_AGEMA_signal_9444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_9447), .Q (new_AGEMA_signal_9448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_9451), .Q (new_AGEMA_signal_9452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_9455), .Q (new_AGEMA_signal_9456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_9459), .Q (new_AGEMA_signal_9460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_9463), .Q (new_AGEMA_signal_9464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_9467), .Q (new_AGEMA_signal_9468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_9471), .Q (new_AGEMA_signal_9472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_9475), .Q (new_AGEMA_signal_9476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_9479), .Q (new_AGEMA_signal_9480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_9483), .Q (new_AGEMA_signal_9484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_9487), .Q (new_AGEMA_signal_9488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_9491), .Q (new_AGEMA_signal_9492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_9495), .Q (new_AGEMA_signal_9496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_9499), .Q (new_AGEMA_signal_9500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_9503), .Q (new_AGEMA_signal_9504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_9507), .Q (new_AGEMA_signal_9508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_9511), .Q (new_AGEMA_signal_9512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_9515), .Q (new_AGEMA_signal_9516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_9519), .Q (new_AGEMA_signal_9520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_9523), .Q (new_AGEMA_signal_9524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_9527), .Q (new_AGEMA_signal_9528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_9531), .Q (new_AGEMA_signal_9532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_9535), .Q (new_AGEMA_signal_9536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_9539), .Q (new_AGEMA_signal_9540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_9543), .Q (new_AGEMA_signal_9544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_9547), .Q (new_AGEMA_signal_9548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_9551), .Q (new_AGEMA_signal_9552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_9555), .Q (new_AGEMA_signal_9556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_9559), .Q (new_AGEMA_signal_9560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_9563), .Q (new_AGEMA_signal_9564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_9567), .Q (new_AGEMA_signal_9568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_9571), .Q (new_AGEMA_signal_9572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_9575), .Q (new_AGEMA_signal_9576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_9579), .Q (new_AGEMA_signal_9580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_9583), .Q (new_AGEMA_signal_9584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_9587), .Q (new_AGEMA_signal_9588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_9591), .Q (new_AGEMA_signal_9592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_9595), .Q (new_AGEMA_signal_9596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_9599), .Q (new_AGEMA_signal_9600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_9603), .Q (new_AGEMA_signal_9604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_9607), .Q (new_AGEMA_signal_9608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_9611), .Q (new_AGEMA_signal_9612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_9615), .Q (new_AGEMA_signal_9616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_9619), .Q (new_AGEMA_signal_9620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_9623), .Q (new_AGEMA_signal_9624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_9627), .Q (new_AGEMA_signal_9628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_9631), .Q (new_AGEMA_signal_9632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_9635), .Q (new_AGEMA_signal_9636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_9639), .Q (new_AGEMA_signal_9640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_9643), .Q (new_AGEMA_signal_9644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_9647), .Q (new_AGEMA_signal_9648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_9651), .Q (new_AGEMA_signal_9652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_9655), .Q (new_AGEMA_signal_9656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_9659), .Q (new_AGEMA_signal_9660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_9663), .Q (new_AGEMA_signal_9664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_9667), .Q (new_AGEMA_signal_9668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_9671), .Q (new_AGEMA_signal_9672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_9675), .Q (new_AGEMA_signal_9676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_9679), .Q (new_AGEMA_signal_9680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_9683), .Q (new_AGEMA_signal_9684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_9687), .Q (new_AGEMA_signal_9688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_9691), .Q (new_AGEMA_signal_9692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_9695), .Q (new_AGEMA_signal_9696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_9699), .Q (new_AGEMA_signal_9700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_9703), .Q (new_AGEMA_signal_9704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_9707), .Q (new_AGEMA_signal_9708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_9711), .Q (new_AGEMA_signal_9712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_9715), .Q (new_AGEMA_signal_9716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4683 ( .C (clk), .D (new_AGEMA_signal_9719), .Q (new_AGEMA_signal_9720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_9723), .Q (new_AGEMA_signal_9724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_9727), .Q (new_AGEMA_signal_9728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_9731), .Q (new_AGEMA_signal_9732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_9735), .Q (new_AGEMA_signal_9736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_9739), .Q (new_AGEMA_signal_9740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_9743), .Q (new_AGEMA_signal_9744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_9747), .Q (new_AGEMA_signal_9748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_9751), .Q (new_AGEMA_signal_9752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_9755), .Q (new_AGEMA_signal_9756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_9759), .Q (new_AGEMA_signal_9760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_9763), .Q (new_AGEMA_signal_9764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_9767), .Q (new_AGEMA_signal_9768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_9771), .Q (new_AGEMA_signal_9772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_9775), .Q (new_AGEMA_signal_9776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_9779), .Q (new_AGEMA_signal_9780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_9783), .Q (new_AGEMA_signal_9784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_9787), .Q (new_AGEMA_signal_9788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_9791), .Q (new_AGEMA_signal_9792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_9795), .Q (new_AGEMA_signal_9796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_9799), .Q (new_AGEMA_signal_9800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_9803), .Q (new_AGEMA_signal_9804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_9807), .Q (new_AGEMA_signal_9808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_9811), .Q (new_AGEMA_signal_9812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4779 ( .C (clk), .D (new_AGEMA_signal_9815), .Q (new_AGEMA_signal_9816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_9819), .Q (new_AGEMA_signal_9820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_9823), .Q (new_AGEMA_signal_9824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_9827), .Q (new_AGEMA_signal_9828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_9831), .Q (new_AGEMA_signal_9832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_9835), .Q (new_AGEMA_signal_9836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4803 ( .C (clk), .D (new_AGEMA_signal_9839), .Q (new_AGEMA_signal_9840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_9843), .Q (new_AGEMA_signal_9844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_9847), .Q (new_AGEMA_signal_9848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_9851), .Q (new_AGEMA_signal_9852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_9855), .Q (new_AGEMA_signal_9856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_9859), .Q (new_AGEMA_signal_9860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4827 ( .C (clk), .D (new_AGEMA_signal_9863), .Q (new_AGEMA_signal_9864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_9867), .Q (new_AGEMA_signal_9868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_9871), .Q (new_AGEMA_signal_9872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_9875), .Q (new_AGEMA_signal_9876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_9879), .Q (new_AGEMA_signal_9880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_9883), .Q (new_AGEMA_signal_9884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4851 ( .C (clk), .D (new_AGEMA_signal_9887), .Q (new_AGEMA_signal_9888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_9891), .Q (new_AGEMA_signal_9892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_9895), .Q (new_AGEMA_signal_9896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_9899), .Q (new_AGEMA_signal_9900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_9903), .Q (new_AGEMA_signal_9904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_9907), .Q (new_AGEMA_signal_9908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4875 ( .C (clk), .D (new_AGEMA_signal_9911), .Q (new_AGEMA_signal_9912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_9915), .Q (new_AGEMA_signal_9916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_9919), .Q (new_AGEMA_signal_9920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_9923), .Q (new_AGEMA_signal_9924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_9927), .Q (new_AGEMA_signal_9928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_9931), .Q (new_AGEMA_signal_9932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4899 ( .C (clk), .D (new_AGEMA_signal_9935), .Q (new_AGEMA_signal_9936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_9939), .Q (new_AGEMA_signal_9940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_9943), .Q (new_AGEMA_signal_9944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_9947), .Q (new_AGEMA_signal_9948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_9951), .Q (new_AGEMA_signal_9952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_9955), .Q (new_AGEMA_signal_9956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4923 ( .C (clk), .D (new_AGEMA_signal_9959), .Q (new_AGEMA_signal_9960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_9963), .Q (new_AGEMA_signal_9964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_9967), .Q (new_AGEMA_signal_9968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_9971), .Q (new_AGEMA_signal_9972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_9975), .Q (new_AGEMA_signal_9976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_9979), .Q (new_AGEMA_signal_9980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4947 ( .C (clk), .D (new_AGEMA_signal_9983), .Q (new_AGEMA_signal_9984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_9987), .Q (new_AGEMA_signal_9988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_9991), .Q (new_AGEMA_signal_9992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_9995), .Q (new_AGEMA_signal_9996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_9999), .Q (new_AGEMA_signal_10000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_10003), .Q (new_AGEMA_signal_10004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4971 ( .C (clk), .D (new_AGEMA_signal_10007), .Q (new_AGEMA_signal_10008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_10011), .Q (new_AGEMA_signal_10012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_10015), .Q (new_AGEMA_signal_10016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_10019), .Q (new_AGEMA_signal_10020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_10023), .Q (new_AGEMA_signal_10024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_10027), .Q (new_AGEMA_signal_10028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4995 ( .C (clk), .D (new_AGEMA_signal_10031), .Q (new_AGEMA_signal_10032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_10035), .Q (new_AGEMA_signal_10036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_10039), .Q (new_AGEMA_signal_10040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_10043), .Q (new_AGEMA_signal_10044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_10047), .Q (new_AGEMA_signal_10048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_10051), .Q (new_AGEMA_signal_10052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5019 ( .C (clk), .D (new_AGEMA_signal_10055), .Q (new_AGEMA_signal_10056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_10059), .Q (new_AGEMA_signal_10060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_10063), .Q (new_AGEMA_signal_10064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_10067), .Q (new_AGEMA_signal_10068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_10071), .Q (new_AGEMA_signal_10072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_10075), .Q (new_AGEMA_signal_10076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5043 ( .C (clk), .D (new_AGEMA_signal_10079), .Q (new_AGEMA_signal_10080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_10083), .Q (new_AGEMA_signal_10084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_10087), .Q (new_AGEMA_signal_10088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_10091), .Q (new_AGEMA_signal_10092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_10095), .Q (new_AGEMA_signal_10096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_10099), .Q (new_AGEMA_signal_10100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5067 ( .C (clk), .D (new_AGEMA_signal_10103), .Q (new_AGEMA_signal_10104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_10107), .Q (new_AGEMA_signal_10108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_10111), .Q (new_AGEMA_signal_10112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_10115), .Q (new_AGEMA_signal_10116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_10119), .Q (new_AGEMA_signal_10120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_10123), .Q (new_AGEMA_signal_10124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5091 ( .C (clk), .D (new_AGEMA_signal_10127), .Q (new_AGEMA_signal_10128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_10131), .Q (new_AGEMA_signal_10132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_10135), .Q (new_AGEMA_signal_10136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_10139), .Q (new_AGEMA_signal_10140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_10143), .Q (new_AGEMA_signal_10144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_10147), .Q (new_AGEMA_signal_10148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5115 ( .C (clk), .D (new_AGEMA_signal_10151), .Q (new_AGEMA_signal_10152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_10155), .Q (new_AGEMA_signal_10156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_10159), .Q (new_AGEMA_signal_10160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_10163), .Q (new_AGEMA_signal_10164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_10167), .Q (new_AGEMA_signal_10168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_10171), .Q (new_AGEMA_signal_10172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5139 ( .C (clk), .D (new_AGEMA_signal_10175), .Q (new_AGEMA_signal_10176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_10179), .Q (new_AGEMA_signal_10180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_10183), .Q (new_AGEMA_signal_10184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_10187), .Q (new_AGEMA_signal_10188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_10191), .Q (new_AGEMA_signal_10192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_10195), .Q (new_AGEMA_signal_10196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5163 ( .C (clk), .D (new_AGEMA_signal_10199), .Q (new_AGEMA_signal_10200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_10203), .Q (new_AGEMA_signal_10204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_10207), .Q (new_AGEMA_signal_10208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_10211), .Q (new_AGEMA_signal_10212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_10215), .Q (new_AGEMA_signal_10216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_10219), .Q (new_AGEMA_signal_10220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5187 ( .C (clk), .D (new_AGEMA_signal_10223), .Q (new_AGEMA_signal_10224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_10227), .Q (new_AGEMA_signal_10228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_10231), .Q (new_AGEMA_signal_10232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_10235), .Q (new_AGEMA_signal_10236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_10239), .Q (new_AGEMA_signal_10240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_10243), .Q (new_AGEMA_signal_10244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5211 ( .C (clk), .D (new_AGEMA_signal_10247), .Q (new_AGEMA_signal_10248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_10251), .Q (new_AGEMA_signal_10252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_10255), .Q (new_AGEMA_signal_10256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_10259), .Q (new_AGEMA_signal_10260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_10263), .Q (new_AGEMA_signal_10264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_10267), .Q (new_AGEMA_signal_10268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5235 ( .C (clk), .D (new_AGEMA_signal_10271), .Q (new_AGEMA_signal_10272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_10275), .Q (new_AGEMA_signal_10276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_10279), .Q (new_AGEMA_signal_10280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_10283), .Q (new_AGEMA_signal_10284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_10287), .Q (new_AGEMA_signal_10288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_10291), .Q (new_AGEMA_signal_10292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5259 ( .C (clk), .D (new_AGEMA_signal_10295), .Q (new_AGEMA_signal_10296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_10299), .Q (new_AGEMA_signal_10300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_10303), .Q (new_AGEMA_signal_10304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_10307), .Q (new_AGEMA_signal_10308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_10311), .Q (new_AGEMA_signal_10312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_10315), .Q (new_AGEMA_signal_10316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5283 ( .C (clk), .D (new_AGEMA_signal_10319), .Q (new_AGEMA_signal_10320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_10323), .Q (new_AGEMA_signal_10324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_10327), .Q (new_AGEMA_signal_10328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_10331), .Q (new_AGEMA_signal_10332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_10335), .Q (new_AGEMA_signal_10336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_10339), .Q (new_AGEMA_signal_10340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5307 ( .C (clk), .D (new_AGEMA_signal_10343), .Q (new_AGEMA_signal_10344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_10347), .Q (new_AGEMA_signal_10348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_10351), .Q (new_AGEMA_signal_10352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_10355), .Q (new_AGEMA_signal_10356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_10359), .Q (new_AGEMA_signal_10360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_10363), .Q (new_AGEMA_signal_10364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5331 ( .C (clk), .D (new_AGEMA_signal_10367), .Q (new_AGEMA_signal_10368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_10371), .Q (new_AGEMA_signal_10372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_10375), .Q (new_AGEMA_signal_10376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_10379), .Q (new_AGEMA_signal_10380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_10383), .Q (new_AGEMA_signal_10384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_10387), .Q (new_AGEMA_signal_10388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5355 ( .C (clk), .D (new_AGEMA_signal_10391), .Q (new_AGEMA_signal_10392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_10395), .Q (new_AGEMA_signal_10396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_10399), .Q (new_AGEMA_signal_10400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_10403), .Q (new_AGEMA_signal_10404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_10407), .Q (new_AGEMA_signal_10408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_10411), .Q (new_AGEMA_signal_10412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5379 ( .C (clk), .D (new_AGEMA_signal_10415), .Q (new_AGEMA_signal_10416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_10419), .Q (new_AGEMA_signal_10420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_10423), .Q (new_AGEMA_signal_10424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_10427), .Q (new_AGEMA_signal_10428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_10431), .Q (new_AGEMA_signal_10432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_10435), .Q (new_AGEMA_signal_10436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_10439), .Q (new_AGEMA_signal_10440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_10443), .Q (new_AGEMA_signal_10444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_10447), .Q (new_AGEMA_signal_10448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_10451), .Q (new_AGEMA_signal_10452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_10455), .Q (new_AGEMA_signal_10456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_10459), .Q (new_AGEMA_signal_10460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_10463), .Q (new_AGEMA_signal_10464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_10467), .Q (new_AGEMA_signal_10468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_10471), .Q (new_AGEMA_signal_10472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_10475), .Q (new_AGEMA_signal_10476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_10479), .Q (new_AGEMA_signal_10480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_10483), .Q (new_AGEMA_signal_10484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_10487), .Q (new_AGEMA_signal_10488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_10491), .Q (new_AGEMA_signal_10492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_10495), .Q (new_AGEMA_signal_10496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_10499), .Q (new_AGEMA_signal_10500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_10503), .Q (new_AGEMA_signal_10504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_10507), .Q (new_AGEMA_signal_10508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_10511), .Q (new_AGEMA_signal_10512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_10515), .Q (new_AGEMA_signal_10516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_10519), .Q (new_AGEMA_signal_10520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_10523), .Q (new_AGEMA_signal_10524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_10527), .Q (new_AGEMA_signal_10528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_10531), .Q (new_AGEMA_signal_10532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_10535), .Q (new_AGEMA_signal_10536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_10539), .Q (new_AGEMA_signal_10540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_10543), .Q (new_AGEMA_signal_10544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_10547), .Q (new_AGEMA_signal_10548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_10551), .Q (new_AGEMA_signal_10552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_10555), .Q (new_AGEMA_signal_10556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_10559), .Q (new_AGEMA_signal_10560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_10563), .Q (new_AGEMA_signal_10564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_10567), .Q (new_AGEMA_signal_10568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_10571), .Q (new_AGEMA_signal_10572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_10575), .Q (new_AGEMA_signal_10576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_10579), .Q (new_AGEMA_signal_10580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_10583), .Q (new_AGEMA_signal_10584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_10587), .Q (new_AGEMA_signal_10588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_10591), .Q (new_AGEMA_signal_10592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_10595), .Q (new_AGEMA_signal_10596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_10599), .Q (new_AGEMA_signal_10600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_10603), .Q (new_AGEMA_signal_10604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_10607), .Q (new_AGEMA_signal_10608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_10611), .Q (new_AGEMA_signal_10612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_10615), .Q (new_AGEMA_signal_10616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_10619), .Q (new_AGEMA_signal_10620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_10623), .Q (new_AGEMA_signal_10624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_10627), .Q (new_AGEMA_signal_10628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_10631), .Q (new_AGEMA_signal_10632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_10635), .Q (new_AGEMA_signal_10636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_10639), .Q (new_AGEMA_signal_10640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_10643), .Q (new_AGEMA_signal_10644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_10647), .Q (new_AGEMA_signal_10648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_10651), .Q (new_AGEMA_signal_10652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_10655), .Q (new_AGEMA_signal_10656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_10659), .Q (new_AGEMA_signal_10660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_10663), .Q (new_AGEMA_signal_10664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_10667), .Q (new_AGEMA_signal_10668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_10671), .Q (new_AGEMA_signal_10672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_10675), .Q (new_AGEMA_signal_10676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_10679), .Q (new_AGEMA_signal_10680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_10683), .Q (new_AGEMA_signal_10684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_10687), .Q (new_AGEMA_signal_10688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_10691), .Q (new_AGEMA_signal_10692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_10695), .Q (new_AGEMA_signal_10696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_10699), .Q (new_AGEMA_signal_10700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_10703), .Q (new_AGEMA_signal_10704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_10707), .Q (new_AGEMA_signal_10708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_10711), .Q (new_AGEMA_signal_10712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_10715), .Q (new_AGEMA_signal_10716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_10719), .Q (new_AGEMA_signal_10720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_10723), .Q (new_AGEMA_signal_10724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_10727), .Q (new_AGEMA_signal_10728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_10731), .Q (new_AGEMA_signal_10732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_10735), .Q (new_AGEMA_signal_10736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_10739), .Q (new_AGEMA_signal_10740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_10743), .Q (new_AGEMA_signal_10744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_10747), .Q (new_AGEMA_signal_10748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_10751), .Q (new_AGEMA_signal_10752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_10755), .Q (new_AGEMA_signal_10756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_10759), .Q (new_AGEMA_signal_10760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_10763), .Q (new_AGEMA_signal_10764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_10767), .Q (new_AGEMA_signal_10768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_10771), .Q (new_AGEMA_signal_10772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_10775), .Q (new_AGEMA_signal_10776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_10779), .Q (new_AGEMA_signal_10780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_10783), .Q (new_AGEMA_signal_10784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5751 ( .C (clk), .D (new_AGEMA_signal_10787), .Q (new_AGEMA_signal_10788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_10791), .Q (new_AGEMA_signal_10792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_10795), .Q (new_AGEMA_signal_10796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5763 ( .C (clk), .D (new_AGEMA_signal_10799), .Q (new_AGEMA_signal_10800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_10803), .Q (new_AGEMA_signal_10804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_10807), .Q (new_AGEMA_signal_10808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5775 ( .C (clk), .D (new_AGEMA_signal_10811), .Q (new_AGEMA_signal_10812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_10815), .Q (new_AGEMA_signal_10816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_10819), .Q (new_AGEMA_signal_10820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5787 ( .C (clk), .D (new_AGEMA_signal_10823), .Q (new_AGEMA_signal_10824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_10827), .Q (new_AGEMA_signal_10828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_10831), .Q (new_AGEMA_signal_10832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5799 ( .C (clk), .D (new_AGEMA_signal_10835), .Q (new_AGEMA_signal_10836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_10839), .Q (new_AGEMA_signal_10840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_10843), .Q (new_AGEMA_signal_10844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5811 ( .C (clk), .D (new_AGEMA_signal_10847), .Q (new_AGEMA_signal_10848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_10851), .Q (new_AGEMA_signal_10852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_10855), .Q (new_AGEMA_signal_10856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5823 ( .C (clk), .D (new_AGEMA_signal_10859), .Q (new_AGEMA_signal_10860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_10863), .Q (new_AGEMA_signal_10864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_10867), .Q (new_AGEMA_signal_10868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5835 ( .C (clk), .D (new_AGEMA_signal_10871), .Q (new_AGEMA_signal_10872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_10875), .Q (new_AGEMA_signal_10876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_10879), .Q (new_AGEMA_signal_10880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5847 ( .C (clk), .D (new_AGEMA_signal_10883), .Q (new_AGEMA_signal_10884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_10887), .Q (new_AGEMA_signal_10888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_10891), .Q (new_AGEMA_signal_10892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5859 ( .C (clk), .D (new_AGEMA_signal_10895), .Q (new_AGEMA_signal_10896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_10899), .Q (new_AGEMA_signal_10900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_10903), .Q (new_AGEMA_signal_10904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5871 ( .C (clk), .D (new_AGEMA_signal_10907), .Q (new_AGEMA_signal_10908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_10911), .Q (new_AGEMA_signal_10912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_10915), .Q (new_AGEMA_signal_10916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5883 ( .C (clk), .D (new_AGEMA_signal_10919), .Q (new_AGEMA_signal_10920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_10923), .Q (new_AGEMA_signal_10924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_10927), .Q (new_AGEMA_signal_10928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5895 ( .C (clk), .D (new_AGEMA_signal_10931), .Q (new_AGEMA_signal_10932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_10935), .Q (new_AGEMA_signal_10936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_10939), .Q (new_AGEMA_signal_10940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5907 ( .C (clk), .D (new_AGEMA_signal_10943), .Q (new_AGEMA_signal_10944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_10947), .Q (new_AGEMA_signal_10948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_10951), .Q (new_AGEMA_signal_10952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5919 ( .C (clk), .D (new_AGEMA_signal_10955), .Q (new_AGEMA_signal_10956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_10959), .Q (new_AGEMA_signal_10960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_10963), .Q (new_AGEMA_signal_10964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5931 ( .C (clk), .D (new_AGEMA_signal_10967), .Q (new_AGEMA_signal_10968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_10971), .Q (new_AGEMA_signal_10972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_10975), .Q (new_AGEMA_signal_10976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5943 ( .C (clk), .D (new_AGEMA_signal_10979), .Q (new_AGEMA_signal_10980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_10983), .Q (new_AGEMA_signal_10984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_10987), .Q (new_AGEMA_signal_10988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5955 ( .C (clk), .D (new_AGEMA_signal_10991), .Q (new_AGEMA_signal_10992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_10995), .Q (new_AGEMA_signal_10996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_10999), .Q (new_AGEMA_signal_11000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5967 ( .C (clk), .D (new_AGEMA_signal_11003), .Q (new_AGEMA_signal_11004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_11007), .Q (new_AGEMA_signal_11008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_11011), .Q (new_AGEMA_signal_11012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5979 ( .C (clk), .D (new_AGEMA_signal_11015), .Q (new_AGEMA_signal_11016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_11019), .Q (new_AGEMA_signal_11020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_11023), .Q (new_AGEMA_signal_11024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5991 ( .C (clk), .D (new_AGEMA_signal_11027), .Q (new_AGEMA_signal_11028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_11031), .Q (new_AGEMA_signal_11032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_11035), .Q (new_AGEMA_signal_11036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6003 ( .C (clk), .D (new_AGEMA_signal_11039), .Q (new_AGEMA_signal_11040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_11043), .Q (new_AGEMA_signal_11044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_11047), .Q (new_AGEMA_signal_11048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6015 ( .C (clk), .D (new_AGEMA_signal_11051), .Q (new_AGEMA_signal_11052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_11055), .Q (new_AGEMA_signal_11056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_11059), .Q (new_AGEMA_signal_11060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6027 ( .C (clk), .D (new_AGEMA_signal_11063), .Q (new_AGEMA_signal_11064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_11067), .Q (new_AGEMA_signal_11068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_11071), .Q (new_AGEMA_signal_11072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6039 ( .C (clk), .D (new_AGEMA_signal_11075), .Q (new_AGEMA_signal_11076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_11079), .Q (new_AGEMA_signal_11080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_11083), .Q (new_AGEMA_signal_11084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6051 ( .C (clk), .D (new_AGEMA_signal_11087), .Q (new_AGEMA_signal_11088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6055 ( .C (clk), .D (new_AGEMA_signal_11091), .Q (new_AGEMA_signal_11092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6059 ( .C (clk), .D (new_AGEMA_signal_11095), .Q (new_AGEMA_signal_11096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6063 ( .C (clk), .D (new_AGEMA_signal_11099), .Q (new_AGEMA_signal_11100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6067 ( .C (clk), .D (new_AGEMA_signal_11103), .Q (new_AGEMA_signal_11104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6071 ( .C (clk), .D (new_AGEMA_signal_11107), .Q (new_AGEMA_signal_11108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6075 ( .C (clk), .D (new_AGEMA_signal_11111), .Q (new_AGEMA_signal_11112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6079 ( .C (clk), .D (new_AGEMA_signal_11115), .Q (new_AGEMA_signal_11116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6083 ( .C (clk), .D (new_AGEMA_signal_11119), .Q (new_AGEMA_signal_11120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6087 ( .C (clk), .D (new_AGEMA_signal_11123), .Q (new_AGEMA_signal_11124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6091 ( .C (clk), .D (new_AGEMA_signal_11127), .Q (new_AGEMA_signal_11128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6095 ( .C (clk), .D (new_AGEMA_signal_11131), .Q (new_AGEMA_signal_11132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6099 ( .C (clk), .D (new_AGEMA_signal_11135), .Q (new_AGEMA_signal_11136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6103 ( .C (clk), .D (new_AGEMA_signal_11139), .Q (new_AGEMA_signal_11140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6107 ( .C (clk), .D (new_AGEMA_signal_11143), .Q (new_AGEMA_signal_11144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6111 ( .C (clk), .D (new_AGEMA_signal_11147), .Q (new_AGEMA_signal_11148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6115 ( .C (clk), .D (new_AGEMA_signal_11151), .Q (new_AGEMA_signal_11152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6119 ( .C (clk), .D (new_AGEMA_signal_11155), .Q (new_AGEMA_signal_11156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6123 ( .C (clk), .D (new_AGEMA_signal_11159), .Q (new_AGEMA_signal_11160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6127 ( .C (clk), .D (new_AGEMA_signal_11163), .Q (new_AGEMA_signal_11164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6131 ( .C (clk), .D (new_AGEMA_signal_11167), .Q (new_AGEMA_signal_11168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6135 ( .C (clk), .D (new_AGEMA_signal_11171), .Q (new_AGEMA_signal_11172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6139 ( .C (clk), .D (new_AGEMA_signal_11175), .Q (new_AGEMA_signal_11176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6143 ( .C (clk), .D (new_AGEMA_signal_11179), .Q (new_AGEMA_signal_11180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6147 ( .C (clk), .D (new_AGEMA_signal_11183), .Q (new_AGEMA_signal_11184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6151 ( .C (clk), .D (new_AGEMA_signal_11187), .Q (new_AGEMA_signal_11188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6155 ( .C (clk), .D (new_AGEMA_signal_11191), .Q (new_AGEMA_signal_11192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6159 ( .C (clk), .D (new_AGEMA_signal_11195), .Q (new_AGEMA_signal_11196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6163 ( .C (clk), .D (new_AGEMA_signal_11199), .Q (new_AGEMA_signal_11200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6167 ( .C (clk), .D (new_AGEMA_signal_11203), .Q (new_AGEMA_signal_11204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6171 ( .C (clk), .D (new_AGEMA_signal_11207), .Q (new_AGEMA_signal_11208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6175 ( .C (clk), .D (new_AGEMA_signal_11211), .Q (new_AGEMA_signal_11212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6179 ( .C (clk), .D (new_AGEMA_signal_11215), .Q (new_AGEMA_signal_11216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6183 ( .C (clk), .D (new_AGEMA_signal_11219), .Q (new_AGEMA_signal_11220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6187 ( .C (clk), .D (new_AGEMA_signal_11223), .Q (new_AGEMA_signal_11224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6191 ( .C (clk), .D (new_AGEMA_signal_11227), .Q (new_AGEMA_signal_11228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6195 ( .C (clk), .D (new_AGEMA_signal_11231), .Q (new_AGEMA_signal_11232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6199 ( .C (clk), .D (new_AGEMA_signal_11235), .Q (new_AGEMA_signal_11236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6203 ( .C (clk), .D (new_AGEMA_signal_11239), .Q (new_AGEMA_signal_11240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6207 ( .C (clk), .D (new_AGEMA_signal_11243), .Q (new_AGEMA_signal_11244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6211 ( .C (clk), .D (new_AGEMA_signal_11247), .Q (new_AGEMA_signal_11248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6215 ( .C (clk), .D (new_AGEMA_signal_11251), .Q (new_AGEMA_signal_11252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6219 ( .C (clk), .D (new_AGEMA_signal_11255), .Q (new_AGEMA_signal_11256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6223 ( .C (clk), .D (new_AGEMA_signal_11259), .Q (new_AGEMA_signal_11260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6227 ( .C (clk), .D (new_AGEMA_signal_11263), .Q (new_AGEMA_signal_11264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6231 ( .C (clk), .D (new_AGEMA_signal_11267), .Q (new_AGEMA_signal_11268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6235 ( .C (clk), .D (new_AGEMA_signal_11271), .Q (new_AGEMA_signal_11272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6239 ( .C (clk), .D (new_AGEMA_signal_11275), .Q (new_AGEMA_signal_11276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6243 ( .C (clk), .D (new_AGEMA_signal_11279), .Q (new_AGEMA_signal_11280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6247 ( .C (clk), .D (new_AGEMA_signal_11283), .Q (new_AGEMA_signal_11284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6251 ( .C (clk), .D (new_AGEMA_signal_11287), .Q (new_AGEMA_signal_11288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6255 ( .C (clk), .D (new_AGEMA_signal_11291), .Q (new_AGEMA_signal_11292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6259 ( .C (clk), .D (new_AGEMA_signal_11295), .Q (new_AGEMA_signal_11296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6263 ( .C (clk), .D (new_AGEMA_signal_11299), .Q (new_AGEMA_signal_11300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6267 ( .C (clk), .D (new_AGEMA_signal_11303), .Q (new_AGEMA_signal_11304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6271 ( .C (clk), .D (new_AGEMA_signal_11307), .Q (new_AGEMA_signal_11308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6275 ( .C (clk), .D (new_AGEMA_signal_11311), .Q (new_AGEMA_signal_11312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6279 ( .C (clk), .D (new_AGEMA_signal_11315), .Q (new_AGEMA_signal_11316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6283 ( .C (clk), .D (new_AGEMA_signal_11319), .Q (new_AGEMA_signal_11320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6287 ( .C (clk), .D (new_AGEMA_signal_11323), .Q (new_AGEMA_signal_11324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6291 ( .C (clk), .D (new_AGEMA_signal_11327), .Q (new_AGEMA_signal_11328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6295 ( .C (clk), .D (new_AGEMA_signal_11331), .Q (new_AGEMA_signal_11332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6299 ( .C (clk), .D (new_AGEMA_signal_11335), .Q (new_AGEMA_signal_11336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6303 ( .C (clk), .D (new_AGEMA_signal_11339), .Q (new_AGEMA_signal_11340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6307 ( .C (clk), .D (new_AGEMA_signal_11343), .Q (new_AGEMA_signal_11344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6311 ( .C (clk), .D (new_AGEMA_signal_11347), .Q (new_AGEMA_signal_11348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6315 ( .C (clk), .D (new_AGEMA_signal_11351), .Q (new_AGEMA_signal_11352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6319 ( .C (clk), .D (new_AGEMA_signal_11355), .Q (new_AGEMA_signal_11356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6323 ( .C (clk), .D (new_AGEMA_signal_11359), .Q (new_AGEMA_signal_11360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6327 ( .C (clk), .D (new_AGEMA_signal_11363), .Q (new_AGEMA_signal_11364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6331 ( .C (clk), .D (new_AGEMA_signal_11367), .Q (new_AGEMA_signal_11368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6335 ( .C (clk), .D (new_AGEMA_signal_11371), .Q (new_AGEMA_signal_11372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6339 ( .C (clk), .D (new_AGEMA_signal_11375), .Q (new_AGEMA_signal_11376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6343 ( .C (clk), .D (new_AGEMA_signal_11379), .Q (new_AGEMA_signal_11380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6347 ( .C (clk), .D (new_AGEMA_signal_11383), .Q (new_AGEMA_signal_11384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6351 ( .C (clk), .D (new_AGEMA_signal_11387), .Q (new_AGEMA_signal_11388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6355 ( .C (clk), .D (new_AGEMA_signal_11391), .Q (new_AGEMA_signal_11392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6359 ( .C (clk), .D (new_AGEMA_signal_11395), .Q (new_AGEMA_signal_11396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6363 ( .C (clk), .D (new_AGEMA_signal_11399), .Q (new_AGEMA_signal_11400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6367 ( .C (clk), .D (new_AGEMA_signal_11403), .Q (new_AGEMA_signal_11404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6371 ( .C (clk), .D (new_AGEMA_signal_11407), .Q (new_AGEMA_signal_11408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6375 ( .C (clk), .D (new_AGEMA_signal_11411), .Q (new_AGEMA_signal_11412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6379 ( .C (clk), .D (new_AGEMA_signal_11415), .Q (new_AGEMA_signal_11416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6383 ( .C (clk), .D (new_AGEMA_signal_11419), .Q (new_AGEMA_signal_11420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6387 ( .C (clk), .D (new_AGEMA_signal_11423), .Q (new_AGEMA_signal_11424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6391 ( .C (clk), .D (new_AGEMA_signal_11427), .Q (new_AGEMA_signal_11428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6395 ( .C (clk), .D (new_AGEMA_signal_11431), .Q (new_AGEMA_signal_11432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6399 ( .C (clk), .D (new_AGEMA_signal_11435), .Q (new_AGEMA_signal_11436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6403 ( .C (clk), .D (new_AGEMA_signal_11439), .Q (new_AGEMA_signal_11440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6407 ( .C (clk), .D (new_AGEMA_signal_11443), .Q (new_AGEMA_signal_11444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6411 ( .C (clk), .D (new_AGEMA_signal_11447), .Q (new_AGEMA_signal_11448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6415 ( .C (clk), .D (new_AGEMA_signal_11451), .Q (new_AGEMA_signal_11452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6419 ( .C (clk), .D (new_AGEMA_signal_11455), .Q (new_AGEMA_signal_11456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6423 ( .C (clk), .D (new_AGEMA_signal_11459), .Q (new_AGEMA_signal_11460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6427 ( .C (clk), .D (new_AGEMA_signal_11463), .Q (new_AGEMA_signal_11464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6431 ( .C (clk), .D (new_AGEMA_signal_11467), .Q (new_AGEMA_signal_11468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6435 ( .C (clk), .D (new_AGEMA_signal_11471), .Q (new_AGEMA_signal_11472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6439 ( .C (clk), .D (new_AGEMA_signal_11475), .Q (new_AGEMA_signal_11476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6443 ( .C (clk), .D (new_AGEMA_signal_11479), .Q (new_AGEMA_signal_11480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6447 ( .C (clk), .D (new_AGEMA_signal_11483), .Q (new_AGEMA_signal_11484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6451 ( .C (clk), .D (new_AGEMA_signal_11487), .Q (new_AGEMA_signal_11488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6455 ( .C (clk), .D (new_AGEMA_signal_11491), .Q (new_AGEMA_signal_11492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6459 ( .C (clk), .D (new_AGEMA_signal_11495), .Q (new_AGEMA_signal_11496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6463 ( .C (clk), .D (new_AGEMA_signal_11499), .Q (new_AGEMA_signal_11500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6467 ( .C (clk), .D (new_AGEMA_signal_11503), .Q (new_AGEMA_signal_11504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6471 ( .C (clk), .D (new_AGEMA_signal_11507), .Q (new_AGEMA_signal_11508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6475 ( .C (clk), .D (new_AGEMA_signal_11511), .Q (new_AGEMA_signal_11512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6479 ( .C (clk), .D (new_AGEMA_signal_11515), .Q (new_AGEMA_signal_11516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6483 ( .C (clk), .D (new_AGEMA_signal_11519), .Q (new_AGEMA_signal_11520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6487 ( .C (clk), .D (new_AGEMA_signal_11523), .Q (new_AGEMA_signal_11524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6491 ( .C (clk), .D (new_AGEMA_signal_11527), .Q (new_AGEMA_signal_11528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6495 ( .C (clk), .D (new_AGEMA_signal_11531), .Q (new_AGEMA_signal_11532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6499 ( .C (clk), .D (new_AGEMA_signal_11535), .Q (new_AGEMA_signal_11536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6503 ( .C (clk), .D (new_AGEMA_signal_11539), .Q (new_AGEMA_signal_11540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6507 ( .C (clk), .D (new_AGEMA_signal_11543), .Q (new_AGEMA_signal_11544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6511 ( .C (clk), .D (new_AGEMA_signal_11547), .Q (new_AGEMA_signal_11548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6515 ( .C (clk), .D (new_AGEMA_signal_11551), .Q (new_AGEMA_signal_11552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6519 ( .C (clk), .D (new_AGEMA_signal_11555), .Q (new_AGEMA_signal_11556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6523 ( .C (clk), .D (new_AGEMA_signal_11559), .Q (new_AGEMA_signal_11560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6527 ( .C (clk), .D (new_AGEMA_signal_11563), .Q (new_AGEMA_signal_11564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6531 ( .C (clk), .D (new_AGEMA_signal_11567), .Q (new_AGEMA_signal_11568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6535 ( .C (clk), .D (new_AGEMA_signal_11571), .Q (new_AGEMA_signal_11572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6539 ( .C (clk), .D (new_AGEMA_signal_11575), .Q (new_AGEMA_signal_11576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6543 ( .C (clk), .D (new_AGEMA_signal_11579), .Q (new_AGEMA_signal_11580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6547 ( .C (clk), .D (new_AGEMA_signal_11583), .Q (new_AGEMA_signal_11584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6551 ( .C (clk), .D (new_AGEMA_signal_11587), .Q (new_AGEMA_signal_11588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6555 ( .C (clk), .D (new_AGEMA_signal_11591), .Q (new_AGEMA_signal_11592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6559 ( .C (clk), .D (new_AGEMA_signal_11595), .Q (new_AGEMA_signal_11596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6563 ( .C (clk), .D (new_AGEMA_signal_11599), .Q (new_AGEMA_signal_11600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6567 ( .C (clk), .D (new_AGEMA_signal_11603), .Q (new_AGEMA_signal_11604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6571 ( .C (clk), .D (new_AGEMA_signal_11607), .Q (new_AGEMA_signal_11608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6575 ( .C (clk), .D (new_AGEMA_signal_11611), .Q (new_AGEMA_signal_11612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6579 ( .C (clk), .D (new_AGEMA_signal_11615), .Q (new_AGEMA_signal_11616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6583 ( .C (clk), .D (new_AGEMA_signal_11619), .Q (new_AGEMA_signal_11620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6587 ( .C (clk), .D (new_AGEMA_signal_11623), .Q (new_AGEMA_signal_11624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6591 ( .C (clk), .D (new_AGEMA_signal_11627), .Q (new_AGEMA_signal_11628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6595 ( .C (clk), .D (new_AGEMA_signal_11631), .Q (new_AGEMA_signal_11632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6599 ( .C (clk), .D (new_AGEMA_signal_11635), .Q (new_AGEMA_signal_11636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6603 ( .C (clk), .D (new_AGEMA_signal_11639), .Q (new_AGEMA_signal_11640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6607 ( .C (clk), .D (new_AGEMA_signal_11643), .Q (new_AGEMA_signal_11644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6611 ( .C (clk), .D (new_AGEMA_signal_11647), .Q (new_AGEMA_signal_11648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6615 ( .C (clk), .D (new_AGEMA_signal_11651), .Q (new_AGEMA_signal_11652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6619 ( .C (clk), .D (new_AGEMA_signal_11655), .Q (new_AGEMA_signal_11656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6623 ( .C (clk), .D (new_AGEMA_signal_11659), .Q (new_AGEMA_signal_11660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6627 ( .C (clk), .D (new_AGEMA_signal_11663), .Q (new_AGEMA_signal_11664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6631 ( .C (clk), .D (new_AGEMA_signal_11667), .Q (new_AGEMA_signal_11668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6635 ( .C (clk), .D (new_AGEMA_signal_11671), .Q (new_AGEMA_signal_11672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6639 ( .C (clk), .D (new_AGEMA_signal_11675), .Q (new_AGEMA_signal_11676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6643 ( .C (clk), .D (new_AGEMA_signal_11679), .Q (new_AGEMA_signal_11680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6647 ( .C (clk), .D (new_AGEMA_signal_11683), .Q (new_AGEMA_signal_11684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6651 ( .C (clk), .D (new_AGEMA_signal_11687), .Q (new_AGEMA_signal_11688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6655 ( .C (clk), .D (new_AGEMA_signal_11691), .Q (new_AGEMA_signal_11692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6659 ( .C (clk), .D (new_AGEMA_signal_11695), .Q (new_AGEMA_signal_11696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6663 ( .C (clk), .D (new_AGEMA_signal_11699), .Q (new_AGEMA_signal_11700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6667 ( .C (clk), .D (new_AGEMA_signal_11703), .Q (new_AGEMA_signal_11704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6671 ( .C (clk), .D (new_AGEMA_signal_11707), .Q (new_AGEMA_signal_11708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6675 ( .C (clk), .D (new_AGEMA_signal_11711), .Q (new_AGEMA_signal_11712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6679 ( .C (clk), .D (new_AGEMA_signal_11715), .Q (new_AGEMA_signal_11716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6683 ( .C (clk), .D (new_AGEMA_signal_11719), .Q (new_AGEMA_signal_11720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6687 ( .C (clk), .D (new_AGEMA_signal_11723), .Q (new_AGEMA_signal_11724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6691 ( .C (clk), .D (new_AGEMA_signal_11727), .Q (new_AGEMA_signal_11728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6695 ( .C (clk), .D (new_AGEMA_signal_11731), .Q (new_AGEMA_signal_11732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6699 ( .C (clk), .D (new_AGEMA_signal_11735), .Q (new_AGEMA_signal_11736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6703 ( .C (clk), .D (new_AGEMA_signal_11739), .Q (new_AGEMA_signal_11740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6707 ( .C (clk), .D (new_AGEMA_signal_11743), .Q (new_AGEMA_signal_11744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6711 ( .C (clk), .D (new_AGEMA_signal_11747), .Q (new_AGEMA_signal_11748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6715 ( .C (clk), .D (new_AGEMA_signal_11751), .Q (new_AGEMA_signal_11752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6719 ( .C (clk), .D (new_AGEMA_signal_11755), .Q (new_AGEMA_signal_11756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6723 ( .C (clk), .D (new_AGEMA_signal_11759), .Q (new_AGEMA_signal_11760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6727 ( .C (clk), .D (new_AGEMA_signal_11763), .Q (new_AGEMA_signal_11764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6731 ( .C (clk), .D (new_AGEMA_signal_11767), .Q (new_AGEMA_signal_11768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6735 ( .C (clk), .D (new_AGEMA_signal_11771), .Q (new_AGEMA_signal_11772) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C (clk), .D (new_AGEMA_signal_11775), .Q (new_AGEMA_signal_11776) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C (clk), .D (new_AGEMA_signal_11779), .Q (new_AGEMA_signal_11780) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C (clk), .D (new_AGEMA_signal_11783), .Q (new_AGEMA_signal_11784) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C (clk), .D (new_AGEMA_signal_11787), .Q (new_AGEMA_signal_11788) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C (clk), .D (new_AGEMA_signal_11791), .Q (new_AGEMA_signal_11792) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C (clk), .D (new_AGEMA_signal_11795), .Q (new_AGEMA_signal_11796) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C (clk), .D (new_AGEMA_signal_11799), .Q (new_AGEMA_signal_11800) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C (clk), .D (new_AGEMA_signal_11803), .Q (new_AGEMA_signal_11804) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C (clk), .D (new_AGEMA_signal_11807), .Q (new_AGEMA_signal_11808) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C (clk), .D (new_AGEMA_signal_11811), .Q (new_AGEMA_signal_11812) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C (clk), .D (new_AGEMA_signal_11815), .Q (new_AGEMA_signal_11816) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C (clk), .D (new_AGEMA_signal_11819), .Q (new_AGEMA_signal_11820) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C (clk), .D (new_AGEMA_signal_11823), .Q (new_AGEMA_signal_11824) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C (clk), .D (new_AGEMA_signal_11827), .Q (new_AGEMA_signal_11828) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C (clk), .D (new_AGEMA_signal_11831), .Q (new_AGEMA_signal_11832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6799 ( .C (clk), .D (new_AGEMA_signal_11835), .Q (new_AGEMA_signal_11836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6803 ( .C (clk), .D (new_AGEMA_signal_11839), .Q (new_AGEMA_signal_11840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6807 ( .C (clk), .D (new_AGEMA_signal_11843), .Q (new_AGEMA_signal_11844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6811 ( .C (clk), .D (new_AGEMA_signal_11847), .Q (new_AGEMA_signal_11848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6815 ( .C (clk), .D (new_AGEMA_signal_11851), .Q (new_AGEMA_signal_11852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6819 ( .C (clk), .D (new_AGEMA_signal_11855), .Q (new_AGEMA_signal_11856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6823 ( .C (clk), .D (new_AGEMA_signal_11859), .Q (new_AGEMA_signal_11860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6827 ( .C (clk), .D (new_AGEMA_signal_11863), .Q (new_AGEMA_signal_11864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6831 ( .C (clk), .D (new_AGEMA_signal_11867), .Q (new_AGEMA_signal_11868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6835 ( .C (clk), .D (new_AGEMA_signal_11871), .Q (new_AGEMA_signal_11872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6839 ( .C (clk), .D (new_AGEMA_signal_11875), .Q (new_AGEMA_signal_11876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6843 ( .C (clk), .D (new_AGEMA_signal_11879), .Q (new_AGEMA_signal_11880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6847 ( .C (clk), .D (new_AGEMA_signal_11883), .Q (new_AGEMA_signal_11884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6851 ( .C (clk), .D (new_AGEMA_signal_11887), .Q (new_AGEMA_signal_11888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6855 ( .C (clk), .D (new_AGEMA_signal_11891), .Q (new_AGEMA_signal_11892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6859 ( .C (clk), .D (new_AGEMA_signal_11895), .Q (new_AGEMA_signal_11896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6863 ( .C (clk), .D (new_AGEMA_signal_11899), .Q (new_AGEMA_signal_11900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6867 ( .C (clk), .D (new_AGEMA_signal_11903), .Q (new_AGEMA_signal_11904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6871 ( .C (clk), .D (new_AGEMA_signal_11907), .Q (new_AGEMA_signal_11908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6875 ( .C (clk), .D (new_AGEMA_signal_11911), .Q (new_AGEMA_signal_11912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6879 ( .C (clk), .D (new_AGEMA_signal_11915), .Q (new_AGEMA_signal_11916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6883 ( .C (clk), .D (new_AGEMA_signal_11919), .Q (new_AGEMA_signal_11920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6887 ( .C (clk), .D (new_AGEMA_signal_11923), .Q (new_AGEMA_signal_11924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6891 ( .C (clk), .D (new_AGEMA_signal_11927), .Q (new_AGEMA_signal_11928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6895 ( .C (clk), .D (new_AGEMA_signal_11931), .Q (new_AGEMA_signal_11932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6899 ( .C (clk), .D (new_AGEMA_signal_11935), .Q (new_AGEMA_signal_11936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6903 ( .C (clk), .D (new_AGEMA_signal_11939), .Q (new_AGEMA_signal_11940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6907 ( .C (clk), .D (new_AGEMA_signal_11943), .Q (new_AGEMA_signal_11944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6911 ( .C (clk), .D (new_AGEMA_signal_11947), .Q (new_AGEMA_signal_11948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6915 ( .C (clk), .D (new_AGEMA_signal_11951), .Q (new_AGEMA_signal_11952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6919 ( .C (clk), .D (new_AGEMA_signal_11955), .Q (new_AGEMA_signal_11956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6923 ( .C (clk), .D (new_AGEMA_signal_11959), .Q (new_AGEMA_signal_11960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6927 ( .C (clk), .D (new_AGEMA_signal_11963), .Q (new_AGEMA_signal_11964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6931 ( .C (clk), .D (new_AGEMA_signal_11967), .Q (new_AGEMA_signal_11968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6935 ( .C (clk), .D (new_AGEMA_signal_11971), .Q (new_AGEMA_signal_11972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6939 ( .C (clk), .D (new_AGEMA_signal_11975), .Q (new_AGEMA_signal_11976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6943 ( .C (clk), .D (new_AGEMA_signal_11979), .Q (new_AGEMA_signal_11980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6947 ( .C (clk), .D (new_AGEMA_signal_11983), .Q (new_AGEMA_signal_11984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6951 ( .C (clk), .D (new_AGEMA_signal_11987), .Q (new_AGEMA_signal_11988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6955 ( .C (clk), .D (new_AGEMA_signal_11991), .Q (new_AGEMA_signal_11992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6959 ( .C (clk), .D (new_AGEMA_signal_11995), .Q (new_AGEMA_signal_11996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6963 ( .C (clk), .D (new_AGEMA_signal_11999), .Q (new_AGEMA_signal_12000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6967 ( .C (clk), .D (new_AGEMA_signal_12003), .Q (new_AGEMA_signal_12004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6971 ( .C (clk), .D (new_AGEMA_signal_12007), .Q (new_AGEMA_signal_12008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6975 ( .C (clk), .D (new_AGEMA_signal_12011), .Q (new_AGEMA_signal_12012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6979 ( .C (clk), .D (new_AGEMA_signal_12015), .Q (new_AGEMA_signal_12016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6983 ( .C (clk), .D (new_AGEMA_signal_12019), .Q (new_AGEMA_signal_12020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6987 ( .C (clk), .D (new_AGEMA_signal_12023), .Q (new_AGEMA_signal_12024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6991 ( .C (clk), .D (new_AGEMA_signal_12027), .Q (new_AGEMA_signal_12028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6995 ( .C (clk), .D (new_AGEMA_signal_12031), .Q (new_AGEMA_signal_12032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6999 ( .C (clk), .D (new_AGEMA_signal_12035), .Q (new_AGEMA_signal_12036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7003 ( .C (clk), .D (new_AGEMA_signal_12039), .Q (new_AGEMA_signal_12040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7007 ( .C (clk), .D (new_AGEMA_signal_12043), .Q (new_AGEMA_signal_12044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7011 ( .C (clk), .D (new_AGEMA_signal_12047), .Q (new_AGEMA_signal_12048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7015 ( .C (clk), .D (new_AGEMA_signal_12051), .Q (new_AGEMA_signal_12052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7019 ( .C (clk), .D (new_AGEMA_signal_12055), .Q (new_AGEMA_signal_12056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7023 ( .C (clk), .D (new_AGEMA_signal_12059), .Q (new_AGEMA_signal_12060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7027 ( .C (clk), .D (new_AGEMA_signal_12063), .Q (new_AGEMA_signal_12064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7031 ( .C (clk), .D (new_AGEMA_signal_12067), .Q (new_AGEMA_signal_12068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7035 ( .C (clk), .D (new_AGEMA_signal_12071), .Q (new_AGEMA_signal_12072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7039 ( .C (clk), .D (new_AGEMA_signal_12075), .Q (new_AGEMA_signal_12076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7043 ( .C (clk), .D (new_AGEMA_signal_12079), .Q (new_AGEMA_signal_12080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7047 ( .C (clk), .D (new_AGEMA_signal_12083), .Q (new_AGEMA_signal_12084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7051 ( .C (clk), .D (new_AGEMA_signal_12087), .Q (new_AGEMA_signal_12088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7055 ( .C (clk), .D (new_AGEMA_signal_12091), .Q (new_AGEMA_signal_12092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7059 ( .C (clk), .D (new_AGEMA_signal_12095), .Q (new_AGEMA_signal_12096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7063 ( .C (clk), .D (new_AGEMA_signal_12099), .Q (new_AGEMA_signal_12100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7067 ( .C (clk), .D (new_AGEMA_signal_12103), .Q (new_AGEMA_signal_12104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7071 ( .C (clk), .D (new_AGEMA_signal_12107), .Q (new_AGEMA_signal_12108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7075 ( .C (clk), .D (new_AGEMA_signal_12111), .Q (new_AGEMA_signal_12112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7079 ( .C (clk), .D (new_AGEMA_signal_12115), .Q (new_AGEMA_signal_12116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7083 ( .C (clk), .D (new_AGEMA_signal_12119), .Q (new_AGEMA_signal_12120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7087 ( .C (clk), .D (new_AGEMA_signal_12123), .Q (new_AGEMA_signal_12124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7091 ( .C (clk), .D (new_AGEMA_signal_12127), .Q (new_AGEMA_signal_12128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7095 ( .C (clk), .D (new_AGEMA_signal_12131), .Q (new_AGEMA_signal_12132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7099 ( .C (clk), .D (new_AGEMA_signal_12135), .Q (new_AGEMA_signal_12136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7103 ( .C (clk), .D (new_AGEMA_signal_12139), .Q (new_AGEMA_signal_12140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7107 ( .C (clk), .D (new_AGEMA_signal_12143), .Q (new_AGEMA_signal_12144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7111 ( .C (clk), .D (new_AGEMA_signal_12147), .Q (new_AGEMA_signal_12148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7115 ( .C (clk), .D (new_AGEMA_signal_12151), .Q (new_AGEMA_signal_12152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7119 ( .C (clk), .D (new_AGEMA_signal_12155), .Q (new_AGEMA_signal_12156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7123 ( .C (clk), .D (new_AGEMA_signal_12159), .Q (new_AGEMA_signal_12160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7127 ( .C (clk), .D (new_AGEMA_signal_12163), .Q (new_AGEMA_signal_12164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7131 ( .C (clk), .D (new_AGEMA_signal_12167), .Q (new_AGEMA_signal_12168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7135 ( .C (clk), .D (new_AGEMA_signal_12171), .Q (new_AGEMA_signal_12172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7139 ( .C (clk), .D (new_AGEMA_signal_12175), .Q (new_AGEMA_signal_12176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7143 ( .C (clk), .D (new_AGEMA_signal_12179), .Q (new_AGEMA_signal_12180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7147 ( .C (clk), .D (new_AGEMA_signal_12183), .Q (new_AGEMA_signal_12184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7151 ( .C (clk), .D (new_AGEMA_signal_12187), .Q (new_AGEMA_signal_12188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7155 ( .C (clk), .D (new_AGEMA_signal_12191), .Q (new_AGEMA_signal_12192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7159 ( .C (clk), .D (new_AGEMA_signal_12195), .Q (new_AGEMA_signal_12196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7163 ( .C (clk), .D (new_AGEMA_signal_12199), .Q (new_AGEMA_signal_12200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7167 ( .C (clk), .D (new_AGEMA_signal_12203), .Q (new_AGEMA_signal_12204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7171 ( .C (clk), .D (new_AGEMA_signal_12207), .Q (new_AGEMA_signal_12208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7175 ( .C (clk), .D (new_AGEMA_signal_12211), .Q (new_AGEMA_signal_12212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7179 ( .C (clk), .D (new_AGEMA_signal_12215), .Q (new_AGEMA_signal_12216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7183 ( .C (clk), .D (new_AGEMA_signal_12219), .Q (new_AGEMA_signal_12220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7187 ( .C (clk), .D (new_AGEMA_signal_12223), .Q (new_AGEMA_signal_12224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7191 ( .C (clk), .D (new_AGEMA_signal_12227), .Q (new_AGEMA_signal_12228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7195 ( .C (clk), .D (new_AGEMA_signal_12231), .Q (new_AGEMA_signal_12232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7199 ( .C (clk), .D (new_AGEMA_signal_12235), .Q (new_AGEMA_signal_12236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7203 ( .C (clk), .D (new_AGEMA_signal_12239), .Q (new_AGEMA_signal_12240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7207 ( .C (clk), .D (new_AGEMA_signal_12243), .Q (new_AGEMA_signal_12244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7211 ( .C (clk), .D (new_AGEMA_signal_12247), .Q (new_AGEMA_signal_12248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7215 ( .C (clk), .D (new_AGEMA_signal_12251), .Q (new_AGEMA_signal_12252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7219 ( .C (clk), .D (new_AGEMA_signal_12255), .Q (new_AGEMA_signal_12256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7223 ( .C (clk), .D (new_AGEMA_signal_12259), .Q (new_AGEMA_signal_12260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7227 ( .C (clk), .D (new_AGEMA_signal_12263), .Q (new_AGEMA_signal_12264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7231 ( .C (clk), .D (new_AGEMA_signal_12267), .Q (new_AGEMA_signal_12268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7235 ( .C (clk), .D (new_AGEMA_signal_12271), .Q (new_AGEMA_signal_12272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7239 ( .C (clk), .D (new_AGEMA_signal_12275), .Q (new_AGEMA_signal_12276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7243 ( .C (clk), .D (new_AGEMA_signal_12279), .Q (new_AGEMA_signal_12280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7247 ( .C (clk), .D (new_AGEMA_signal_12283), .Q (new_AGEMA_signal_12284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7251 ( .C (clk), .D (new_AGEMA_signal_12287), .Q (new_AGEMA_signal_12288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7255 ( .C (clk), .D (new_AGEMA_signal_12291), .Q (new_AGEMA_signal_12292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7259 ( .C (clk), .D (new_AGEMA_signal_12295), .Q (new_AGEMA_signal_12296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7263 ( .C (clk), .D (new_AGEMA_signal_12299), .Q (new_AGEMA_signal_12300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7267 ( .C (clk), .D (new_AGEMA_signal_12303), .Q (new_AGEMA_signal_12304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7271 ( .C (clk), .D (new_AGEMA_signal_12307), .Q (new_AGEMA_signal_12308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7275 ( .C (clk), .D (new_AGEMA_signal_12311), .Q (new_AGEMA_signal_12312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7279 ( .C (clk), .D (new_AGEMA_signal_12315), .Q (new_AGEMA_signal_12316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7283 ( .C (clk), .D (new_AGEMA_signal_12319), .Q (new_AGEMA_signal_12320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7287 ( .C (clk), .D (new_AGEMA_signal_12323), .Q (new_AGEMA_signal_12324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7291 ( .C (clk), .D (new_AGEMA_signal_12327), .Q (new_AGEMA_signal_12328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7295 ( .C (clk), .D (new_AGEMA_signal_12331), .Q (new_AGEMA_signal_12332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7299 ( .C (clk), .D (new_AGEMA_signal_12335), .Q (new_AGEMA_signal_12336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7303 ( .C (clk), .D (new_AGEMA_signal_12339), .Q (new_AGEMA_signal_12340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7307 ( .C (clk), .D (new_AGEMA_signal_12343), .Q (new_AGEMA_signal_12344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7311 ( .C (clk), .D (new_AGEMA_signal_12347), .Q (new_AGEMA_signal_12348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7315 ( .C (clk), .D (new_AGEMA_signal_12351), .Q (new_AGEMA_signal_12352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7319 ( .C (clk), .D (new_AGEMA_signal_12355), .Q (new_AGEMA_signal_12356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7323 ( .C (clk), .D (new_AGEMA_signal_12359), .Q (new_AGEMA_signal_12360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7327 ( .C (clk), .D (new_AGEMA_signal_12363), .Q (new_AGEMA_signal_12364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7331 ( .C (clk), .D (new_AGEMA_signal_12367), .Q (new_AGEMA_signal_12368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7335 ( .C (clk), .D (new_AGEMA_signal_12371), .Q (new_AGEMA_signal_12372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7339 ( .C (clk), .D (new_AGEMA_signal_12375), .Q (new_AGEMA_signal_12376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7343 ( .C (clk), .D (new_AGEMA_signal_12379), .Q (new_AGEMA_signal_12380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7347 ( .C (clk), .D (new_AGEMA_signal_12383), .Q (new_AGEMA_signal_12384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7351 ( .C (clk), .D (new_AGEMA_signal_12387), .Q (new_AGEMA_signal_12388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7355 ( .C (clk), .D (new_AGEMA_signal_12391), .Q (new_AGEMA_signal_12392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7359 ( .C (clk), .D (new_AGEMA_signal_12395), .Q (new_AGEMA_signal_12396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7363 ( .C (clk), .D (new_AGEMA_signal_12399), .Q (new_AGEMA_signal_12400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7367 ( .C (clk), .D (new_AGEMA_signal_12403), .Q (new_AGEMA_signal_12404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7371 ( .C (clk), .D (new_AGEMA_signal_12407), .Q (new_AGEMA_signal_12408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7375 ( .C (clk), .D (new_AGEMA_signal_12411), .Q (new_AGEMA_signal_12412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7379 ( .C (clk), .D (new_AGEMA_signal_12415), .Q (new_AGEMA_signal_12416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7383 ( .C (clk), .D (new_AGEMA_signal_12419), .Q (new_AGEMA_signal_12420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7387 ( .C (clk), .D (new_AGEMA_signal_12423), .Q (new_AGEMA_signal_12424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7391 ( .C (clk), .D (new_AGEMA_signal_12427), .Q (new_AGEMA_signal_12428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7395 ( .C (clk), .D (new_AGEMA_signal_12431), .Q (new_AGEMA_signal_12432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7399 ( .C (clk), .D (new_AGEMA_signal_12435), .Q (new_AGEMA_signal_12436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7403 ( .C (clk), .D (new_AGEMA_signal_12439), .Q (new_AGEMA_signal_12440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7407 ( .C (clk), .D (new_AGEMA_signal_12443), .Q (new_AGEMA_signal_12444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7411 ( .C (clk), .D (new_AGEMA_signal_12447), .Q (new_AGEMA_signal_12448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7415 ( .C (clk), .D (new_AGEMA_signal_12451), .Q (new_AGEMA_signal_12452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7419 ( .C (clk), .D (new_AGEMA_signal_12455), .Q (new_AGEMA_signal_12456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7423 ( .C (clk), .D (new_AGEMA_signal_12459), .Q (new_AGEMA_signal_12460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7427 ( .C (clk), .D (new_AGEMA_signal_12463), .Q (new_AGEMA_signal_12464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7431 ( .C (clk), .D (new_AGEMA_signal_12467), .Q (new_AGEMA_signal_12468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7435 ( .C (clk), .D (new_AGEMA_signal_12471), .Q (new_AGEMA_signal_12472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7439 ( .C (clk), .D (new_AGEMA_signal_12475), .Q (new_AGEMA_signal_12476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7443 ( .C (clk), .D (new_AGEMA_signal_12479), .Q (new_AGEMA_signal_12480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7447 ( .C (clk), .D (new_AGEMA_signal_12483), .Q (new_AGEMA_signal_12484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7451 ( .C (clk), .D (new_AGEMA_signal_12487), .Q (new_AGEMA_signal_12488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7455 ( .C (clk), .D (new_AGEMA_signal_12491), .Q (new_AGEMA_signal_12492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7459 ( .C (clk), .D (new_AGEMA_signal_12495), .Q (new_AGEMA_signal_12496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7463 ( .C (clk), .D (new_AGEMA_signal_12499), .Q (new_AGEMA_signal_12500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7467 ( .C (clk), .D (new_AGEMA_signal_12503), .Q (new_AGEMA_signal_12504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7471 ( .C (clk), .D (new_AGEMA_signal_12507), .Q (new_AGEMA_signal_12508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7475 ( .C (clk), .D (new_AGEMA_signal_12511), .Q (new_AGEMA_signal_12512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7479 ( .C (clk), .D (new_AGEMA_signal_12515), .Q (new_AGEMA_signal_12516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7483 ( .C (clk), .D (new_AGEMA_signal_12519), .Q (new_AGEMA_signal_12520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7487 ( .C (clk), .D (new_AGEMA_signal_12523), .Q (new_AGEMA_signal_12524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7491 ( .C (clk), .D (new_AGEMA_signal_12527), .Q (new_AGEMA_signal_12528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7495 ( .C (clk), .D (new_AGEMA_signal_12531), .Q (new_AGEMA_signal_12532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7499 ( .C (clk), .D (new_AGEMA_signal_12535), .Q (new_AGEMA_signal_12536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7503 ( .C (clk), .D (new_AGEMA_signal_12539), .Q (new_AGEMA_signal_12540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7507 ( .C (clk), .D (new_AGEMA_signal_12543), .Q (new_AGEMA_signal_12544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7511 ( .C (clk), .D (new_AGEMA_signal_12547), .Q (new_AGEMA_signal_12548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7515 ( .C (clk), .D (new_AGEMA_signal_12551), .Q (new_AGEMA_signal_12552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7519 ( .C (clk), .D (new_AGEMA_signal_12555), .Q (new_AGEMA_signal_12556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7523 ( .C (clk), .D (new_AGEMA_signal_12559), .Q (new_AGEMA_signal_12560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7527 ( .C (clk), .D (new_AGEMA_signal_12563), .Q (new_AGEMA_signal_12564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7531 ( .C (clk), .D (new_AGEMA_signal_12567), .Q (new_AGEMA_signal_12568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7535 ( .C (clk), .D (new_AGEMA_signal_12571), .Q (new_AGEMA_signal_12572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7539 ( .C (clk), .D (new_AGEMA_signal_12575), .Q (new_AGEMA_signal_12576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7543 ( .C (clk), .D (new_AGEMA_signal_12579), .Q (new_AGEMA_signal_12580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7547 ( .C (clk), .D (new_AGEMA_signal_12583), .Q (new_AGEMA_signal_12584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7551 ( .C (clk), .D (new_AGEMA_signal_12587), .Q (new_AGEMA_signal_12588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7555 ( .C (clk), .D (new_AGEMA_signal_12591), .Q (new_AGEMA_signal_12592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7559 ( .C (clk), .D (new_AGEMA_signal_12595), .Q (new_AGEMA_signal_12596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7563 ( .C (clk), .D (new_AGEMA_signal_12599), .Q (new_AGEMA_signal_12600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7567 ( .C (clk), .D (new_AGEMA_signal_12603), .Q (new_AGEMA_signal_12604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7571 ( .C (clk), .D (new_AGEMA_signal_12607), .Q (new_AGEMA_signal_12608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7575 ( .C (clk), .D (new_AGEMA_signal_12611), .Q (new_AGEMA_signal_12612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7579 ( .C (clk), .D (new_AGEMA_signal_12615), .Q (new_AGEMA_signal_12616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7583 ( .C (clk), .D (new_AGEMA_signal_12619), .Q (new_AGEMA_signal_12620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7587 ( .C (clk), .D (new_AGEMA_signal_12623), .Q (new_AGEMA_signal_12624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7591 ( .C (clk), .D (new_AGEMA_signal_12627), .Q (new_AGEMA_signal_12628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7595 ( .C (clk), .D (new_AGEMA_signal_12631), .Q (new_AGEMA_signal_12632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7599 ( .C (clk), .D (new_AGEMA_signal_12635), .Q (new_AGEMA_signal_12636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7603 ( .C (clk), .D (new_AGEMA_signal_12639), .Q (new_AGEMA_signal_12640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7607 ( .C (clk), .D (new_AGEMA_signal_12643), .Q (new_AGEMA_signal_12644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7611 ( .C (clk), .D (new_AGEMA_signal_12647), .Q (new_AGEMA_signal_12648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7615 ( .C (clk), .D (new_AGEMA_signal_12651), .Q (new_AGEMA_signal_12652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7619 ( .C (clk), .D (new_AGEMA_signal_12655), .Q (new_AGEMA_signal_12656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7623 ( .C (clk), .D (new_AGEMA_signal_12659), .Q (new_AGEMA_signal_12660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7627 ( .C (clk), .D (new_AGEMA_signal_12663), .Q (new_AGEMA_signal_12664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7631 ( .C (clk), .D (new_AGEMA_signal_12667), .Q (new_AGEMA_signal_12668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7635 ( .C (clk), .D (new_AGEMA_signal_12671), .Q (new_AGEMA_signal_12672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7639 ( .C (clk), .D (new_AGEMA_signal_12675), .Q (new_AGEMA_signal_12676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7643 ( .C (clk), .D (new_AGEMA_signal_12679), .Q (new_AGEMA_signal_12680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7647 ( .C (clk), .D (new_AGEMA_signal_12683), .Q (new_AGEMA_signal_12684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7651 ( .C (clk), .D (new_AGEMA_signal_12687), .Q (new_AGEMA_signal_12688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7655 ( .C (clk), .D (new_AGEMA_signal_12691), .Q (new_AGEMA_signal_12692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7659 ( .C (clk), .D (new_AGEMA_signal_12695), .Q (new_AGEMA_signal_12696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7663 ( .C (clk), .D (new_AGEMA_signal_12699), .Q (new_AGEMA_signal_12700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7667 ( .C (clk), .D (new_AGEMA_signal_12703), .Q (new_AGEMA_signal_12704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7671 ( .C (clk), .D (new_AGEMA_signal_12707), .Q (new_AGEMA_signal_12708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7675 ( .C (clk), .D (new_AGEMA_signal_12711), .Q (new_AGEMA_signal_12712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7679 ( .C (clk), .D (new_AGEMA_signal_12715), .Q (new_AGEMA_signal_12716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7683 ( .C (clk), .D (new_AGEMA_signal_12719), .Q (new_AGEMA_signal_12720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7687 ( .C (clk), .D (new_AGEMA_signal_12723), .Q (new_AGEMA_signal_12724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7691 ( .C (clk), .D (new_AGEMA_signal_12727), .Q (new_AGEMA_signal_12728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7695 ( .C (clk), .D (new_AGEMA_signal_12731), .Q (new_AGEMA_signal_12732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7699 ( .C (clk), .D (new_AGEMA_signal_12735), .Q (new_AGEMA_signal_12736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7703 ( .C (clk), .D (new_AGEMA_signal_12739), .Q (new_AGEMA_signal_12740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7707 ( .C (clk), .D (new_AGEMA_signal_12743), .Q (new_AGEMA_signal_12744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7711 ( .C (clk), .D (new_AGEMA_signal_12747), .Q (new_AGEMA_signal_12748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7715 ( .C (clk), .D (new_AGEMA_signal_12751), .Q (new_AGEMA_signal_12752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7719 ( .C (clk), .D (new_AGEMA_signal_12755), .Q (new_AGEMA_signal_12756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7723 ( .C (clk), .D (new_AGEMA_signal_12759), .Q (new_AGEMA_signal_12760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7727 ( .C (clk), .D (new_AGEMA_signal_12763), .Q (new_AGEMA_signal_12764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7731 ( .C (clk), .D (new_AGEMA_signal_12767), .Q (new_AGEMA_signal_12768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7735 ( .C (clk), .D (new_AGEMA_signal_12771), .Q (new_AGEMA_signal_12772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7739 ( .C (clk), .D (new_AGEMA_signal_12775), .Q (new_AGEMA_signal_12776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7743 ( .C (clk), .D (new_AGEMA_signal_12779), .Q (new_AGEMA_signal_12780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7747 ( .C (clk), .D (new_AGEMA_signal_12783), .Q (new_AGEMA_signal_12784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7751 ( .C (clk), .D (new_AGEMA_signal_12787), .Q (new_AGEMA_signal_12788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7755 ( .C (clk), .D (new_AGEMA_signal_12791), .Q (new_AGEMA_signal_12792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7759 ( .C (clk), .D (new_AGEMA_signal_12795), .Q (new_AGEMA_signal_12796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7763 ( .C (clk), .D (new_AGEMA_signal_12799), .Q (new_AGEMA_signal_12800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7767 ( .C (clk), .D (new_AGEMA_signal_12803), .Q (new_AGEMA_signal_12804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7771 ( .C (clk), .D (new_AGEMA_signal_12807), .Q (new_AGEMA_signal_12808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7775 ( .C (clk), .D (new_AGEMA_signal_12811), .Q (new_AGEMA_signal_12812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7779 ( .C (clk), .D (new_AGEMA_signal_12815), .Q (new_AGEMA_signal_12816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7783 ( .C (clk), .D (new_AGEMA_signal_12819), .Q (new_AGEMA_signal_12820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7787 ( .C (clk), .D (new_AGEMA_signal_12823), .Q (new_AGEMA_signal_12824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7791 ( .C (clk), .D (new_AGEMA_signal_12827), .Q (new_AGEMA_signal_12828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7795 ( .C (clk), .D (new_AGEMA_signal_12831), .Q (new_AGEMA_signal_12832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7799 ( .C (clk), .D (new_AGEMA_signal_12835), .Q (new_AGEMA_signal_12836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7803 ( .C (clk), .D (new_AGEMA_signal_12839), .Q (new_AGEMA_signal_12840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7807 ( .C (clk), .D (new_AGEMA_signal_12843), .Q (new_AGEMA_signal_12844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7811 ( .C (clk), .D (new_AGEMA_signal_12847), .Q (new_AGEMA_signal_12848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7815 ( .C (clk), .D (new_AGEMA_signal_12851), .Q (new_AGEMA_signal_12852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7819 ( .C (clk), .D (new_AGEMA_signal_12855), .Q (new_AGEMA_signal_12856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7823 ( .C (clk), .D (new_AGEMA_signal_12859), .Q (new_AGEMA_signal_12860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7827 ( .C (clk), .D (new_AGEMA_signal_12863), .Q (new_AGEMA_signal_12864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7831 ( .C (clk), .D (new_AGEMA_signal_12867), .Q (new_AGEMA_signal_12868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7835 ( .C (clk), .D (new_AGEMA_signal_12871), .Q (new_AGEMA_signal_12872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7839 ( .C (clk), .D (new_AGEMA_signal_12875), .Q (new_AGEMA_signal_12876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7843 ( .C (clk), .D (new_AGEMA_signal_12879), .Q (new_AGEMA_signal_12880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7847 ( .C (clk), .D (new_AGEMA_signal_12883), .Q (new_AGEMA_signal_12884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7851 ( .C (clk), .D (new_AGEMA_signal_12887), .Q (new_AGEMA_signal_12888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7855 ( .C (clk), .D (new_AGEMA_signal_12891), .Q (new_AGEMA_signal_12892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7859 ( .C (clk), .D (new_AGEMA_signal_12895), .Q (new_AGEMA_signal_12896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7863 ( .C (clk), .D (new_AGEMA_signal_12899), .Q (new_AGEMA_signal_12900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7867 ( .C (clk), .D (new_AGEMA_signal_12903), .Q (new_AGEMA_signal_12904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7871 ( .C (clk), .D (new_AGEMA_signal_12907), .Q (new_AGEMA_signal_12908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7875 ( .C (clk), .D (new_AGEMA_signal_12911), .Q (new_AGEMA_signal_12912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7879 ( .C (clk), .D (new_AGEMA_signal_12915), .Q (new_AGEMA_signal_12916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7883 ( .C (clk), .D (new_AGEMA_signal_12919), .Q (new_AGEMA_signal_12920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7887 ( .C (clk), .D (new_AGEMA_signal_12923), .Q (new_AGEMA_signal_12924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7891 ( .C (clk), .D (new_AGEMA_signal_12927), .Q (new_AGEMA_signal_12928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7895 ( .C (clk), .D (new_AGEMA_signal_12931), .Q (new_AGEMA_signal_12932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7899 ( .C (clk), .D (new_AGEMA_signal_12935), .Q (new_AGEMA_signal_12936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7903 ( .C (clk), .D (new_AGEMA_signal_12939), .Q (new_AGEMA_signal_12940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7907 ( .C (clk), .D (new_AGEMA_signal_12943), .Q (new_AGEMA_signal_12944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7911 ( .C (clk), .D (new_AGEMA_signal_12947), .Q (new_AGEMA_signal_12948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7915 ( .C (clk), .D (new_AGEMA_signal_12951), .Q (new_AGEMA_signal_12952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7919 ( .C (clk), .D (new_AGEMA_signal_12955), .Q (new_AGEMA_signal_12956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7923 ( .C (clk), .D (new_AGEMA_signal_12959), .Q (new_AGEMA_signal_12960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7927 ( .C (clk), .D (new_AGEMA_signal_12963), .Q (new_AGEMA_signal_12964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7931 ( .C (clk), .D (new_AGEMA_signal_12967), .Q (new_AGEMA_signal_12968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7935 ( .C (clk), .D (new_AGEMA_signal_12971), .Q (new_AGEMA_signal_12972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7939 ( .C (clk), .D (new_AGEMA_signal_12975), .Q (new_AGEMA_signal_12976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7943 ( .C (clk), .D (new_AGEMA_signal_12979), .Q (new_AGEMA_signal_12980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7947 ( .C (clk), .D (new_AGEMA_signal_12983), .Q (new_AGEMA_signal_12984) ) ;
    buf_clk new_AGEMA_reg_buffer_7951 ( .C (clk), .D (new_AGEMA_signal_12987), .Q (new_AGEMA_signal_12988) ) ;
    buf_clk new_AGEMA_reg_buffer_7955 ( .C (clk), .D (new_AGEMA_signal_12991), .Q (new_AGEMA_signal_12992) ) ;
    buf_clk new_AGEMA_reg_buffer_7959 ( .C (clk), .D (new_AGEMA_signal_12995), .Q (new_AGEMA_signal_12996) ) ;
    buf_clk new_AGEMA_reg_buffer_7963 ( .C (clk), .D (new_AGEMA_signal_12999), .Q (new_AGEMA_signal_13000) ) ;
    buf_clk new_AGEMA_reg_buffer_7967 ( .C (clk), .D (new_AGEMA_signal_13003), .Q (new_AGEMA_signal_13004) ) ;
    buf_clk new_AGEMA_reg_buffer_7971 ( .C (clk), .D (new_AGEMA_signal_13007), .Q (new_AGEMA_signal_13008) ) ;
    buf_clk new_AGEMA_reg_buffer_7975 ( .C (clk), .D (new_AGEMA_signal_13011), .Q (new_AGEMA_signal_13012) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, RoundOutput[0]}), .a ({new_AGEMA_signal_7257, new_AGEMA_signal_7253, new_AGEMA_signal_7249}), .c ({new_AGEMA_signal_5975, new_AGEMA_signal_5974, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6053, new_AGEMA_signal_6052, RoundOutput[1]}), .a ({new_AGEMA_signal_7269, new_AGEMA_signal_7265, new_AGEMA_signal_7261}), .c ({new_AGEMA_signal_6209, new_AGEMA_signal_6208, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5735, new_AGEMA_signal_5734, RoundOutput[2]}), .a ({new_AGEMA_signal_7281, new_AGEMA_signal_7277, new_AGEMA_signal_7273}), .c ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, RoundOutput[3]}), .a ({new_AGEMA_signal_7293, new_AGEMA_signal_7289, new_AGEMA_signal_7285}), .c ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, RoundOutput[4]}), .a ({new_AGEMA_signal_7305, new_AGEMA_signal_7301, new_AGEMA_signal_7297}), .c ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, RoundOutput[5]}), .a ({new_AGEMA_signal_7317, new_AGEMA_signal_7313, new_AGEMA_signal_7309}), .c ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, RoundOutput[6]}), .a ({new_AGEMA_signal_7329, new_AGEMA_signal_7325, new_AGEMA_signal_7321}), .c ({new_AGEMA_signal_5987, new_AGEMA_signal_5986, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5741, new_AGEMA_signal_5740, RoundOutput[7]}), .a ({new_AGEMA_signal_7341, new_AGEMA_signal_7337, new_AGEMA_signal_7333}), .c ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, RoundOutput[8]}), .a ({new_AGEMA_signal_7353, new_AGEMA_signal_7349, new_AGEMA_signal_7345}), .c ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6059, new_AGEMA_signal_6058, RoundOutput[9]}), .a ({new_AGEMA_signal_7365, new_AGEMA_signal_7361, new_AGEMA_signal_7357}), .c ({new_AGEMA_signal_6221, new_AGEMA_signal_6220, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, RoundOutput[10]}), .a ({new_AGEMA_signal_7377, new_AGEMA_signal_7373, new_AGEMA_signal_7369}), .c ({new_AGEMA_signal_5999, new_AGEMA_signal_5998, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, RoundOutput[11]}), .a ({new_AGEMA_signal_7389, new_AGEMA_signal_7385, new_AGEMA_signal_7381}), .c ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, RoundOutput[12]}), .a ({new_AGEMA_signal_7401, new_AGEMA_signal_7397, new_AGEMA_signal_7393}), .c ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5747, new_AGEMA_signal_5746, RoundOutput[13]}), .a ({new_AGEMA_signal_7413, new_AGEMA_signal_7409, new_AGEMA_signal_7405}), .c ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, RoundOutput[14]}), .a ({new_AGEMA_signal_7425, new_AGEMA_signal_7421, new_AGEMA_signal_7417}), .c ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, RoundOutput[15]}), .a ({new_AGEMA_signal_7437, new_AGEMA_signal_7433, new_AGEMA_signal_7429}), .c ({new_AGEMA_signal_6011, new_AGEMA_signal_6010, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5753, new_AGEMA_signal_5752, RoundOutput[16]}), .a ({new_AGEMA_signal_7449, new_AGEMA_signal_7445, new_AGEMA_signal_7441}), .c ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6065, new_AGEMA_signal_6064, RoundOutput[17]}), .a ({new_AGEMA_signal_7461, new_AGEMA_signal_7457, new_AGEMA_signal_7453}), .c ({new_AGEMA_signal_6233, new_AGEMA_signal_6232, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, RoundOutput[18]}), .a ({new_AGEMA_signal_7473, new_AGEMA_signal_7469, new_AGEMA_signal_7465}), .c ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, RoundOutput[19]}), .a ({new_AGEMA_signal_7485, new_AGEMA_signal_7481, new_AGEMA_signal_7477}), .c ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, RoundOutput[20]}), .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7493, new_AGEMA_signal_7489}), .c ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, RoundOutput[21]}), .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7505, new_AGEMA_signal_7501}), .c ({new_AGEMA_signal_6023, new_AGEMA_signal_6022, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5759, new_AGEMA_signal_5758, RoundOutput[22]}), .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7517, new_AGEMA_signal_7513}), .c ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, RoundOutput[23]}), .a ({new_AGEMA_signal_7533, new_AGEMA_signal_7529, new_AGEMA_signal_7525}), .c ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, RoundOutput[24]}), .a ({new_AGEMA_signal_7545, new_AGEMA_signal_7541, new_AGEMA_signal_7537}), .c ({new_AGEMA_signal_6035, new_AGEMA_signal_6034, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6071, new_AGEMA_signal_6070, RoundOutput[25]}), .a ({new_AGEMA_signal_7557, new_AGEMA_signal_7553, new_AGEMA_signal_7549}), .c ({new_AGEMA_signal_6245, new_AGEMA_signal_6244, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5765, new_AGEMA_signal_5764, RoundOutput[26]}), .a ({new_AGEMA_signal_7569, new_AGEMA_signal_7565, new_AGEMA_signal_7561}), .c ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, RoundOutput[27]}), .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7577, new_AGEMA_signal_7573}), .c ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, RoundOutput[28]}), .a ({new_AGEMA_signal_7593, new_AGEMA_signal_7589, new_AGEMA_signal_7585}), .c ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, RoundOutput[29]}), .a ({new_AGEMA_signal_7605, new_AGEMA_signal_7601, new_AGEMA_signal_7597}), .c ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, RoundOutput[30]}), .a ({new_AGEMA_signal_7617, new_AGEMA_signal_7613, new_AGEMA_signal_7609}), .c ({new_AGEMA_signal_6047, new_AGEMA_signal_6046, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5771, new_AGEMA_signal_5770, RoundOutput[31]}), .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7625, new_AGEMA_signal_7621}), .c ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7635, new_AGEMA_signal_7632}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7644, new_AGEMA_signal_7641}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_4291, new_AGEMA_signal_4290, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_7656, new_AGEMA_signal_7653, new_AGEMA_signal_7650}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7662, new_AGEMA_signal_7659}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_7674, new_AGEMA_signal_7671, new_AGEMA_signal_7668}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7683, new_AGEMA_signal_7680, new_AGEMA_signal_7677}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_7692, new_AGEMA_signal_7689, new_AGEMA_signal_7686}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_7701, new_AGEMA_signal_7698, new_AGEMA_signal_7695}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_7710, new_AGEMA_signal_7707, new_AGEMA_signal_7704}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7716, new_AGEMA_signal_7713}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_7728, new_AGEMA_signal_7725, new_AGEMA_signal_7722}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_7737, new_AGEMA_signal_7734, new_AGEMA_signal_7731}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7743, new_AGEMA_signal_7740}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_7755, new_AGEMA_signal_7752, new_AGEMA_signal_7749}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_7764, new_AGEMA_signal_7761, new_AGEMA_signal_7758}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7770, new_AGEMA_signal_7767}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_7782, new_AGEMA_signal_7779, new_AGEMA_signal_7776}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_7791, new_AGEMA_signal_7788, new_AGEMA_signal_7785}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_4291, new_AGEMA_signal_4290, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_4487, new_AGEMA_signal_4486, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_4643, new_AGEMA_signal_4642, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_4631, new_AGEMA_signal_4630, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_4571, new_AGEMA_signal_4570, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7797, new_AGEMA_signal_7794}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_7809, new_AGEMA_signal_7806, new_AGEMA_signal_7803}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_7818, new_AGEMA_signal_7815, new_AGEMA_signal_7812}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_7827, new_AGEMA_signal_7824, new_AGEMA_signal_7821}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_7836, new_AGEMA_signal_7833, new_AGEMA_signal_7830}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7845, new_AGEMA_signal_7842, new_AGEMA_signal_7839}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_7854, new_AGEMA_signal_7851, new_AGEMA_signal_7848}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_7863, new_AGEMA_signal_7860, new_AGEMA_signal_7857}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_7872, new_AGEMA_signal_7869, new_AGEMA_signal_7866}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_7881, new_AGEMA_signal_7878, new_AGEMA_signal_7875}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_7890, new_AGEMA_signal_7887, new_AGEMA_signal_7884}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_7899, new_AGEMA_signal_7896, new_AGEMA_signal_7893}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7905, new_AGEMA_signal_7902}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_7917, new_AGEMA_signal_7914, new_AGEMA_signal_7911}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_4327, new_AGEMA_signal_4326, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_7926, new_AGEMA_signal_7923, new_AGEMA_signal_7920}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7932, new_AGEMA_signal_7929}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_7944, new_AGEMA_signal_7941, new_AGEMA_signal_7938}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_7953, new_AGEMA_signal_7950, new_AGEMA_signal_7947}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_4327, new_AGEMA_signal_4326, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_4511, new_AGEMA_signal_4510, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_4667, new_AGEMA_signal_4666, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_4661, new_AGEMA_signal_4660, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4655, new_AGEMA_signal_4654, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_4667, new_AGEMA_signal_4666, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7959, new_AGEMA_signal_7956}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_7971, new_AGEMA_signal_7968, new_AGEMA_signal_7965}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_7980, new_AGEMA_signal_7977, new_AGEMA_signal_7974}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7986, new_AGEMA_signal_7983}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_7998, new_AGEMA_signal_7995, new_AGEMA_signal_7992}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_8007, new_AGEMA_signal_8004, new_AGEMA_signal_8001}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_8016, new_AGEMA_signal_8013, new_AGEMA_signal_8010}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_8025, new_AGEMA_signal_8022, new_AGEMA_signal_8019}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_8034, new_AGEMA_signal_8031, new_AGEMA_signal_8028}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_8043, new_AGEMA_signal_8040, new_AGEMA_signal_8037}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_8052, new_AGEMA_signal_8049, new_AGEMA_signal_8046}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_8061, new_AGEMA_signal_8058, new_AGEMA_signal_8055}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8067, new_AGEMA_signal_8064}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_8079, new_AGEMA_signal_8076, new_AGEMA_signal_8073}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_8088, new_AGEMA_signal_8085, new_AGEMA_signal_8082}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_8097, new_AGEMA_signal_8094, new_AGEMA_signal_8091}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_8106, new_AGEMA_signal_8103, new_AGEMA_signal_8100}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_8115, new_AGEMA_signal_8112, new_AGEMA_signal_8109}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_4673, new_AGEMA_signal_4672, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_4685, new_AGEMA_signal_4684, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4679, new_AGEMA_signal_4678, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_4673, new_AGEMA_signal_4672, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_4685, new_AGEMA_signal_4684, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_4607, new_AGEMA_signal_4606, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_8124, new_AGEMA_signal_8121, new_AGEMA_signal_8118}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_8133, new_AGEMA_signal_8130, new_AGEMA_signal_8127}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_4363, new_AGEMA_signal_4362, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_8142, new_AGEMA_signal_8139, new_AGEMA_signal_8136}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_8151, new_AGEMA_signal_8148, new_AGEMA_signal_8145}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_8160, new_AGEMA_signal_8157, new_AGEMA_signal_8154}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_8169, new_AGEMA_signal_8166, new_AGEMA_signal_8163}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_8178, new_AGEMA_signal_8175, new_AGEMA_signal_8172}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_8187, new_AGEMA_signal_8184, new_AGEMA_signal_8181}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_8196, new_AGEMA_signal_8193, new_AGEMA_signal_8190}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_8205, new_AGEMA_signal_8202, new_AGEMA_signal_8199}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_8214, new_AGEMA_signal_8211, new_AGEMA_signal_8208}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_8223, new_AGEMA_signal_8220, new_AGEMA_signal_8217}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_8232, new_AGEMA_signal_8229, new_AGEMA_signal_8226}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_8241, new_AGEMA_signal_8238, new_AGEMA_signal_8235}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_8250, new_AGEMA_signal_8247, new_AGEMA_signal_8244}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_8259, new_AGEMA_signal_8256, new_AGEMA_signal_8253}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_8268, new_AGEMA_signal_8265, new_AGEMA_signal_8262}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_8277, new_AGEMA_signal_8274, new_AGEMA_signal_8271}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_4363, new_AGEMA_signal_4362, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_4697, new_AGEMA_signal_4696, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_4703, new_AGEMA_signal_4702, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_4547, new_AGEMA_signal_4546, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_4709, new_AGEMA_signal_4708, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_4697, new_AGEMA_signal_4696, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_4703, new_AGEMA_signal_4702, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U96 ( .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, MixColumnsIns_n64}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_5395, new_AGEMA_signal_5394, MixColumnsOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U95 ( .a ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, MixColumnsIns_n63}), .b ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, MixColumnsIns_n62}), .c ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, MixColumnsIns_n64}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U94 ( .a ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, MixColumnsIns_n61}), .b ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, MixColumnsIns_n60}), .c ({new_AGEMA_signal_5105, new_AGEMA_signal_5104, MixColumnsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U93 ( .a ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, MixColumnsIns_n59}), .b ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, MixColumnsIns_n61}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U92 ( .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, MixColumnsIns_n58}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, MixColumnsIns_n57}), .c ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, MixColumnsOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U91 ( .a ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, MixColumnsIns_n56}), .b ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, MixColumnsIns_n58}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U90 ( .a ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, MixColumnsIns_n55}), .b ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, MixColumnsIns_n54}), .c ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, MixColumnsOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U89 ( .a ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, MixColumnsIns_n53}), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, MixColumnsIns_n55}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U88 ( .a ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, MixColumnsIns_n52}), .b ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, MixColumnsIns_n51}), .c ({new_AGEMA_signal_5111, new_AGEMA_signal_5110, MixColumnsOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U87 ( .a ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, MixColumnsIns_n50}), .b ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, MixColumnsIns_n52}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U86 ( .a ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, MixColumnsIns_n49}), .b ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, MixColumnsIns_n48}), .c ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, MixColumnsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U85 ( .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, MixColumnsIns_n47}), .b ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, MixColumnsIns_n49}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U84 ( .a ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, MixColumnsIns_n46}), .b ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, MixColumnsIns_n45}), .c ({new_AGEMA_signal_5399, new_AGEMA_signal_5398, MixColumnsOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U83 ( .a ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, MixColumnsIns_n44}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, MixColumnsIns_n46}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U82 ( .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, MixColumnsIns_n43}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, MixColumnsIns_n57}), .c ({new_AGEMA_signal_5117, new_AGEMA_signal_5116, MixColumnsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U81 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, MixColumnsIns_n57}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U80 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, MixColumnsIns_n42}), .c ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, MixColumnsIns_n43}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U79 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, MixColumnsIns_n41}), .b ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, MixColumnsIns_n54}), .c ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, MixColumnsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U78 ( .a ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, MixColumnsIns_n54}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U77 ( .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, MixColumnsIns_n40}), .c ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, MixColumnsIns_n41}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U76 ( .a ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, MixColumnsIns_n39}), .b ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, MixColumnsIns_n38}), .c ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, MixColumnsOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U75 ( .a ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, MixColumnsIns_n37}), .b ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, MixColumnsIns_n39}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U74 ( .a ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, MixColumnsIns_n36}), .b ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, MixColumnsIns_n51}), .c ({new_AGEMA_signal_5123, new_AGEMA_signal_5122, MixColumnsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U73 ( .a ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .b ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, MixColumnsIns_n51}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U72 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, MixColumnsIns_n35}), .c ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, MixColumnsIns_n36}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U71 ( .a ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, MixColumnsIns_n34}), .b ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, MixColumnsIns_n48}), .c ({new_AGEMA_signal_5401, new_AGEMA_signal_5400, MixColumnsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U70 ( .a ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .b ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, MixColumnsIns_DoubleBytes[28]}), .c ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, MixColumnsIns_n48}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U69 ( .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, MixColumnsIns_n33}), .c ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, MixColumnsIns_n34}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U68 ( .a ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, MixColumnsIns_n32}), .b ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, MixColumnsIns_n45}), .c ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, MixColumnsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U67 ( .a ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .b ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, MixColumnsIns_DoubleBytes[27]}), .c ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, MixColumnsIns_n45}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U66 ( .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .b ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, MixColumnsIns_n31}), .c ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, MixColumnsIns_n32}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U65 ( .a ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, MixColumnsIns_n30}), .b ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, MixColumnsIns_n38}), .c ({new_AGEMA_signal_5129, new_AGEMA_signal_5128, MixColumnsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U64 ( .a ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .b ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, MixColumnsIns_n38}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U63 ( .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .b ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, MixColumnsIns_n29}), .c ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, MixColumnsIns_n30}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U62 ( .a ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, MixColumnsIns_n28}), .b ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, MixColumnsIns_n27}), .c ({new_AGEMA_signal_5405, new_AGEMA_signal_5404, MixColumnsOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U61 ( .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, MixColumnsIns_n26}), .c ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, MixColumnsIns_n28}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U60 ( .a ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, MixColumnsIns_n25}), .b ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, MixColumnsIns_n24}), .c ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, MixColumnsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U59 ( .a ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, MixColumnsIns_n23}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, MixColumnsIns_n25}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U58 ( .a ({new_AGEMA_signal_4937, new_AGEMA_signal_4936, MixColumnsIns_n22}), .b ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, MixColumnsIns_n42}), .c ({new_AGEMA_signal_5135, new_AGEMA_signal_5134, MixColumnsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U57 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, MixColumnsIns_n42}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U56 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, MixColumnsIns_n21}), .c ({new_AGEMA_signal_4937, new_AGEMA_signal_4936, MixColumnsIns_n22}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U55 ( .a ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, MixColumnsIns_n20}), .b ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, MixColumnsIns_n40}), .c ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, MixColumnsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U54 ( .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .b ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, MixColumnsIns_n40}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U53 ( .a ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .b ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, MixColumnsIns_n19}), .c ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, MixColumnsIns_n20}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U52 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, MixColumnsIns_n18}), .b ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, MixColumnsIns_n35}), .c ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, MixColumnsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U51 ( .a ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, MixColumnsIns_n35}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U50 ( .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .b ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, MixColumnsIns_n17}), .c ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, MixColumnsIns_n18}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U49 ( .a ({new_AGEMA_signal_5141, new_AGEMA_signal_5140, MixColumnsIns_n16}), .b ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, MixColumnsIns_n33}), .c ({new_AGEMA_signal_5407, new_AGEMA_signal_5406, MixColumnsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U48 ( .a ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .b ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, MixColumnsIns_DoubleBytes[20]}), .c ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, MixColumnsIns_n33}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U47 ( .a ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, MixColumnsIns_n15}), .c ({new_AGEMA_signal_5141, new_AGEMA_signal_5140, MixColumnsIns_n16}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U46 ( .a ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, MixColumnsIns_n14}), .b ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, MixColumnsIns_n27}), .c ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, MixColumnsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U45 ( .a ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .b ({new_AGEMA_signal_4823, new_AGEMA_signal_4822, MixColumnsIns_DoubleBytes[25]}), .c ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, MixColumnsIns_n27}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U44 ( .a ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .b ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, MixColumnsIns_n62}), .c ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, MixColumnsIns_n14}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U43 ( .a ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .b ({new_AGEMA_signal_4841, new_AGEMA_signal_4840, MixColumnsIns_DoubleBytes[1]}), .c ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, MixColumnsIns_n62}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U42 ( .a ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, MixColumnsIns_n13}), .b ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, MixColumnsIns_n31}), .c ({new_AGEMA_signal_5411, new_AGEMA_signal_5410, MixColumnsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U41 ( .a ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .b ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, MixColumnsIns_DoubleBytes[19]}), .c ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, MixColumnsIns_n31}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U40 ( .a ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .b ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, MixColumnsIns_n12}), .c ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, MixColumnsIns_n13}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U39 ( .a ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, MixColumnsIns_n11}), .b ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, MixColumnsIns_n29}), .c ({new_AGEMA_signal_5147, new_AGEMA_signal_5146, MixColumnsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U38 ( .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, MixColumnsIns_n29}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U37 ( .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .b ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, MixColumnsIns_n10}), .c ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, MixColumnsIns_n11}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U36 ( .a ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, MixColumnsIns_n9}), .b ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, MixColumnsIns_n26}), .c ({new_AGEMA_signal_5413, new_AGEMA_signal_5412, MixColumnsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U35 ( .a ({new_AGEMA_signal_4829, new_AGEMA_signal_4828, MixColumnsIns_DoubleBytes[17]}), .b ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, MixColumnsIns_n26}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U34 ( .a ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, MixColumnsIns_n63}), .b ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, MixColumnsIns_n9}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U33 ( .a ({new_AGEMA_signal_4835, new_AGEMA_signal_4834, MixColumnsIns_DoubleBytes[9]}), .b ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, MixColumnsIns_n63}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U32 ( .a ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, MixColumnsIns_n8}), .b ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, MixColumnsIns_n24}), .c ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, MixColumnsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U31 ( .a ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, MixColumnsIns_n24}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U30 ( .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .b ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, MixColumnsIns_n60}), .c ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, MixColumnsIns_n8}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U29 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, MixColumnsIns_n60}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U28 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, MixColumnsIns_n7}), .b ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, MixColumnsIns_n21}), .c ({new_AGEMA_signal_5153, new_AGEMA_signal_5152, MixColumnsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U27 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, MixColumnsIns_n21}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U26 ( .a ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, MixColumnsIns_n56}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, MixColumnsIns_n7}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U25 ( .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, MixColumnsIns_n56}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U24 ( .a ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, MixColumnsIns_n6}), .b ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, MixColumnsIns_n19}), .c ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, MixColumnsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U23 ( .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, MixColumnsIns_n19}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U22 ( .a ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, MixColumnsIns_n53}), .b ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, MixColumnsIns_n6}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U21 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, MixColumnsIns_n53}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U20 ( .a ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, MixColumnsIns_n5}), .b ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, MixColumnsIns_n17}), .c ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, MixColumnsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U19 ( .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, MixColumnsIns_n17}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U18 ( .a ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, MixColumnsIns_n50}), .b ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, MixColumnsIns_n5}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U17 ( .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, MixColumnsIns_n50}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U16 ( .a ({new_AGEMA_signal_5159, new_AGEMA_signal_5158, MixColumnsIns_n4}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, MixColumnsIns_n15}), .c ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, MixColumnsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U15 ( .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, MixColumnsIns_DoubleBytes[12]}), .c ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, MixColumnsIns_n15}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U14 ( .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, MixColumnsIns_n47}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_5159, new_AGEMA_signal_5158, MixColumnsIns_n4}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U13 ( .a ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, MixColumnsIns_DoubleBytes[4]}), .b ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, MixColumnsIns_n47}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U12 ( .a ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, MixColumnsIns_n3}), .b ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, MixColumnsIns_n12}), .c ({new_AGEMA_signal_5417, new_AGEMA_signal_5416, MixColumnsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U11 ( .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .b ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, MixColumnsIns_DoubleBytes[11]}), .c ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, MixColumnsIns_n12}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U10 ( .a ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, MixColumnsIns_n44}), .b ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, MixColumnsIns_n3}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U9 ( .a ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, MixColumnsIns_DoubleBytes[3]}), .b ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, MixColumnsIns_n44}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U8 ( .a ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, MixColumnsIns_n2}), .b ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, MixColumnsIns_n10}), .c ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, MixColumnsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U7 ( .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .b ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, MixColumnsIns_n10}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U6 ( .a ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, MixColumnsIns_n37}), .b ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, MixColumnsIns_n2}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U5 ( .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, MixColumnsIns_n37}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U4 ( .a ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, MixColumnsIns_n1}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_5165, new_AGEMA_signal_5164, MixColumnsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U3 ( .a ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, MixColumnsIns_n59}), .b ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, MixColumnsIns_n23}), .c ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, MixColumnsIns_n1}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U2 ( .a ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .b ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, MixColumnsIns_n23}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_U1 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, MixColumnsIns_n59}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, MixColumnsIns_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, MixColumnsIns_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_4823, new_AGEMA_signal_4822, MixColumnsIns_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, MixColumnsIns_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, MixColumnsIns_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_4829, new_AGEMA_signal_4828, MixColumnsIns_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, MixColumnsIns_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, MixColumnsIns_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_4835, new_AGEMA_signal_4834, MixColumnsIns_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .c ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, MixColumnsIns_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .c ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, MixColumnsIns_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4841, new_AGEMA_signal_4840, MixColumnsIns_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_0_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5165, new_AGEMA_signal_5164, MixColumnsOutput[0]}), .a ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_5419, new_AGEMA_signal_5418, ColumnOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_1_U1 ( .s (new_AGEMA_signal_8285), .b ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, MixColumnsOutput[1]}), .a ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, ColumnOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_2_U1 ( .s (new_AGEMA_signal_8285), .b ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, MixColumnsOutput[2]}), .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .c ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, ColumnOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_3_U1 ( .s (new_AGEMA_signal_8285), .b ({new_AGEMA_signal_5399, new_AGEMA_signal_5398, MixColumnsOutput[3]}), .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .c ({new_AGEMA_signal_5711, new_AGEMA_signal_5710, ColumnOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_4_U1 ( .s (new_AGEMA_signal_8285), .b ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, MixColumnsOutput[4]}), .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, ColumnOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_5_U1 ( .s (new_AGEMA_signal_8285), .b ({new_AGEMA_signal_5111, new_AGEMA_signal_5110, MixColumnsOutput[5]}), .a ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_5423, new_AGEMA_signal_5422, ColumnOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_6_U1 ( .s (new_AGEMA_signal_8285), .b ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, MixColumnsOutput[6]}), .a ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_5425, new_AGEMA_signal_5424, ColumnOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_7_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, MixColumnsOutput[7]}), .a ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, ColumnOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_8_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5105, new_AGEMA_signal_5104, MixColumnsOutput[8]}), .a ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_5429, new_AGEMA_signal_5428, ColumnOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_9_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5395, new_AGEMA_signal_5394, MixColumnsOutput[9]}), .a ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, ColumnOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_10_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, MixColumnsOutput[10]}), .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_5431, new_AGEMA_signal_5430, ColumnOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_11_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5417, new_AGEMA_signal_5416, MixColumnsOutput[11]}), .a ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_5717, new_AGEMA_signal_5716, ColumnOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_12_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, MixColumnsOutput[12]}), .a ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, ColumnOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_13_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, MixColumnsOutput[13]}), .a ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, ColumnOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_14_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, MixColumnsOutput[14]}), .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_5435, new_AGEMA_signal_5434, ColumnOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_15_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5153, new_AGEMA_signal_5152, MixColumnsOutput[15]}), .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_5437, new_AGEMA_signal_5436, ColumnOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_16_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, MixColumnsOutput[16]}), .a ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, ColumnOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_17_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5413, new_AGEMA_signal_5412, MixColumnsOutput[17]}), .a ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, ColumnOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_18_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5147, new_AGEMA_signal_5146, MixColumnsOutput[18]}), .a ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_5441, new_AGEMA_signal_5440, ColumnOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_19_U1 ( .s (new_AGEMA_signal_8281), .b ({new_AGEMA_signal_5411, new_AGEMA_signal_5410, MixColumnsOutput[19]}), .a ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_5723, new_AGEMA_signal_5722, ColumnOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_20_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5407, new_AGEMA_signal_5406, MixColumnsOutput[20]}), .a ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, ColumnOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_21_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, MixColumnsOutput[21]}), .a ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_5443, new_AGEMA_signal_5442, ColumnOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_22_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, MixColumnsOutput[22]}), .a ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, ColumnOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_23_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5135, new_AGEMA_signal_5134, MixColumnsOutput[23]}), .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_5447, new_AGEMA_signal_5446, ColumnOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_24_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, MixColumnsOutput[24]}), .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_5449, new_AGEMA_signal_5448, ColumnOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_25_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5405, new_AGEMA_signal_5404, MixColumnsOutput[25]}), .a ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, ColumnOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_26_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5129, new_AGEMA_signal_5128, MixColumnsOutput[26]}), .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, ColumnOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_27_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5403, new_AGEMA_signal_5402, MixColumnsOutput[27]}), .a ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_5729, new_AGEMA_signal_5728, ColumnOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_28_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5401, new_AGEMA_signal_5400, MixColumnsOutput[28]}), .a ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, ColumnOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_29_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5123, new_AGEMA_signal_5122, MixColumnsOutput[29]}), .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_5453, new_AGEMA_signal_5452, ColumnOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_30_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, MixColumnsOutput[30]}), .a ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_5455, new_AGEMA_signal_5454, ColumnOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxMCOut_mux_inst_31_U1 ( .s (new_AGEMA_signal_8289), .b ({new_AGEMA_signal_5117, new_AGEMA_signal_5116, MixColumnsOutput[31]}), .a ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, ColumnOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_0_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5419, new_AGEMA_signal_5418, ColumnOutput[0]}), .a ({new_AGEMA_signal_8305, new_AGEMA_signal_8301, new_AGEMA_signal_8297}), .c ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_1_U1 ( .s (new_AGEMA_signal_8309), .b ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, ColumnOutput[1]}), .a ({new_AGEMA_signal_8321, new_AGEMA_signal_8317, new_AGEMA_signal_8313}), .c ({new_AGEMA_signal_6053, new_AGEMA_signal_6052, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_2_U1 ( .s (new_AGEMA_signal_8325), .b ({new_AGEMA_signal_5421, new_AGEMA_signal_5420, ColumnOutput[2]}), .a ({new_AGEMA_signal_8337, new_AGEMA_signal_8333, new_AGEMA_signal_8329}), .c ({new_AGEMA_signal_5735, new_AGEMA_signal_5734, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_3_U1 ( .s (new_AGEMA_signal_8341), .b ({new_AGEMA_signal_5711, new_AGEMA_signal_5710, ColumnOutput[3]}), .a ({new_AGEMA_signal_8353, new_AGEMA_signal_8349, new_AGEMA_signal_8345}), .c ({new_AGEMA_signal_6055, new_AGEMA_signal_6054, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_4_U1 ( .s (new_AGEMA_signal_8357), .b ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, ColumnOutput[4]}), .a ({new_AGEMA_signal_8369, new_AGEMA_signal_8365, new_AGEMA_signal_8361}), .c ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_5_U1 ( .s (new_AGEMA_signal_8373), .b ({new_AGEMA_signal_5423, new_AGEMA_signal_5422, ColumnOutput[5]}), .a ({new_AGEMA_signal_8385, new_AGEMA_signal_8381, new_AGEMA_signal_8377}), .c ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_6_U1 ( .s (new_AGEMA_signal_8389), .b ({new_AGEMA_signal_5425, new_AGEMA_signal_5424, ColumnOutput[6]}), .a ({new_AGEMA_signal_8401, new_AGEMA_signal_8397, new_AGEMA_signal_8393}), .c ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_7_U1 ( .s (new_AGEMA_signal_8309), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, ColumnOutput[7]}), .a ({new_AGEMA_signal_8413, new_AGEMA_signal_8409, new_AGEMA_signal_8405}), .c ({new_AGEMA_signal_5741, new_AGEMA_signal_5740, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_8_U1 ( .s (new_AGEMA_signal_8357), .b ({new_AGEMA_signal_5429, new_AGEMA_signal_5428, ColumnOutput[8]}), .a ({new_AGEMA_signal_8425, new_AGEMA_signal_8421, new_AGEMA_signal_8417}), .c ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_9_U1 ( .s (new_AGEMA_signal_8309), .b ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, ColumnOutput[9]}), .a ({new_AGEMA_signal_8437, new_AGEMA_signal_8433, new_AGEMA_signal_8429}), .c ({new_AGEMA_signal_6059, new_AGEMA_signal_6058, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_10_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5431, new_AGEMA_signal_5430, ColumnOutput[10]}), .a ({new_AGEMA_signal_8449, new_AGEMA_signal_8445, new_AGEMA_signal_8441}), .c ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_11_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5717, new_AGEMA_signal_5716, ColumnOutput[11]}), .a ({new_AGEMA_signal_8461, new_AGEMA_signal_8457, new_AGEMA_signal_8453}), .c ({new_AGEMA_signal_6061, new_AGEMA_signal_6060, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_12_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, ColumnOutput[12]}), .a ({new_AGEMA_signal_8473, new_AGEMA_signal_8469, new_AGEMA_signal_8465}), .c ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_13_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, ColumnOutput[13]}), .a ({new_AGEMA_signal_8485, new_AGEMA_signal_8481, new_AGEMA_signal_8477}), .c ({new_AGEMA_signal_5747, new_AGEMA_signal_5746, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_14_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5435, new_AGEMA_signal_5434, ColumnOutput[14]}), .a ({new_AGEMA_signal_8497, new_AGEMA_signal_8493, new_AGEMA_signal_8489}), .c ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_15_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5437, new_AGEMA_signal_5436, ColumnOutput[15]}), .a ({new_AGEMA_signal_8509, new_AGEMA_signal_8505, new_AGEMA_signal_8501}), .c ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_16_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5439, new_AGEMA_signal_5438, ColumnOutput[16]}), .a ({new_AGEMA_signal_8521, new_AGEMA_signal_8517, new_AGEMA_signal_8513}), .c ({new_AGEMA_signal_5753, new_AGEMA_signal_5752, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_17_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, ColumnOutput[17]}), .a ({new_AGEMA_signal_8533, new_AGEMA_signal_8529, new_AGEMA_signal_8525}), .c ({new_AGEMA_signal_6065, new_AGEMA_signal_6064, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_18_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5441, new_AGEMA_signal_5440, ColumnOutput[18]}), .a ({new_AGEMA_signal_8545, new_AGEMA_signal_8541, new_AGEMA_signal_8537}), .c ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_19_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5723, new_AGEMA_signal_5722, ColumnOutput[19]}), .a ({new_AGEMA_signal_8557, new_AGEMA_signal_8553, new_AGEMA_signal_8549}), .c ({new_AGEMA_signal_6067, new_AGEMA_signal_6066, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_20_U1 ( .s (new_AGEMA_signal_8325), .b ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, ColumnOutput[20]}), .a ({new_AGEMA_signal_8569, new_AGEMA_signal_8565, new_AGEMA_signal_8561}), .c ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_21_U1 ( .s (new_AGEMA_signal_8341), .b ({new_AGEMA_signal_5443, new_AGEMA_signal_5442, ColumnOutput[21]}), .a ({new_AGEMA_signal_8581, new_AGEMA_signal_8577, new_AGEMA_signal_8573}), .c ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_22_U1 ( .s (new_AGEMA_signal_8357), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, ColumnOutput[22]}), .a ({new_AGEMA_signal_8593, new_AGEMA_signal_8589, new_AGEMA_signal_8585}), .c ({new_AGEMA_signal_5759, new_AGEMA_signal_5758, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_23_U1 ( .s (new_AGEMA_signal_8373), .b ({new_AGEMA_signal_5447, new_AGEMA_signal_5446, ColumnOutput[23]}), .a ({new_AGEMA_signal_8605, new_AGEMA_signal_8601, new_AGEMA_signal_8597}), .c ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_24_U1 ( .s (new_AGEMA_signal_8389), .b ({new_AGEMA_signal_5449, new_AGEMA_signal_5448, ColumnOutput[24]}), .a ({new_AGEMA_signal_8617, new_AGEMA_signal_8613, new_AGEMA_signal_8609}), .c ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_25_U1 ( .s (new_AGEMA_signal_8357), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, ColumnOutput[25]}), .a ({new_AGEMA_signal_8629, new_AGEMA_signal_8625, new_AGEMA_signal_8621}), .c ({new_AGEMA_signal_6071, new_AGEMA_signal_6070, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_26_U1 ( .s (new_AGEMA_signal_8373), .b ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, ColumnOutput[26]}), .a ({new_AGEMA_signal_8641, new_AGEMA_signal_8637, new_AGEMA_signal_8633}), .c ({new_AGEMA_signal_5765, new_AGEMA_signal_5764, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_27_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5729, new_AGEMA_signal_5728, ColumnOutput[27]}), .a ({new_AGEMA_signal_8653, new_AGEMA_signal_8649, new_AGEMA_signal_8645}), .c ({new_AGEMA_signal_6073, new_AGEMA_signal_6072, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_28_U1 ( .s (new_AGEMA_signal_8293), .b ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, ColumnOutput[28]}), .a ({new_AGEMA_signal_8665, new_AGEMA_signal_8661, new_AGEMA_signal_8657}), .c ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_29_U1 ( .s (new_AGEMA_signal_8309), .b ({new_AGEMA_signal_5453, new_AGEMA_signal_5452, ColumnOutput[29]}), .a ({new_AGEMA_signal_8677, new_AGEMA_signal_8673, new_AGEMA_signal_8669}), .c ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_30_U1 ( .s (new_AGEMA_signal_8325), .b ({new_AGEMA_signal_5455, new_AGEMA_signal_5454, ColumnOutput[30]}), .a ({new_AGEMA_signal_8689, new_AGEMA_signal_8685, new_AGEMA_signal_8681}), .c ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxRound_mux_inst_31_U1 ( .s (new_AGEMA_signal_8341), .b ({new_AGEMA_signal_5457, new_AGEMA_signal_5456, ColumnOutput[31]}), .a ({new_AGEMA_signal_8701, new_AGEMA_signal_8697, new_AGEMA_signal_8693}), .c ({new_AGEMA_signal_5771, new_AGEMA_signal_5770, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5645, new_AGEMA_signal_5644, RoundKeyOutput[0]}), .a ({new_AGEMA_signal_8713, new_AGEMA_signal_8709, new_AGEMA_signal_8705}), .c ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5915, new_AGEMA_signal_5914, RoundKeyOutput[1]}), .a ({new_AGEMA_signal_8725, new_AGEMA_signal_8721, new_AGEMA_signal_8717}), .c ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, RoundKeyOutput[2]}), .a ({new_AGEMA_signal_8737, new_AGEMA_signal_8733, new_AGEMA_signal_8729}), .c ({new_AGEMA_signal_6083, new_AGEMA_signal_6082, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, RoundKeyOutput[3]}), .a ({new_AGEMA_signal_8749, new_AGEMA_signal_8745, new_AGEMA_signal_8741}), .c ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5921, new_AGEMA_signal_5920, RoundKeyOutput[4]}), .a ({new_AGEMA_signal_8761, new_AGEMA_signal_8757, new_AGEMA_signal_8753}), .c ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, RoundKeyOutput[5]}), .a ({new_AGEMA_signal_8773, new_AGEMA_signal_8769, new_AGEMA_signal_8765}), .c ({new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, RoundKeyOutput[6]}), .a ({new_AGEMA_signal_8785, new_AGEMA_signal_8781, new_AGEMA_signal_8777}), .c ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5927, new_AGEMA_signal_5926, RoundKeyOutput[7]}), .a ({new_AGEMA_signal_8797, new_AGEMA_signal_8793, new_AGEMA_signal_8789}), .c ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, RoundKeyOutput[8]}), .a ({new_AGEMA_signal_8809, new_AGEMA_signal_8805, new_AGEMA_signal_8801}), .c ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, RoundKeyOutput[9]}), .a ({new_AGEMA_signal_8821, new_AGEMA_signal_8817, new_AGEMA_signal_8813}), .c ({new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, RoundKeyOutput[10]}), .a ({new_AGEMA_signal_8833, new_AGEMA_signal_8829, new_AGEMA_signal_8825}), .c ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5933, new_AGEMA_signal_5932, RoundKeyOutput[11]}), .a ({new_AGEMA_signal_8845, new_AGEMA_signal_8841, new_AGEMA_signal_8837}), .c ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, RoundKeyOutput[12]}), .a ({new_AGEMA_signal_8857, new_AGEMA_signal_8853, new_AGEMA_signal_8849}), .c ({new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, RoundKeyOutput[13]}), .a ({new_AGEMA_signal_8869, new_AGEMA_signal_8865, new_AGEMA_signal_8861}), .c ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5939, new_AGEMA_signal_5938, RoundKeyOutput[14]}), .a ({new_AGEMA_signal_8881, new_AGEMA_signal_8877, new_AGEMA_signal_8873}), .c ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, RoundKeyOutput[15]}), .a ({new_AGEMA_signal_8893, new_AGEMA_signal_8889, new_AGEMA_signal_8885}), .c ({new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, RoundKeyOutput[16]}), .a ({new_AGEMA_signal_8905, new_AGEMA_signal_8901, new_AGEMA_signal_8897}), .c ({new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, RoundKeyOutput[17]}), .a ({new_AGEMA_signal_8917, new_AGEMA_signal_8913, new_AGEMA_signal_8909}), .c ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5945, new_AGEMA_signal_5944, RoundKeyOutput[18]}), .a ({new_AGEMA_signal_8929, new_AGEMA_signal_8925, new_AGEMA_signal_8921}), .c ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, RoundKeyOutput[19]}), .a ({new_AGEMA_signal_8941, new_AGEMA_signal_8937, new_AGEMA_signal_8933}), .c ({new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, RoundKeyOutput[20]}), .a ({new_AGEMA_signal_8953, new_AGEMA_signal_8949, new_AGEMA_signal_8945}), .c ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5951, new_AGEMA_signal_5950, RoundKeyOutput[21]}), .a ({new_AGEMA_signal_8965, new_AGEMA_signal_8961, new_AGEMA_signal_8957}), .c ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, RoundKeyOutput[22]}), .a ({new_AGEMA_signal_8977, new_AGEMA_signal_8973, new_AGEMA_signal_8969}), .c ({new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, RoundKeyOutput[23]}), .a ({new_AGEMA_signal_8989, new_AGEMA_signal_8985, new_AGEMA_signal_8981}), .c ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5957, new_AGEMA_signal_5956, RoundKeyOutput[24]}), .a ({new_AGEMA_signal_9001, new_AGEMA_signal_8997, new_AGEMA_signal_8993}), .c ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, RoundKeyOutput[25]}), .a ({new_AGEMA_signal_9013, new_AGEMA_signal_9009, new_AGEMA_signal_9005}), .c ({new_AGEMA_signal_6257, new_AGEMA_signal_6256, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, RoundKeyOutput[26]}), .a ({new_AGEMA_signal_9025, new_AGEMA_signal_9021, new_AGEMA_signal_9017}), .c ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6197, new_AGEMA_signal_6196, RoundKeyOutput[27]}), .a ({new_AGEMA_signal_9037, new_AGEMA_signal_9033, new_AGEMA_signal_9029}), .c ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, RoundKeyOutput[28]}), .a ({new_AGEMA_signal_9049, new_AGEMA_signal_9045, new_AGEMA_signal_9041}), .c ({new_AGEMA_signal_6269, new_AGEMA_signal_6268, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, RoundKeyOutput[29]}), .a ({new_AGEMA_signal_9061, new_AGEMA_signal_9057, new_AGEMA_signal_9053}), .c ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6203, new_AGEMA_signal_6202, RoundKeyOutput[30]}), .a ({new_AGEMA_signal_9073, new_AGEMA_signal_9069, new_AGEMA_signal_9065}), .c ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, RoundKeyOutput[31]}), .a ({new_AGEMA_signal_9085, new_AGEMA_signal_9081, new_AGEMA_signal_9077}), .c ({new_AGEMA_signal_6281, new_AGEMA_signal_6280, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, RoundKeyOutput[32]}), .a ({new_AGEMA_signal_9097, new_AGEMA_signal_9093, new_AGEMA_signal_9089}), .c ({new_AGEMA_signal_5461, new_AGEMA_signal_5460, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKeyOutput[33]}), .a ({new_AGEMA_signal_9109, new_AGEMA_signal_9105, new_AGEMA_signal_9101}), .c ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, RoundKeyOutput[34]}), .a ({new_AGEMA_signal_9121, new_AGEMA_signal_9117, new_AGEMA_signal_9113}), .c ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5655, new_AGEMA_signal_5654, RoundKeyOutput[35]}), .a ({new_AGEMA_signal_9133, new_AGEMA_signal_9129, new_AGEMA_signal_9125}), .c ({new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundKeyOutput[36]}), .a ({new_AGEMA_signal_9145, new_AGEMA_signal_9141, new_AGEMA_signal_9137}), .c ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, RoundKeyOutput[37]}), .a ({new_AGEMA_signal_9157, new_AGEMA_signal_9153, new_AGEMA_signal_9149}), .c ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, RoundKeyOutput[38]}), .a ({new_AGEMA_signal_9169, new_AGEMA_signal_9165, new_AGEMA_signal_9161}), .c ({new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5663, new_AGEMA_signal_5662, RoundKeyOutput[39]}), .a ({new_AGEMA_signal_9181, new_AGEMA_signal_9177, new_AGEMA_signal_9173}), .c ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundKeyOutput[40]}), .a ({new_AGEMA_signal_9193, new_AGEMA_signal_9189, new_AGEMA_signal_9185}), .c ({new_AGEMA_signal_5465, new_AGEMA_signal_5464, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, RoundKeyOutput[41]}), .a ({new_AGEMA_signal_9205, new_AGEMA_signal_9201, new_AGEMA_signal_9197}), .c ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, RoundKeyOutput[42]}), .a ({new_AGEMA_signal_9217, new_AGEMA_signal_9213, new_AGEMA_signal_9209}), .c ({new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKeyOutput[43]}), .a ({new_AGEMA_signal_9229, new_AGEMA_signal_9225, new_AGEMA_signal_9221}), .c ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, RoundKeyOutput[44]}), .a ({new_AGEMA_signal_9241, new_AGEMA_signal_9237, new_AGEMA_signal_9233}), .c ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, RoundKeyOutput[45]}), .a ({new_AGEMA_signal_9253, new_AGEMA_signal_9249, new_AGEMA_signal_9245}), .c ({new_AGEMA_signal_5831, new_AGEMA_signal_5830, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundKeyOutput[46]}), .a ({new_AGEMA_signal_9265, new_AGEMA_signal_9261, new_AGEMA_signal_9257}), .c ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, RoundKeyOutput[47]}), .a ({new_AGEMA_signal_9277, new_AGEMA_signal_9273, new_AGEMA_signal_9269}), .c ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5335, new_AGEMA_signal_5334, RoundKeyOutput[48]}), .a ({new_AGEMA_signal_9289, new_AGEMA_signal_9285, new_AGEMA_signal_9281}), .c ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, RoundKeyOutput[49]}), .a ({new_AGEMA_signal_9301, new_AGEMA_signal_9297, new_AGEMA_signal_9293}), .c ({new_AGEMA_signal_5843, new_AGEMA_signal_5842, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5681, new_AGEMA_signal_5680, RoundKeyOutput[50]}), .a ({new_AGEMA_signal_9313, new_AGEMA_signal_9309, new_AGEMA_signal_9305}), .c ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, RoundKeyOutput[51]}), .a ({new_AGEMA_signal_9325, new_AGEMA_signal_9321, new_AGEMA_signal_9317}), .c ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, RoundKeyOutput[52]}), .a ({new_AGEMA_signal_9337, new_AGEMA_signal_9333, new_AGEMA_signal_9329}), .c ({new_AGEMA_signal_5855, new_AGEMA_signal_5854, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKeyOutput[53]}), .a ({new_AGEMA_signal_9349, new_AGEMA_signal_9345, new_AGEMA_signal_9341}), .c ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, RoundKeyOutput[54]}), .a ({new_AGEMA_signal_9361, new_AGEMA_signal_9357, new_AGEMA_signal_9353}), .c ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, RoundKeyOutput[55]}), .a ({new_AGEMA_signal_9373, new_AGEMA_signal_9369, new_AGEMA_signal_9365}), .c ({new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundKeyOutput[56]}), .a ({new_AGEMA_signal_9385, new_AGEMA_signal_9381, new_AGEMA_signal_9377}), .c ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, RoundKeyOutput[57]}), .a ({new_AGEMA_signal_9397, new_AGEMA_signal_9393, new_AGEMA_signal_9389}), .c ({new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, RoundKeyOutput[58]}), .a ({new_AGEMA_signal_9409, new_AGEMA_signal_9405, new_AGEMA_signal_9401}), .c ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5963, new_AGEMA_signal_5962, RoundKeyOutput[59]}), .a ({new_AGEMA_signal_9421, new_AGEMA_signal_9417, new_AGEMA_signal_9413}), .c ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, RoundKeyOutput[60]}), .a ({new_AGEMA_signal_9433, new_AGEMA_signal_9429, new_AGEMA_signal_9425}), .c ({new_AGEMA_signal_6179, new_AGEMA_signal_6178, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, RoundKeyOutput[61]}), .a ({new_AGEMA_signal_9445, new_AGEMA_signal_9441, new_AGEMA_signal_9437}), .c ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5969, new_AGEMA_signal_5968, RoundKeyOutput[62]}), .a ({new_AGEMA_signal_9457, new_AGEMA_signal_9453, new_AGEMA_signal_9449}), .c ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, RoundKeyOutput[63]}), .a ({new_AGEMA_signal_9469, new_AGEMA_signal_9465, new_AGEMA_signal_9461}), .c ({new_AGEMA_signal_6191, new_AGEMA_signal_6190, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, RoundKeyOutput[64]}), .a ({new_AGEMA_signal_9481, new_AGEMA_signal_9477, new_AGEMA_signal_9473}), .c ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, RoundKeyOutput[65]}), .a ({new_AGEMA_signal_9493, new_AGEMA_signal_9489, new_AGEMA_signal_9485}), .c ({new_AGEMA_signal_5473, new_AGEMA_signal_5472, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5339, new_AGEMA_signal_5338, RoundKeyOutput[66]}), .a ({new_AGEMA_signal_9505, new_AGEMA_signal_9501, new_AGEMA_signal_9497}), .c ({new_AGEMA_signal_5477, new_AGEMA_signal_5476, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5341, new_AGEMA_signal_5340, RoundKeyOutput[67]}), .a ({new_AGEMA_signal_9517, new_AGEMA_signal_9513, new_AGEMA_signal_9509}), .c ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, RoundKeyOutput[68]}), .a ({new_AGEMA_signal_9529, new_AGEMA_signal_9525, new_AGEMA_signal_9521}), .c ({new_AGEMA_signal_5485, new_AGEMA_signal_5484, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKeyOutput[69]}), .a ({new_AGEMA_signal_9541, new_AGEMA_signal_9537, new_AGEMA_signal_9533}), .c ({new_AGEMA_signal_5489, new_AGEMA_signal_5488, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5347, new_AGEMA_signal_5346, RoundKeyOutput[70]}), .a ({new_AGEMA_signal_9553, new_AGEMA_signal_9549, new_AGEMA_signal_9545}), .c ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, RoundKeyOutput[71]}), .a ({new_AGEMA_signal_9565, new_AGEMA_signal_9561, new_AGEMA_signal_9557}), .c ({new_AGEMA_signal_5497, new_AGEMA_signal_5496, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, RoundKeyOutput[72]}), .a ({new_AGEMA_signal_9577, new_AGEMA_signal_9573, new_AGEMA_signal_9569}), .c ({new_AGEMA_signal_5173, new_AGEMA_signal_5172, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundKeyOutput[73]}), .a ({new_AGEMA_signal_9589, new_AGEMA_signal_9585, new_AGEMA_signal_9581}), .c ({new_AGEMA_signal_5501, new_AGEMA_signal_5500, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5353, new_AGEMA_signal_5352, RoundKeyOutput[74]}), .a ({new_AGEMA_signal_9601, new_AGEMA_signal_9597, new_AGEMA_signal_9593}), .c ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, RoundKeyOutput[75]}), .a ({new_AGEMA_signal_9613, new_AGEMA_signal_9609, new_AGEMA_signal_9605}), .c ({new_AGEMA_signal_5509, new_AGEMA_signal_5508, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5357, new_AGEMA_signal_5356, RoundKeyOutput[76]}), .a ({new_AGEMA_signal_9625, new_AGEMA_signal_9621, new_AGEMA_signal_9617}), .c ({new_AGEMA_signal_5513, new_AGEMA_signal_5512, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5359, new_AGEMA_signal_5358, RoundKeyOutput[77]}), .a ({new_AGEMA_signal_9637, new_AGEMA_signal_9633, new_AGEMA_signal_9629}), .c ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, RoundKeyOutput[78]}), .a ({new_AGEMA_signal_9649, new_AGEMA_signal_9645, new_AGEMA_signal_9641}), .c ({new_AGEMA_signal_5521, new_AGEMA_signal_5520, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKeyOutput[79]}), .a ({new_AGEMA_signal_9661, new_AGEMA_signal_9657, new_AGEMA_signal_9653}), .c ({new_AGEMA_signal_5525, new_AGEMA_signal_5524, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKeyOutput[80]}), .a ({new_AGEMA_signal_9673, new_AGEMA_signal_9669, new_AGEMA_signal_9665}), .c ({new_AGEMA_signal_5177, new_AGEMA_signal_5176, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5365, new_AGEMA_signal_5364, RoundKeyOutput[81]}), .a ({new_AGEMA_signal_9685, new_AGEMA_signal_9681, new_AGEMA_signal_9677}), .c ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, RoundKeyOutput[82]}), .a ({new_AGEMA_signal_9697, new_AGEMA_signal_9693, new_AGEMA_signal_9689}), .c ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundKeyOutput[83]}), .a ({new_AGEMA_signal_9709, new_AGEMA_signal_9705, new_AGEMA_signal_9701}), .c ({new_AGEMA_signal_5537, new_AGEMA_signal_5536, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5371, new_AGEMA_signal_5370, RoundKeyOutput[84]}), .a ({new_AGEMA_signal_9721, new_AGEMA_signal_9717, new_AGEMA_signal_9713}), .c ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, RoundKeyOutput[85]}), .a ({new_AGEMA_signal_9733, new_AGEMA_signal_9729, new_AGEMA_signal_9725}), .c ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5375, new_AGEMA_signal_5374, RoundKeyOutput[86]}), .a ({new_AGEMA_signal_9745, new_AGEMA_signal_9741, new_AGEMA_signal_9737}), .c ({new_AGEMA_signal_5549, new_AGEMA_signal_5548, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5377, new_AGEMA_signal_5376, RoundKeyOutput[87]}), .a ({new_AGEMA_signal_9757, new_AGEMA_signal_9753, new_AGEMA_signal_9749}), .c ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, RoundKeyOutput[88]}), .a ({new_AGEMA_signal_9769, new_AGEMA_signal_9765, new_AGEMA_signal_9761}), .c ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, RoundKeyOutput[89]}), .a ({new_AGEMA_signal_9781, new_AGEMA_signal_9777, new_AGEMA_signal_9773}), .c ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, RoundKeyOutput[90]}), .a ({new_AGEMA_signal_9793, new_AGEMA_signal_9789, new_AGEMA_signal_9785}), .c ({new_AGEMA_signal_5879, new_AGEMA_signal_5878, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5699, new_AGEMA_signal_5698, RoundKeyOutput[91]}), .a ({new_AGEMA_signal_9805, new_AGEMA_signal_9801, new_AGEMA_signal_9797}), .c ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, RoundKeyOutput[92]}), .a ({new_AGEMA_signal_9817, new_AGEMA_signal_9813, new_AGEMA_signal_9809}), .c ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, RoundKeyOutput[93]}), .a ({new_AGEMA_signal_9829, new_AGEMA_signal_9825, new_AGEMA_signal_9821}), .c ({new_AGEMA_signal_5891, new_AGEMA_signal_5890, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5705, new_AGEMA_signal_5704, RoundKeyOutput[94]}), .a ({new_AGEMA_signal_9841, new_AGEMA_signal_9837, new_AGEMA_signal_9833}), .c ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, RoundKeyOutput[95]}), .a ({new_AGEMA_signal_9853, new_AGEMA_signal_9849, new_AGEMA_signal_9845}), .c ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_4907, new_AGEMA_signal_4906, RoundKeyOutput[96]}), .a ({new_AGEMA_signal_9865, new_AGEMA_signal_9861, new_AGEMA_signal_9857}), .c ({new_AGEMA_signal_4979, new_AGEMA_signal_4978, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, RoundKeyOutput[97]}), .a ({new_AGEMA_signal_9877, new_AGEMA_signal_9873, new_AGEMA_signal_9869}), .c ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, RoundKeyOutput[98]}), .a ({new_AGEMA_signal_9889, new_AGEMA_signal_9885, new_AGEMA_signal_9881}), .c ({new_AGEMA_signal_5185, new_AGEMA_signal_5184, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundKeyOutput[99]}), .a ({new_AGEMA_signal_9901, new_AGEMA_signal_9897, new_AGEMA_signal_9893}), .c ({new_AGEMA_signal_5189, new_AGEMA_signal_5188, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, RoundKeyOutput[100]}), .a ({new_AGEMA_signal_9913, new_AGEMA_signal_9909, new_AGEMA_signal_9905}), .c ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, RoundKeyOutput[101]}), .a ({new_AGEMA_signal_9925, new_AGEMA_signal_9921, new_AGEMA_signal_9917}), .c ({new_AGEMA_signal_5197, new_AGEMA_signal_5196, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5069, new_AGEMA_signal_5068, RoundKeyOutput[102]}), .a ({new_AGEMA_signal_9937, new_AGEMA_signal_9933, new_AGEMA_signal_9929}), .c ({new_AGEMA_signal_5201, new_AGEMA_signal_5200, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, RoundKeyOutput[103]}), .a ({new_AGEMA_signal_9949, new_AGEMA_signal_9945, new_AGEMA_signal_9941}), .c ({new_AGEMA_signal_5205, new_AGEMA_signal_5204, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, RoundKeyOutput[104]}), .a ({new_AGEMA_signal_9961, new_AGEMA_signal_9957, new_AGEMA_signal_9953}), .c ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, RoundKeyOutput[105]}), .a ({new_AGEMA_signal_9973, new_AGEMA_signal_9969, new_AGEMA_signal_9965}), .c ({new_AGEMA_signal_5209, new_AGEMA_signal_5208, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKeyOutput[106]}), .a ({new_AGEMA_signal_9985, new_AGEMA_signal_9981, new_AGEMA_signal_9977}), .c ({new_AGEMA_signal_5213, new_AGEMA_signal_5212, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, RoundKeyOutput[107]}), .a ({new_AGEMA_signal_9997, new_AGEMA_signal_9993, new_AGEMA_signal_9989}), .c ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, RoundKeyOutput[108]}), .a ({new_AGEMA_signal_10009, new_AGEMA_signal_10005, new_AGEMA_signal_10001}), .c ({new_AGEMA_signal_5221, new_AGEMA_signal_5220, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundKeyOutput[109]}), .a ({new_AGEMA_signal_10021, new_AGEMA_signal_10017, new_AGEMA_signal_10013}), .c ({new_AGEMA_signal_5225, new_AGEMA_signal_5224, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, RoundKeyOutput[110]}), .a ({new_AGEMA_signal_10033, new_AGEMA_signal_10029, new_AGEMA_signal_10025}), .c ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, RoundKeyOutput[111]}), .a ({new_AGEMA_signal_10045, new_AGEMA_signal_10041, new_AGEMA_signal_10037}), .c ({new_AGEMA_signal_5233, new_AGEMA_signal_5232, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, RoundKeyOutput[112]}), .a ({new_AGEMA_signal_10057, new_AGEMA_signal_10053, new_AGEMA_signal_10049}), .c ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5087, new_AGEMA_signal_5086, RoundKeyOutput[113]}), .a ({new_AGEMA_signal_10069, new_AGEMA_signal_10065, new_AGEMA_signal_10061}), .c ({new_AGEMA_signal_5237, new_AGEMA_signal_5236, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, RoundKeyOutput[114]}), .a ({new_AGEMA_signal_10081, new_AGEMA_signal_10077, new_AGEMA_signal_10073}), .c ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, RoundKeyOutput[115]}), .a ({new_AGEMA_signal_10093, new_AGEMA_signal_10089, new_AGEMA_signal_10085}), .c ({new_AGEMA_signal_5245, new_AGEMA_signal_5244, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKeyOutput[116]}), .a ({new_AGEMA_signal_10105, new_AGEMA_signal_10101, new_AGEMA_signal_10097}), .c ({new_AGEMA_signal_5249, new_AGEMA_signal_5248, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, RoundKeyOutput[117]}), .a ({new_AGEMA_signal_10117, new_AGEMA_signal_10113, new_AGEMA_signal_10109}), .c ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, RoundKeyOutput[118]}), .a ({new_AGEMA_signal_10129, new_AGEMA_signal_10125, new_AGEMA_signal_10121}), .c ({new_AGEMA_signal_5257, new_AGEMA_signal_5256, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundKeyOutput[119]}), .a ({new_AGEMA_signal_10141, new_AGEMA_signal_10137, new_AGEMA_signal_10133}), .c ({new_AGEMA_signal_5261, new_AGEMA_signal_5260, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, RoundKeyOutput[120]}), .a ({new_AGEMA_signal_10153, new_AGEMA_signal_10149, new_AGEMA_signal_10145}), .c ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKeyOutput[121]}), .a ({new_AGEMA_signal_10165, new_AGEMA_signal_10161, new_AGEMA_signal_10157}), .c ({new_AGEMA_signal_5561, new_AGEMA_signal_5560, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5383, new_AGEMA_signal_5382, RoundKeyOutput[122]}), .a ({new_AGEMA_signal_10177, new_AGEMA_signal_10173, new_AGEMA_signal_10169}), .c ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, RoundKeyOutput[123]}), .a ({new_AGEMA_signal_10189, new_AGEMA_signal_10185, new_AGEMA_signal_10181}), .c ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundKeyOutput[124]}), .a ({new_AGEMA_signal_10201, new_AGEMA_signal_10197, new_AGEMA_signal_10193}), .c ({new_AGEMA_signal_5573, new_AGEMA_signal_5572, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5389, new_AGEMA_signal_5388, RoundKeyOutput[125]}), .a ({new_AGEMA_signal_10213, new_AGEMA_signal_10209, new_AGEMA_signal_10205}), .c ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, RoundKeyOutput[126]}), .a ({new_AGEMA_signal_10225, new_AGEMA_signal_10221, new_AGEMA_signal_10217}), .c ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_7245), .b ({new_AGEMA_signal_5393, new_AGEMA_signal_5392, RoundKeyOutput[127]}), .a ({new_AGEMA_signal_10237, new_AGEMA_signal_10233, new_AGEMA_signal_10229}), .c ({new_AGEMA_signal_5585, new_AGEMA_signal_5584, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_10249, new_AGEMA_signal_10245, new_AGEMA_signal_10241}), .b ({new_AGEMA_signal_5269, new_AGEMA_signal_5268, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, KeyExpansionOutput[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_10261, new_AGEMA_signal_10257, new_AGEMA_signal_10253}), .b ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_5267, new_AGEMA_signal_5266, KeyExpansionOutput[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_10273, new_AGEMA_signal_10269, new_AGEMA_signal_10265}), .b ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, KeyExpansionOutput[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_10285, new_AGEMA_signal_10281, new_AGEMA_signal_10277}), .b ({new_AGEMA_signal_5273, new_AGEMA_signal_5272, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_5591, new_AGEMA_signal_5590, KeyExpansionOutput[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_10297, new_AGEMA_signal_10293, new_AGEMA_signal_10289}), .b ({new_AGEMA_signal_5275, new_AGEMA_signal_5274, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, KeyExpansionOutput[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_10309, new_AGEMA_signal_10305, new_AGEMA_signal_10301}), .b ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, KeyExpansionOutput[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_10321, new_AGEMA_signal_10317, new_AGEMA_signal_10313}), .b ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_5269, new_AGEMA_signal_5268, KeyExpansionOutput[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_10333, new_AGEMA_signal_10329, new_AGEMA_signal_10325}), .b ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyExpansionOutput[73]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_10345, new_AGEMA_signal_10341, new_AGEMA_signal_10337}), .b ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, KeyExpansionOutput[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_10357, new_AGEMA_signal_10353, new_AGEMA_signal_10349}), .b ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyExpansionOutput[72]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_10369, new_AGEMA_signal_10365, new_AGEMA_signal_10361}), .b ({new_AGEMA_signal_5279, new_AGEMA_signal_5278, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_5597, new_AGEMA_signal_5596, KeyExpansionOutput[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_10381, new_AGEMA_signal_10377, new_AGEMA_signal_10373}), .b ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, KeyExpansionOutput[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_10393, new_AGEMA_signal_10389, new_AGEMA_signal_10385}), .b ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, KeyExpansionOutput[71]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_10405, new_AGEMA_signal_10401, new_AGEMA_signal_10397}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_5273, new_AGEMA_signal_5272, KeyExpansionOutput[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_10417, new_AGEMA_signal_10413, new_AGEMA_signal_10409}), .b ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyExpansionOutput[70]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_10429, new_AGEMA_signal_10425, new_AGEMA_signal_10421}), .b ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_5275, new_AGEMA_signal_5274, KeyExpansionOutput[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_10441, new_AGEMA_signal_10437, new_AGEMA_signal_10433}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, KeyExpansionOutput[69]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_10453, new_AGEMA_signal_10449, new_AGEMA_signal_10445}), .b ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, KeyExpansionOutput[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_10465, new_AGEMA_signal_10461, new_AGEMA_signal_10457}), .b ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, KeyExpansionOutput[68]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_10477, new_AGEMA_signal_10473, new_AGEMA_signal_10469}), .b ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_5279, new_AGEMA_signal_5278, KeyExpansionOutput[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_10489, new_AGEMA_signal_10485, new_AGEMA_signal_10481}), .b ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyExpansionOutput[67]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_10501, new_AGEMA_signal_10497, new_AGEMA_signal_10493}), .b ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyExpansionOutput[99]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_10513, new_AGEMA_signal_10509, new_AGEMA_signal_10505}), .b ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, KeyExpansionOutput[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_10525, new_AGEMA_signal_10521, new_AGEMA_signal_10517}), .b ({new_AGEMA_signal_5281, new_AGEMA_signal_5280, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, KeyExpansionOutput[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_10537, new_AGEMA_signal_10533, new_AGEMA_signal_10529}), .b ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_5281, new_AGEMA_signal_5280, KeyExpansionOutput[95]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_10549, new_AGEMA_signal_10545, new_AGEMA_signal_10541}), .b ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_5903, new_AGEMA_signal_5902, KeyExpansionOutput[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_10561, new_AGEMA_signal_10557, new_AGEMA_signal_10553}), .b ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, KeyExpansionOutput[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_10573, new_AGEMA_signal_10569, new_AGEMA_signal_10565}), .b ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, KeyExpansionOutput[94]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_10585, new_AGEMA_signal_10581, new_AGEMA_signal_10577}), .b ({new_AGEMA_signal_5285, new_AGEMA_signal_5284, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_5603, new_AGEMA_signal_5602, KeyExpansionOutput[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_10597, new_AGEMA_signal_10593, new_AGEMA_signal_10589}), .b ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_5285, new_AGEMA_signal_5284, KeyExpansionOutput[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_10609, new_AGEMA_signal_10605, new_AGEMA_signal_10601}), .b ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, KeyExpansionOutput[66]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_10621, new_AGEMA_signal_10617, new_AGEMA_signal_10613}), .b ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyExpansionOutput[98]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_10633, new_AGEMA_signal_10629, new_AGEMA_signal_10625}), .b ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, KeyExpansionOutput[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_10645, new_AGEMA_signal_10641, new_AGEMA_signal_10637}), .b ({new_AGEMA_signal_5287, new_AGEMA_signal_5286, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, KeyExpansionOutput[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_10657, new_AGEMA_signal_10653, new_AGEMA_signal_10649}), .b ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_5287, new_AGEMA_signal_5286, KeyExpansionOutput[93]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_10669, new_AGEMA_signal_10665, new_AGEMA_signal_10661}), .b ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, KeyExpansionOutput[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_10681, new_AGEMA_signal_10677, new_AGEMA_signal_10673}), .b ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, KeyExpansionOutput[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_10693, new_AGEMA_signal_10689, new_AGEMA_signal_10685}), .b ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, KeyExpansionOutput[92]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_10705, new_AGEMA_signal_10701, new_AGEMA_signal_10697}), .b ({new_AGEMA_signal_5609, new_AGEMA_signal_5608, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_5909, new_AGEMA_signal_5908, KeyExpansionOutput[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_10717, new_AGEMA_signal_10713, new_AGEMA_signal_10709}), .b ({new_AGEMA_signal_5291, new_AGEMA_signal_5290, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_5609, new_AGEMA_signal_5608, KeyExpansionOutput[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_10729, new_AGEMA_signal_10725, new_AGEMA_signal_10721}), .b ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_5291, new_AGEMA_signal_5290, KeyExpansionOutput[91]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_10741, new_AGEMA_signal_10737, new_AGEMA_signal_10733}), .b ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, KeyExpansionOutput[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_10753, new_AGEMA_signal_10749, new_AGEMA_signal_10745}), .b ({new_AGEMA_signal_5293, new_AGEMA_signal_5292, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, KeyExpansionOutput[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_10765, new_AGEMA_signal_10761, new_AGEMA_signal_10757}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_5293, new_AGEMA_signal_5292, KeyExpansionOutput[90]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_10777, new_AGEMA_signal_10773, new_AGEMA_signal_10769}), .b ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, KeyExpansionOutput[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_10789, new_AGEMA_signal_10785, new_AGEMA_signal_10781}), .b ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, KeyExpansionOutput[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_10801, new_AGEMA_signal_10797, new_AGEMA_signal_10793}), .b ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, KeyExpansionOutput[89]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_10813, new_AGEMA_signal_10809, new_AGEMA_signal_10805}), .b ({new_AGEMA_signal_5297, new_AGEMA_signal_5296, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_5615, new_AGEMA_signal_5614, KeyExpansionOutput[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_10825, new_AGEMA_signal_10821, new_AGEMA_signal_10817}), .b ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_5297, new_AGEMA_signal_5296, KeyExpansionOutput[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_10837, new_AGEMA_signal_10833, new_AGEMA_signal_10829}), .b ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, KeyExpansionOutput[88]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_10849, new_AGEMA_signal_10845, new_AGEMA_signal_10841}), .b ({new_AGEMA_signal_5299, new_AGEMA_signal_5298, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, KeyExpansionOutput[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_10861, new_AGEMA_signal_10857, new_AGEMA_signal_10853}), .b ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_5299, new_AGEMA_signal_5298, KeyExpansionOutput[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_10873, new_AGEMA_signal_10869, new_AGEMA_signal_10865}), .b ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyExpansionOutput[87]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_10885, new_AGEMA_signal_10881, new_AGEMA_signal_10877}), .b ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_5619, new_AGEMA_signal_5618, KeyExpansionOutput[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_10897, new_AGEMA_signal_10893, new_AGEMA_signal_10889}), .b ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, KeyExpansionOutput[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_10909, new_AGEMA_signal_10905, new_AGEMA_signal_10901}), .b ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, KeyExpansionOutput[86]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_10921, new_AGEMA_signal_10917, new_AGEMA_signal_10913}), .b ({new_AGEMA_signal_5303, new_AGEMA_signal_5302, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_5621, new_AGEMA_signal_5620, KeyExpansionOutput[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_10933, new_AGEMA_signal_10929, new_AGEMA_signal_10925}), .b ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_5303, new_AGEMA_signal_5302, KeyExpansionOutput[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_10945, new_AGEMA_signal_10941, new_AGEMA_signal_10937}), .b ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, KeyExpansionOutput[85]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_10957, new_AGEMA_signal_10953, new_AGEMA_signal_10949}), .b ({new_AGEMA_signal_5305, new_AGEMA_signal_5304, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, KeyExpansionOutput[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_10969, new_AGEMA_signal_10965, new_AGEMA_signal_10961}), .b ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_5305, new_AGEMA_signal_5304, KeyExpansionOutput[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_10981, new_AGEMA_signal_10977, new_AGEMA_signal_10973}), .b ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyExpansionOutput[84]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_10993, new_AGEMA_signal_10989, new_AGEMA_signal_10985}), .b ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, KeyExpansionOutput[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_11005, new_AGEMA_signal_11001, new_AGEMA_signal_10997}), .b ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, KeyExpansionOutput[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_11017, new_AGEMA_signal_11013, new_AGEMA_signal_11009}), .b ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, KeyExpansionOutput[65]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_11029, new_AGEMA_signal_11025, new_AGEMA_signal_11021}), .b ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyExpansionOutput[97]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_11041, new_AGEMA_signal_11037, new_AGEMA_signal_11033}), .b ({new_AGEMA_signal_5309, new_AGEMA_signal_5308, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_5627, new_AGEMA_signal_5626, KeyExpansionOutput[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_11053, new_AGEMA_signal_11049, new_AGEMA_signal_11045}), .b ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_5309, new_AGEMA_signal_5308, KeyExpansionOutput[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_11065, new_AGEMA_signal_11061, new_AGEMA_signal_11057}), .b ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, KeyExpansionOutput[83]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_11077, new_AGEMA_signal_11073, new_AGEMA_signal_11069}), .b ({new_AGEMA_signal_5311, new_AGEMA_signal_5310, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, KeyExpansionOutput[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_11089, new_AGEMA_signal_11085, new_AGEMA_signal_11081}), .b ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_5311, new_AGEMA_signal_5310, KeyExpansionOutput[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_11101, new_AGEMA_signal_11097, new_AGEMA_signal_11093}), .b ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyExpansionOutput[82]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_11113, new_AGEMA_signal_11109, new_AGEMA_signal_11105}), .b ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, KeyExpansionOutput[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_11125, new_AGEMA_signal_11121, new_AGEMA_signal_11117}), .b ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, KeyExpansionOutput[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_11137, new_AGEMA_signal_11133, new_AGEMA_signal_11129}), .b ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, KeyExpansionOutput[81]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_11149, new_AGEMA_signal_11145, new_AGEMA_signal_11141}), .b ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_5315, new_AGEMA_signal_5314, KeyExpansionOutput[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_11161, new_AGEMA_signal_11157, new_AGEMA_signal_11153}), .b ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, KeyExpansionOutput[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_11173, new_AGEMA_signal_11169, new_AGEMA_signal_11165}), .b ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyExpansionOutput[80]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_11185, new_AGEMA_signal_11181, new_AGEMA_signal_11177}), .b ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_5633, new_AGEMA_signal_5632, KeyExpansionOutput[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_11197, new_AGEMA_signal_11193, new_AGEMA_signal_11189}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, KeyExpansionOutput[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_11209, new_AGEMA_signal_11205, new_AGEMA_signal_11201}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyExpansionOutput[79]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_11221, new_AGEMA_signal_11217, new_AGEMA_signal_11213}), .b ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, KeyExpansionOutput[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_11233, new_AGEMA_signal_11229, new_AGEMA_signal_11225}), .b ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyExpansionOutput[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_11245, new_AGEMA_signal_11241, new_AGEMA_signal_11237}), .b ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, KeyExpansionOutput[78]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_11257, new_AGEMA_signal_11253, new_AGEMA_signal_11249}), .b ({new_AGEMA_signal_5321, new_AGEMA_signal_5320, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, KeyExpansionOutput[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_11269, new_AGEMA_signal_11265, new_AGEMA_signal_11261}), .b ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_5321, new_AGEMA_signal_5320, KeyExpansionOutput[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_11281, new_AGEMA_signal_11277, new_AGEMA_signal_11273}), .b ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyExpansionOutput[77]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_11293, new_AGEMA_signal_11289, new_AGEMA_signal_11285}), .b ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_5639, new_AGEMA_signal_5638, KeyExpansionOutput[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_11305, new_AGEMA_signal_11301, new_AGEMA_signal_11297}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, KeyExpansionOutput[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_11317, new_AGEMA_signal_11313, new_AGEMA_signal_11309}), .b ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyExpansionOutput[76]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_11329, new_AGEMA_signal_11325, new_AGEMA_signal_11321}), .b ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, KeyExpansionOutput[127]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_11341, new_AGEMA_signal_11337, new_AGEMA_signal_11333}), .b ({new_AGEMA_signal_4895, new_AGEMA_signal_4894, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, KeyExpansionOutput[126]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_11353, new_AGEMA_signal_11349, new_AGEMA_signal_11345}), .b ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, KeyExpansionOutput[125]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_11365, new_AGEMA_signal_11361, new_AGEMA_signal_11357}), .b ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, KeyExpansionOutput[124]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_11377, new_AGEMA_signal_11373, new_AGEMA_signal_11369}), .b ({new_AGEMA_signal_4901, new_AGEMA_signal_4900, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, KeyExpansionOutput[123]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_11389, new_AGEMA_signal_11385, new_AGEMA_signal_11381}), .b ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, KeyExpansionOutput[122]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_11401, new_AGEMA_signal_11397, new_AGEMA_signal_11393}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, KeyExpansionOutput[121]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_11413, new_AGEMA_signal_11409, new_AGEMA_signal_11405}), .b ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyExpansionOutput[120]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_11425, new_AGEMA_signal_11421, new_AGEMA_signal_11417}), .b ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, KeyExpansionOutput[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_11437, new_AGEMA_signal_11433, new_AGEMA_signal_11429}), .b ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyExpansionOutput[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_11449, new_AGEMA_signal_11445, new_AGEMA_signal_11441}), .b ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, KeyExpansionOutput[75]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_11461, new_AGEMA_signal_11457, new_AGEMA_signal_11453}), .b ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyExpansionOutput[119]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_11473, new_AGEMA_signal_11469, new_AGEMA_signal_11465}), .b ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyExpansionOutput[118]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_11485, new_AGEMA_signal_11481, new_AGEMA_signal_11477}), .b ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, KeyExpansionOutput[117]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_11497, new_AGEMA_signal_11493, new_AGEMA_signal_11489}), .b ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, KeyExpansionOutput[116]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_11509, new_AGEMA_signal_11505, new_AGEMA_signal_11501}), .b ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyExpansionOutput[115]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_11521, new_AGEMA_signal_11517, new_AGEMA_signal_11513}), .b ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, KeyExpansionOutput[114]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_11533, new_AGEMA_signal_11529, new_AGEMA_signal_11525}), .b ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyExpansionOutput[113]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_11545, new_AGEMA_signal_11541, new_AGEMA_signal_11537}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyExpansionOutput[112]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_11557, new_AGEMA_signal_11553, new_AGEMA_signal_11549}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyExpansionOutput[111]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_11569, new_AGEMA_signal_11565, new_AGEMA_signal_11561}), .b ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyExpansionOutput[110]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_11581, new_AGEMA_signal_11577, new_AGEMA_signal_11573}), .b ({new_AGEMA_signal_5327, new_AGEMA_signal_5326, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, KeyExpansionOutput[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_11593, new_AGEMA_signal_11589, new_AGEMA_signal_11585}), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_5327, new_AGEMA_signal_5326, KeyExpansionOutput[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_11605, new_AGEMA_signal_11601, new_AGEMA_signal_11597}), .b ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, KeyExpansionOutput[74]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_11617, new_AGEMA_signal_11613, new_AGEMA_signal_11609}), .b ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyExpansionOutput[109]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_11629, new_AGEMA_signal_11625, new_AGEMA_signal_11621}), .b ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyExpansionOutput[108]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_11641, new_AGEMA_signal_11637, new_AGEMA_signal_11633}), .b ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyExpansionOutput[107]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_11653, new_AGEMA_signal_11649, new_AGEMA_signal_11645}), .b ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyExpansionOutput[106]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_11665, new_AGEMA_signal_11661, new_AGEMA_signal_11657}), .b ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyExpansionOutput[105]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_11677, new_AGEMA_signal_11673, new_AGEMA_signal_11669}), .b ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyExpansionOutput[104]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_11689, new_AGEMA_signal_11685, new_AGEMA_signal_11681}), .b ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, KeyExpansionOutput[103]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_11701, new_AGEMA_signal_11697, new_AGEMA_signal_11693}), .b ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, KeyExpansionOutput[102]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_11713, new_AGEMA_signal_11709, new_AGEMA_signal_11705}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyExpansionOutput[101]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_11725, new_AGEMA_signal_11721, new_AGEMA_signal_11717}), .b ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, KeyExpansionOutput[100]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_11737, new_AGEMA_signal_11733, new_AGEMA_signal_11729}), .b ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_5329, new_AGEMA_signal_5328, KeyExpansionOutput[0]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_11749, new_AGEMA_signal_11745, new_AGEMA_signal_11741}), .b ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, KeyExpansionOutput[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_11761, new_AGEMA_signal_11757, new_AGEMA_signal_11753}), .b ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, KeyExpansionOutput[64]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_11773, new_AGEMA_signal_11769, new_AGEMA_signal_11765}), .b ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyExpansionOutput[96]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11777}), .b ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11781}), .b ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_4895, new_AGEMA_signal_4894, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11785}), .b ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11789}), .b ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11793}), .b ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, SubBytesOutput[3]}), .c ({new_AGEMA_signal_4901, new_AGEMA_signal_4900, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11797}), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, SubBytesOutput[2]}), .c ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11801}), .b ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({1'b0, 1'b0, new_AGEMA_signal_11805}), .b ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, SubBytesOutput[0]}), .c ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, KeyExpansionIns_tmp[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_0_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11737, new_AGEMA_signal_11733, new_AGEMA_signal_11729}), .a ({new_AGEMA_signal_5329, new_AGEMA_signal_5328, KeyExpansionOutput[0]}), .c ({new_AGEMA_signal_5645, new_AGEMA_signal_5644, RoundKeyOutput[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_1_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10993, new_AGEMA_signal_10989, new_AGEMA_signal_10985}), .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, KeyExpansionOutput[1]}), .c ({new_AGEMA_signal_5915, new_AGEMA_signal_5914, RoundKeyOutput[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_2_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10585, new_AGEMA_signal_10581, new_AGEMA_signal_10577}), .a ({new_AGEMA_signal_5603, new_AGEMA_signal_5602, KeyExpansionOutput[2]}), .c ({new_AGEMA_signal_5917, new_AGEMA_signal_5916, RoundKeyOutput[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_3_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10369, new_AGEMA_signal_10365, new_AGEMA_signal_10361}), .a ({new_AGEMA_signal_5597, new_AGEMA_signal_5596, KeyExpansionOutput[3]}), .c ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, RoundKeyOutput[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_4_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10309, new_AGEMA_signal_10305, new_AGEMA_signal_10301}), .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, KeyExpansionOutput[4]}), .c ({new_AGEMA_signal_5921, new_AGEMA_signal_5920, RoundKeyOutput[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_5_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10297, new_AGEMA_signal_10293, new_AGEMA_signal_10289}), .a ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, KeyExpansionOutput[5]}), .c ({new_AGEMA_signal_5923, new_AGEMA_signal_5922, RoundKeyOutput[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_6_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10285, new_AGEMA_signal_10281, new_AGEMA_signal_10277}), .a ({new_AGEMA_signal_5591, new_AGEMA_signal_5590, KeyExpansionOutput[6]}), .c ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, RoundKeyOutput[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_7_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10273, new_AGEMA_signal_10269, new_AGEMA_signal_10265}), .a ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, KeyExpansionOutput[7]}), .c ({new_AGEMA_signal_5927, new_AGEMA_signal_5926, RoundKeyOutput[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_8_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_10261, new_AGEMA_signal_10257, new_AGEMA_signal_10253}), .a ({new_AGEMA_signal_5267, new_AGEMA_signal_5266, KeyExpansionOutput[8]}), .c ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, RoundKeyOutput[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_9_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10249, new_AGEMA_signal_10245, new_AGEMA_signal_10241}), .a ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, KeyExpansionOutput[9]}), .c ({new_AGEMA_signal_5929, new_AGEMA_signal_5928, RoundKeyOutput[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_10_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11581, new_AGEMA_signal_11577, new_AGEMA_signal_11573}), .a ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, KeyExpansionOutput[10]}), .c ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, RoundKeyOutput[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_11_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11425, new_AGEMA_signal_11421, new_AGEMA_signal_11417}), .a ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, KeyExpansionOutput[11]}), .c ({new_AGEMA_signal_5933, new_AGEMA_signal_5932, RoundKeyOutput[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_12_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_11293, new_AGEMA_signal_11289, new_AGEMA_signal_11285}), .a ({new_AGEMA_signal_5639, new_AGEMA_signal_5638, KeyExpansionOutput[12]}), .c ({new_AGEMA_signal_5935, new_AGEMA_signal_5934, RoundKeyOutput[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_13_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11257, new_AGEMA_signal_11253, new_AGEMA_signal_11249}), .a ({new_AGEMA_signal_5637, new_AGEMA_signal_5636, KeyExpansionOutput[13]}), .c ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, RoundKeyOutput[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_14_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_11221, new_AGEMA_signal_11217, new_AGEMA_signal_11213}), .a ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, KeyExpansionOutput[14]}), .c ({new_AGEMA_signal_5939, new_AGEMA_signal_5938, RoundKeyOutput[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_15_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_11185, new_AGEMA_signal_11181, new_AGEMA_signal_11177}), .a ({new_AGEMA_signal_5633, new_AGEMA_signal_5632, KeyExpansionOutput[15]}), .c ({new_AGEMA_signal_5941, new_AGEMA_signal_5940, RoundKeyOutput[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_16_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11149, new_AGEMA_signal_11145, new_AGEMA_signal_11141}), .a ({new_AGEMA_signal_5315, new_AGEMA_signal_5314, KeyExpansionOutput[16]}), .c ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, RoundKeyOutput[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_17_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11113, new_AGEMA_signal_11109, new_AGEMA_signal_11105}), .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, KeyExpansionOutput[17]}), .c ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, RoundKeyOutput[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_18_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11077, new_AGEMA_signal_11073, new_AGEMA_signal_11069}), .a ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, KeyExpansionOutput[18]}), .c ({new_AGEMA_signal_5945, new_AGEMA_signal_5944, RoundKeyOutput[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_19_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11041, new_AGEMA_signal_11037, new_AGEMA_signal_11033}), .a ({new_AGEMA_signal_5627, new_AGEMA_signal_5626, KeyExpansionOutput[19]}), .c ({new_AGEMA_signal_5947, new_AGEMA_signal_5946, RoundKeyOutput[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_20_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10957, new_AGEMA_signal_10953, new_AGEMA_signal_10949}), .a ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, KeyExpansionOutput[20]}), .c ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, RoundKeyOutput[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_21_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10921, new_AGEMA_signal_10917, new_AGEMA_signal_10913}), .a ({new_AGEMA_signal_5621, new_AGEMA_signal_5620, KeyExpansionOutput[21]}), .c ({new_AGEMA_signal_5951, new_AGEMA_signal_5950, RoundKeyOutput[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_22_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_10885, new_AGEMA_signal_10881, new_AGEMA_signal_10877}), .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5618, KeyExpansionOutput[22]}), .c ({new_AGEMA_signal_5953, new_AGEMA_signal_5952, RoundKeyOutput[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_23_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10849, new_AGEMA_signal_10845, new_AGEMA_signal_10841}), .a ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, KeyExpansionOutput[23]}), .c ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, RoundKeyOutput[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_24_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10813, new_AGEMA_signal_10809, new_AGEMA_signal_10805}), .a ({new_AGEMA_signal_5615, new_AGEMA_signal_5614, KeyExpansionOutput[24]}), .c ({new_AGEMA_signal_5957, new_AGEMA_signal_5956, RoundKeyOutput[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_25_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10777, new_AGEMA_signal_10773, new_AGEMA_signal_10769}), .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, KeyExpansionOutput[25]}), .c ({new_AGEMA_signal_6193, new_AGEMA_signal_6192, RoundKeyOutput[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_26_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10741, new_AGEMA_signal_10737, new_AGEMA_signal_10733}), .a ({new_AGEMA_signal_5911, new_AGEMA_signal_5910, KeyExpansionOutput[26]}), .c ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, RoundKeyOutput[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_27_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10705, new_AGEMA_signal_10701, new_AGEMA_signal_10697}), .a ({new_AGEMA_signal_5909, new_AGEMA_signal_5908, KeyExpansionOutput[27]}), .c ({new_AGEMA_signal_6197, new_AGEMA_signal_6196, RoundKeyOutput[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_28_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_10669, new_AGEMA_signal_10665, new_AGEMA_signal_10661}), .a ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, KeyExpansionOutput[28]}), .c ({new_AGEMA_signal_6199, new_AGEMA_signal_6198, RoundKeyOutput[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_29_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_10633, new_AGEMA_signal_10629, new_AGEMA_signal_10625}), .a ({new_AGEMA_signal_5905, new_AGEMA_signal_5904, KeyExpansionOutput[29]}), .c ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, RoundKeyOutput[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_30_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10549, new_AGEMA_signal_10545, new_AGEMA_signal_10541}), .a ({new_AGEMA_signal_5903, new_AGEMA_signal_5902, KeyExpansionOutput[30]}), .c ({new_AGEMA_signal_6203, new_AGEMA_signal_6202, RoundKeyOutput[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_31_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10513, new_AGEMA_signal_10509, new_AGEMA_signal_10505}), .a ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, KeyExpansionOutput[31]}), .c ({new_AGEMA_signal_6205, new_AGEMA_signal_6204, RoundKeyOutput[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_32_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11749, new_AGEMA_signal_11745, new_AGEMA_signal_11741}), .a ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_5331, new_AGEMA_signal_5330, RoundKeyOutput[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_33_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11005, new_AGEMA_signal_11001, new_AGEMA_signal_10997}), .a ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKeyOutput[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_34_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10597, new_AGEMA_signal_10593, new_AGEMA_signal_10589}), .a ({new_AGEMA_signal_5285, new_AGEMA_signal_5284, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, RoundKeyOutput[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_35_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10477, new_AGEMA_signal_10473, new_AGEMA_signal_10469}), .a ({new_AGEMA_signal_5279, new_AGEMA_signal_5278, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_5655, new_AGEMA_signal_5654, RoundKeyOutput[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_36_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10453, new_AGEMA_signal_10449, new_AGEMA_signal_10445}), .a ({new_AGEMA_signal_5277, new_AGEMA_signal_5276, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundKeyOutput[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_37_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_10429, new_AGEMA_signal_10425, new_AGEMA_signal_10421}), .a ({new_AGEMA_signal_5275, new_AGEMA_signal_5274, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, RoundKeyOutput[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_38_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10405, new_AGEMA_signal_10401, new_AGEMA_signal_10397}), .a ({new_AGEMA_signal_5273, new_AGEMA_signal_5272, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, RoundKeyOutput[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_39_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10381, new_AGEMA_signal_10377, new_AGEMA_signal_10373}), .a ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_5663, new_AGEMA_signal_5662, RoundKeyOutput[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_40_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10345, new_AGEMA_signal_10341, new_AGEMA_signal_10337}), .a ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundKeyOutput[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_41_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10321, new_AGEMA_signal_10317, new_AGEMA_signal_10313}), .a ({new_AGEMA_signal_5269, new_AGEMA_signal_5268, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, RoundKeyOutput[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_42_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11593, new_AGEMA_signal_11589, new_AGEMA_signal_11585}), .a ({new_AGEMA_signal_5327, new_AGEMA_signal_5326, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, RoundKeyOutput[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_43_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11437, new_AGEMA_signal_11433, new_AGEMA_signal_11429}), .a ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKeyOutput[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_44_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11305, new_AGEMA_signal_11301, new_AGEMA_signal_11297}), .a ({new_AGEMA_signal_5323, new_AGEMA_signal_5322, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, RoundKeyOutput[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_45_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11269, new_AGEMA_signal_11265, new_AGEMA_signal_11261}), .a ({new_AGEMA_signal_5321, new_AGEMA_signal_5320, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_5673, new_AGEMA_signal_5672, RoundKeyOutput[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_46_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11233, new_AGEMA_signal_11229, new_AGEMA_signal_11225}), .a ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundKeyOutput[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_47_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11197, new_AGEMA_signal_11193, new_AGEMA_signal_11189}), .a ({new_AGEMA_signal_5317, new_AGEMA_signal_5316, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, RoundKeyOutput[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_48_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11161, new_AGEMA_signal_11157, new_AGEMA_signal_11153}), .a ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_5335, new_AGEMA_signal_5334, RoundKeyOutput[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_49_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11125, new_AGEMA_signal_11121, new_AGEMA_signal_11117}), .a ({new_AGEMA_signal_5313, new_AGEMA_signal_5312, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, RoundKeyOutput[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_50_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11089, new_AGEMA_signal_11085, new_AGEMA_signal_11081}), .a ({new_AGEMA_signal_5311, new_AGEMA_signal_5310, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_5681, new_AGEMA_signal_5680, RoundKeyOutput[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_51_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_11053, new_AGEMA_signal_11049, new_AGEMA_signal_11045}), .a ({new_AGEMA_signal_5309, new_AGEMA_signal_5308, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, RoundKeyOutput[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_52_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10969, new_AGEMA_signal_10965, new_AGEMA_signal_10961}), .a ({new_AGEMA_signal_5305, new_AGEMA_signal_5304, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, RoundKeyOutput[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_53_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10933, new_AGEMA_signal_10929, new_AGEMA_signal_10925}), .a ({new_AGEMA_signal_5303, new_AGEMA_signal_5302, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKeyOutput[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_54_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10897, new_AGEMA_signal_10893, new_AGEMA_signal_10889}), .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, RoundKeyOutput[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_55_U1 ( .s (new_AGEMA_signal_11829), .b ({new_AGEMA_signal_10861, new_AGEMA_signal_10857, new_AGEMA_signal_10853}), .a ({new_AGEMA_signal_5299, new_AGEMA_signal_5298, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_5691, new_AGEMA_signal_5690, RoundKeyOutput[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_56_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10825, new_AGEMA_signal_10821, new_AGEMA_signal_10817}), .a ({new_AGEMA_signal_5297, new_AGEMA_signal_5296, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundKeyOutput[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_57_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10789, new_AGEMA_signal_10785, new_AGEMA_signal_10781}), .a ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_5959, new_AGEMA_signal_5958, RoundKeyOutput[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_58_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10753, new_AGEMA_signal_10749, new_AGEMA_signal_10745}), .a ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, RoundKeyOutput[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_59_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10717, new_AGEMA_signal_10713, new_AGEMA_signal_10709}), .a ({new_AGEMA_signal_5609, new_AGEMA_signal_5608, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_5963, new_AGEMA_signal_5962, RoundKeyOutput[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_60_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10681, new_AGEMA_signal_10677, new_AGEMA_signal_10673}), .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_5965, new_AGEMA_signal_5964, RoundKeyOutput[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_61_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10645, new_AGEMA_signal_10641, new_AGEMA_signal_10637}), .a ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, RoundKeyOutput[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_62_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10561, new_AGEMA_signal_10557, new_AGEMA_signal_10553}), .a ({new_AGEMA_signal_5601, new_AGEMA_signal_5600, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_5969, new_AGEMA_signal_5968, RoundKeyOutput[62]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_63_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10525, new_AGEMA_signal_10521, new_AGEMA_signal_10517}), .a ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_5971, new_AGEMA_signal_5970, RoundKeyOutput[63]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_64_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_11761, new_AGEMA_signal_11757, new_AGEMA_signal_11753}), .a ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, RoundKeyOutput[64]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_65_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_11017, new_AGEMA_signal_11013, new_AGEMA_signal_11009}), .a ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, RoundKeyOutput[65]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_66_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10609, new_AGEMA_signal_10605, new_AGEMA_signal_10601}), .a ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_5339, new_AGEMA_signal_5338, RoundKeyOutput[66]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_67_U1 ( .s (new_AGEMA_signal_11825), .b ({new_AGEMA_signal_10489, new_AGEMA_signal_10485, new_AGEMA_signal_10481}), .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_5341, new_AGEMA_signal_5340, RoundKeyOutput[67]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_68_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10465, new_AGEMA_signal_10461, new_AGEMA_signal_10457}), .a ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, RoundKeyOutput[68]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_69_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10441, new_AGEMA_signal_10437, new_AGEMA_signal_10433}), .a ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKeyOutput[69]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_70_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10417, new_AGEMA_signal_10413, new_AGEMA_signal_10409}), .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_5347, new_AGEMA_signal_5346, RoundKeyOutput[70]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_71_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10393, new_AGEMA_signal_10389, new_AGEMA_signal_10385}), .a ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_5349, new_AGEMA_signal_5348, RoundKeyOutput[71]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_72_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10357, new_AGEMA_signal_10353, new_AGEMA_signal_10349}), .a ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, RoundKeyOutput[72]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_73_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_10333, new_AGEMA_signal_10329, new_AGEMA_signal_10325}), .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundKeyOutput[73]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_74_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11605, new_AGEMA_signal_11601, new_AGEMA_signal_11597}), .a ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_5353, new_AGEMA_signal_5352, RoundKeyOutput[74]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_75_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11449, new_AGEMA_signal_11445, new_AGEMA_signal_11441}), .a ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, RoundKeyOutput[75]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_76_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11317, new_AGEMA_signal_11313, new_AGEMA_signal_11309}), .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_5357, new_AGEMA_signal_5356, RoundKeyOutput[76]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_77_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11281, new_AGEMA_signal_11277, new_AGEMA_signal_11273}), .a ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_5359, new_AGEMA_signal_5358, RoundKeyOutput[77]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_78_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11245, new_AGEMA_signal_11241, new_AGEMA_signal_11237}), .a ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, RoundKeyOutput[78]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_79_U1 ( .s (new_AGEMA_signal_11821), .b ({new_AGEMA_signal_11209, new_AGEMA_signal_11205, new_AGEMA_signal_11201}), .a ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKeyOutput[79]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_80_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11173, new_AGEMA_signal_11169, new_AGEMA_signal_11165}), .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKeyOutput[80]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_81_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11137, new_AGEMA_signal_11133, new_AGEMA_signal_11129}), .a ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_5365, new_AGEMA_signal_5364, RoundKeyOutput[81]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_82_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11101, new_AGEMA_signal_11097, new_AGEMA_signal_11093}), .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_5367, new_AGEMA_signal_5366, RoundKeyOutput[82]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_83_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_11065, new_AGEMA_signal_11061, new_AGEMA_signal_11057}), .a ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundKeyOutput[83]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_84_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10981, new_AGEMA_signal_10977, new_AGEMA_signal_10973}), .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_5371, new_AGEMA_signal_5370, RoundKeyOutput[84]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_85_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10945, new_AGEMA_signal_10941, new_AGEMA_signal_10937}), .a ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, RoundKeyOutput[85]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_86_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10909, new_AGEMA_signal_10905, new_AGEMA_signal_10901}), .a ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_5375, new_AGEMA_signal_5374, RoundKeyOutput[86]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_87_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10873, new_AGEMA_signal_10869, new_AGEMA_signal_10865}), .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_5377, new_AGEMA_signal_5376, RoundKeyOutput[87]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_88_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10837, new_AGEMA_signal_10833, new_AGEMA_signal_10829}), .a ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, RoundKeyOutput[88]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_89_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10801, new_AGEMA_signal_10797, new_AGEMA_signal_10793}), .a ({new_AGEMA_signal_5295, new_AGEMA_signal_5294, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, RoundKeyOutput[89]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_90_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10765, new_AGEMA_signal_10761, new_AGEMA_signal_10757}), .a ({new_AGEMA_signal_5293, new_AGEMA_signal_5292, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, RoundKeyOutput[90]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_91_U1 ( .s (new_AGEMA_signal_11817), .b ({new_AGEMA_signal_10729, new_AGEMA_signal_10725, new_AGEMA_signal_10721}), .a ({new_AGEMA_signal_5291, new_AGEMA_signal_5290, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_5699, new_AGEMA_signal_5698, RoundKeyOutput[91]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_92_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10693, new_AGEMA_signal_10689, new_AGEMA_signal_10685}), .a ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, RoundKeyOutput[92]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_93_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10657, new_AGEMA_signal_10653, new_AGEMA_signal_10649}), .a ({new_AGEMA_signal_5287, new_AGEMA_signal_5286, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, RoundKeyOutput[93]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_94_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10573, new_AGEMA_signal_10569, new_AGEMA_signal_10565}), .a ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_5705, new_AGEMA_signal_5704, RoundKeyOutput[94]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_95_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10537, new_AGEMA_signal_10533, new_AGEMA_signal_10529}), .a ({new_AGEMA_signal_5281, new_AGEMA_signal_5280, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, RoundKeyOutput[95]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_96_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11773, new_AGEMA_signal_11769, new_AGEMA_signal_11765}), .a ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_4907, new_AGEMA_signal_4906, RoundKeyOutput[96]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_97_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11029, new_AGEMA_signal_11025, new_AGEMA_signal_11021}), .a ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, RoundKeyOutput[97]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_98_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10621, new_AGEMA_signal_10617, new_AGEMA_signal_10613}), .a ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, RoundKeyOutput[98]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_99_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_10501, new_AGEMA_signal_10497, new_AGEMA_signal_10493}), .a ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundKeyOutput[99]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_100_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11725, new_AGEMA_signal_11721, new_AGEMA_signal_11717}), .a ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, RoundKeyOutput[100]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_101_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11713, new_AGEMA_signal_11709, new_AGEMA_signal_11705}), .a ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, RoundKeyOutput[101]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_102_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11701, new_AGEMA_signal_11697, new_AGEMA_signal_11693}), .a ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_5069, new_AGEMA_signal_5068, RoundKeyOutput[102]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_103_U1 ( .s (new_AGEMA_signal_11813), .b ({new_AGEMA_signal_11689, new_AGEMA_signal_11685, new_AGEMA_signal_11681}), .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, RoundKeyOutput[103]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_104_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11677, new_AGEMA_signal_11673, new_AGEMA_signal_11669}), .a ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, RoundKeyOutput[104]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_105_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11665, new_AGEMA_signal_11661, new_AGEMA_signal_11657}), .a ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, RoundKeyOutput[105]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_106_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11653, new_AGEMA_signal_11649, new_AGEMA_signal_11645}), .a ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKeyOutput[106]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_107_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11641, new_AGEMA_signal_11637, new_AGEMA_signal_11633}), .a ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, RoundKeyOutput[107]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_108_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11629, new_AGEMA_signal_11625, new_AGEMA_signal_11621}), .a ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, RoundKeyOutput[108]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_109_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11617, new_AGEMA_signal_11613, new_AGEMA_signal_11609}), .a ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundKeyOutput[109]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_110_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11569, new_AGEMA_signal_11565, new_AGEMA_signal_11561}), .a ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, RoundKeyOutput[110]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_111_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11557, new_AGEMA_signal_11553, new_AGEMA_signal_11549}), .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, RoundKeyOutput[111]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_112_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11545, new_AGEMA_signal_11541, new_AGEMA_signal_11537}), .a ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, RoundKeyOutput[112]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_113_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11533, new_AGEMA_signal_11529, new_AGEMA_signal_11525}), .a ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_5087, new_AGEMA_signal_5086, RoundKeyOutput[113]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_114_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11521, new_AGEMA_signal_11517, new_AGEMA_signal_11513}), .a ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, RoundKeyOutput[114]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_115_U1 ( .s (new_AGEMA_signal_11809), .b ({new_AGEMA_signal_11509, new_AGEMA_signal_11505, new_AGEMA_signal_11501}), .a ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, RoundKeyOutput[115]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_116_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11497, new_AGEMA_signal_11493, new_AGEMA_signal_11489}), .a ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKeyOutput[116]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_117_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11485, new_AGEMA_signal_11481, new_AGEMA_signal_11477}), .a ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, RoundKeyOutput[117]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_118_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11473, new_AGEMA_signal_11469, new_AGEMA_signal_11465}), .a ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, RoundKeyOutput[118]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_119_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11461, new_AGEMA_signal_11457, new_AGEMA_signal_11453}), .a ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundKeyOutput[119]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_120_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11413, new_AGEMA_signal_11409, new_AGEMA_signal_11405}), .a ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, RoundKeyOutput[120]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_121_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11401, new_AGEMA_signal_11397, new_AGEMA_signal_11393}), .a ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKeyOutput[121]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_122_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11389, new_AGEMA_signal_11385, new_AGEMA_signal_11381}), .a ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_5383, new_AGEMA_signal_5382, RoundKeyOutput[122]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_123_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11377, new_AGEMA_signal_11373, new_AGEMA_signal_11369}), .a ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_5385, new_AGEMA_signal_5384, RoundKeyOutput[123]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_124_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11365, new_AGEMA_signal_11361, new_AGEMA_signal_11357}), .a ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundKeyOutput[124]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_125_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11353, new_AGEMA_signal_11349, new_AGEMA_signal_11345}), .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_5389, new_AGEMA_signal_5388, RoundKeyOutput[125]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_126_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11341, new_AGEMA_signal_11337, new_AGEMA_signal_11333}), .a ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, RoundKeyOutput[126]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) MuxKeyExpansion_mux_inst_127_U1 ( .s (new_AGEMA_signal_11833), .b ({new_AGEMA_signal_11329, new_AGEMA_signal_11325, new_AGEMA_signal_11321}), .a ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_5393, new_AGEMA_signal_5392, RoundKeyOutput[127]}) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_7244), .Q (new_AGEMA_signal_7245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_7248), .Q (new_AGEMA_signal_7249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_7252), .Q (new_AGEMA_signal_7253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_7256), .Q (new_AGEMA_signal_7257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_7260), .Q (new_AGEMA_signal_7261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_7264), .Q (new_AGEMA_signal_7265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_7268), .Q (new_AGEMA_signal_7269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_7272), .Q (new_AGEMA_signal_7273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_7276), .Q (new_AGEMA_signal_7277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_7280), .Q (new_AGEMA_signal_7281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_7284), .Q (new_AGEMA_signal_7285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_7288), .Q (new_AGEMA_signal_7289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_7292), .Q (new_AGEMA_signal_7293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_7296), .Q (new_AGEMA_signal_7297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_7300), .Q (new_AGEMA_signal_7301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_7304), .Q (new_AGEMA_signal_7305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_7308), .Q (new_AGEMA_signal_7309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_7312), .Q (new_AGEMA_signal_7313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_7316), .Q (new_AGEMA_signal_7317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_7320), .Q (new_AGEMA_signal_7321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_7324), .Q (new_AGEMA_signal_7325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_7328), .Q (new_AGEMA_signal_7329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_7332), .Q (new_AGEMA_signal_7333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_7336), .Q (new_AGEMA_signal_7337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_7340), .Q (new_AGEMA_signal_7341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_7344), .Q (new_AGEMA_signal_7345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_7348), .Q (new_AGEMA_signal_7349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_7352), .Q (new_AGEMA_signal_7353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_7356), .Q (new_AGEMA_signal_7357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_7360), .Q (new_AGEMA_signal_7361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_7364), .Q (new_AGEMA_signal_7365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_7368), .Q (new_AGEMA_signal_7369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_7372), .Q (new_AGEMA_signal_7373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_7376), .Q (new_AGEMA_signal_7377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_7380), .Q (new_AGEMA_signal_7381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_7384), .Q (new_AGEMA_signal_7385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_7388), .Q (new_AGEMA_signal_7389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_7392), .Q (new_AGEMA_signal_7393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_7396), .Q (new_AGEMA_signal_7397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_7400), .Q (new_AGEMA_signal_7401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_7404), .Q (new_AGEMA_signal_7405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_7408), .Q (new_AGEMA_signal_7409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_7412), .Q (new_AGEMA_signal_7413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_7416), .Q (new_AGEMA_signal_7417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_7420), .Q (new_AGEMA_signal_7421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_7424), .Q (new_AGEMA_signal_7425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_7428), .Q (new_AGEMA_signal_7429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_7432), .Q (new_AGEMA_signal_7433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_7436), .Q (new_AGEMA_signal_7437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_7440), .Q (new_AGEMA_signal_7441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_7445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_7449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_7453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_7457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_7461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_7465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_7469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_7472), .Q (new_AGEMA_signal_7473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_7477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_7480), .Q (new_AGEMA_signal_7481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_7485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_7489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_7493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_7497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_7501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_7504), .Q (new_AGEMA_signal_7505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_7509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_7512), .Q (new_AGEMA_signal_7513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_7517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_7520), .Q (new_AGEMA_signal_7521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_7524), .Q (new_AGEMA_signal_7525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_7529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_7532), .Q (new_AGEMA_signal_7533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_7537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_7540), .Q (new_AGEMA_signal_7541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_7544), .Q (new_AGEMA_signal_7545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_7548), .Q (new_AGEMA_signal_7549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_7552), .Q (new_AGEMA_signal_7553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_7556), .Q (new_AGEMA_signal_7557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_7560), .Q (new_AGEMA_signal_7561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_7564), .Q (new_AGEMA_signal_7565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_7568), .Q (new_AGEMA_signal_7569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_7572), .Q (new_AGEMA_signal_7573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_7576), .Q (new_AGEMA_signal_7577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_7580), .Q (new_AGEMA_signal_7581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_7584), .Q (new_AGEMA_signal_7585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_7589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_7592), .Q (new_AGEMA_signal_7593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_7596), .Q (new_AGEMA_signal_7597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_7600), .Q (new_AGEMA_signal_7601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_7604), .Q (new_AGEMA_signal_7605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_7608), .Q (new_AGEMA_signal_7609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_7612), .Q (new_AGEMA_signal_7613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_7617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_7620), .Q (new_AGEMA_signal_7621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_7624), .Q (new_AGEMA_signal_7625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_7628), .Q (new_AGEMA_signal_7629) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_8280), .Q (new_AGEMA_signal_8281) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_8284), .Q (new_AGEMA_signal_8285) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_8288), .Q (new_AGEMA_signal_8289) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_8292), .Q (new_AGEMA_signal_8293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_8296), .Q (new_AGEMA_signal_8297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_8300), .Q (new_AGEMA_signal_8301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_8304), .Q (new_AGEMA_signal_8305) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_8308), .Q (new_AGEMA_signal_8309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_8312), .Q (new_AGEMA_signal_8313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_8316), .Q (new_AGEMA_signal_8317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_8320), .Q (new_AGEMA_signal_8321) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_8324), .Q (new_AGEMA_signal_8325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_8328), .Q (new_AGEMA_signal_8329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_8332), .Q (new_AGEMA_signal_8333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_8336), .Q (new_AGEMA_signal_8337) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_8340), .Q (new_AGEMA_signal_8341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_8344), .Q (new_AGEMA_signal_8345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_8348), .Q (new_AGEMA_signal_8349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_8352), .Q (new_AGEMA_signal_8353) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_8356), .Q (new_AGEMA_signal_8357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_8360), .Q (new_AGEMA_signal_8361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_8364), .Q (new_AGEMA_signal_8365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_8368), .Q (new_AGEMA_signal_8369) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_8372), .Q (new_AGEMA_signal_8373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_8376), .Q (new_AGEMA_signal_8377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_8380), .Q (new_AGEMA_signal_8381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_8384), .Q (new_AGEMA_signal_8385) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_8388), .Q (new_AGEMA_signal_8389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_8392), .Q (new_AGEMA_signal_8393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_8396), .Q (new_AGEMA_signal_8397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_8400), .Q (new_AGEMA_signal_8401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_8404), .Q (new_AGEMA_signal_8405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_8408), .Q (new_AGEMA_signal_8409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_8412), .Q (new_AGEMA_signal_8413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_8416), .Q (new_AGEMA_signal_8417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_8420), .Q (new_AGEMA_signal_8421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_8424), .Q (new_AGEMA_signal_8425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_8428), .Q (new_AGEMA_signal_8429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_8432), .Q (new_AGEMA_signal_8433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_8436), .Q (new_AGEMA_signal_8437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_8440), .Q (new_AGEMA_signal_8441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_8444), .Q (new_AGEMA_signal_8445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_8448), .Q (new_AGEMA_signal_8449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_8452), .Q (new_AGEMA_signal_8453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_8456), .Q (new_AGEMA_signal_8457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_8460), .Q (new_AGEMA_signal_8461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_8464), .Q (new_AGEMA_signal_8465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_8468), .Q (new_AGEMA_signal_8469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_8472), .Q (new_AGEMA_signal_8473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_8476), .Q (new_AGEMA_signal_8477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_8480), .Q (new_AGEMA_signal_8481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_8484), .Q (new_AGEMA_signal_8485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_8488), .Q (new_AGEMA_signal_8489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_8492), .Q (new_AGEMA_signal_8493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_8496), .Q (new_AGEMA_signal_8497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_8500), .Q (new_AGEMA_signal_8501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_8504), .Q (new_AGEMA_signal_8505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_8508), .Q (new_AGEMA_signal_8509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_8512), .Q (new_AGEMA_signal_8513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_8516), .Q (new_AGEMA_signal_8517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_8520), .Q (new_AGEMA_signal_8521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_8524), .Q (new_AGEMA_signal_8525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_8528), .Q (new_AGEMA_signal_8529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_8532), .Q (new_AGEMA_signal_8533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_8536), .Q (new_AGEMA_signal_8537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_8540), .Q (new_AGEMA_signal_8541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_8544), .Q (new_AGEMA_signal_8545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_8548), .Q (new_AGEMA_signal_8549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_8552), .Q (new_AGEMA_signal_8553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_8556), .Q (new_AGEMA_signal_8557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_8560), .Q (new_AGEMA_signal_8561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_8564), .Q (new_AGEMA_signal_8565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_8568), .Q (new_AGEMA_signal_8569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_8572), .Q (new_AGEMA_signal_8573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_8576), .Q (new_AGEMA_signal_8577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_8580), .Q (new_AGEMA_signal_8581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_8584), .Q (new_AGEMA_signal_8585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_8588), .Q (new_AGEMA_signal_8589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_8592), .Q (new_AGEMA_signal_8593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_8596), .Q (new_AGEMA_signal_8597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_8600), .Q (new_AGEMA_signal_8601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_8604), .Q (new_AGEMA_signal_8605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_8608), .Q (new_AGEMA_signal_8609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_8612), .Q (new_AGEMA_signal_8613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_8616), .Q (new_AGEMA_signal_8617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_8620), .Q (new_AGEMA_signal_8621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_8624), .Q (new_AGEMA_signal_8625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_8628), .Q (new_AGEMA_signal_8629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_8632), .Q (new_AGEMA_signal_8633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_8636), .Q (new_AGEMA_signal_8637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_8640), .Q (new_AGEMA_signal_8641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_8644), .Q (new_AGEMA_signal_8645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_8648), .Q (new_AGEMA_signal_8649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_8652), .Q (new_AGEMA_signal_8653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_8656), .Q (new_AGEMA_signal_8657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_8660), .Q (new_AGEMA_signal_8661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_8664), .Q (new_AGEMA_signal_8665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_8668), .Q (new_AGEMA_signal_8669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_8672), .Q (new_AGEMA_signal_8673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_8676), .Q (new_AGEMA_signal_8677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_8680), .Q (new_AGEMA_signal_8681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_8684), .Q (new_AGEMA_signal_8685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_8688), .Q (new_AGEMA_signal_8689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_8692), .Q (new_AGEMA_signal_8693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_8696), .Q (new_AGEMA_signal_8697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_8700), .Q (new_AGEMA_signal_8701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_8704), .Q (new_AGEMA_signal_8705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_8708), .Q (new_AGEMA_signal_8709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_8712), .Q (new_AGEMA_signal_8713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_8716), .Q (new_AGEMA_signal_8717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_8720), .Q (new_AGEMA_signal_8721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_8724), .Q (new_AGEMA_signal_8725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_8728), .Q (new_AGEMA_signal_8729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_8732), .Q (new_AGEMA_signal_8733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_8736), .Q (new_AGEMA_signal_8737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_8740), .Q (new_AGEMA_signal_8741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_8744), .Q (new_AGEMA_signal_8745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_8748), .Q (new_AGEMA_signal_8749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_8752), .Q (new_AGEMA_signal_8753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_8756), .Q (new_AGEMA_signal_8757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_8760), .Q (new_AGEMA_signal_8761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_8764), .Q (new_AGEMA_signal_8765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_8768), .Q (new_AGEMA_signal_8769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_8772), .Q (new_AGEMA_signal_8773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_8776), .Q (new_AGEMA_signal_8777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_8780), .Q (new_AGEMA_signal_8781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_8784), .Q (new_AGEMA_signal_8785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_8788), .Q (new_AGEMA_signal_8789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_8792), .Q (new_AGEMA_signal_8793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_8796), .Q (new_AGEMA_signal_8797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_8800), .Q (new_AGEMA_signal_8801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_8804), .Q (new_AGEMA_signal_8805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_8808), .Q (new_AGEMA_signal_8809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_8812), .Q (new_AGEMA_signal_8813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_8816), .Q (new_AGEMA_signal_8817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_8820), .Q (new_AGEMA_signal_8821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_8824), .Q (new_AGEMA_signal_8825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_8828), .Q (new_AGEMA_signal_8829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_8832), .Q (new_AGEMA_signal_8833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_8836), .Q (new_AGEMA_signal_8837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_8840), .Q (new_AGEMA_signal_8841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_8844), .Q (new_AGEMA_signal_8845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_8848), .Q (new_AGEMA_signal_8849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_8852), .Q (new_AGEMA_signal_8853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_8856), .Q (new_AGEMA_signal_8857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_8860), .Q (new_AGEMA_signal_8861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_8864), .Q (new_AGEMA_signal_8865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_8868), .Q (new_AGEMA_signal_8869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_8872), .Q (new_AGEMA_signal_8873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_8876), .Q (new_AGEMA_signal_8877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_8880), .Q (new_AGEMA_signal_8881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_8884), .Q (new_AGEMA_signal_8885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_8888), .Q (new_AGEMA_signal_8889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_8892), .Q (new_AGEMA_signal_8893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_8896), .Q (new_AGEMA_signal_8897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_8900), .Q (new_AGEMA_signal_8901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_8904), .Q (new_AGEMA_signal_8905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_8908), .Q (new_AGEMA_signal_8909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_8912), .Q (new_AGEMA_signal_8913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_8916), .Q (new_AGEMA_signal_8917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_8920), .Q (new_AGEMA_signal_8921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_8924), .Q (new_AGEMA_signal_8925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_8928), .Q (new_AGEMA_signal_8929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_8932), .Q (new_AGEMA_signal_8933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_8936), .Q (new_AGEMA_signal_8937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_8940), .Q (new_AGEMA_signal_8941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_8944), .Q (new_AGEMA_signal_8945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_8948), .Q (new_AGEMA_signal_8949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_8952), .Q (new_AGEMA_signal_8953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_8956), .Q (new_AGEMA_signal_8957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_8960), .Q (new_AGEMA_signal_8961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_8964), .Q (new_AGEMA_signal_8965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_8968), .Q (new_AGEMA_signal_8969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_8972), .Q (new_AGEMA_signal_8973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_8976), .Q (new_AGEMA_signal_8977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_8980), .Q (new_AGEMA_signal_8981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_8984), .Q (new_AGEMA_signal_8985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_8988), .Q (new_AGEMA_signal_8989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_8992), .Q (new_AGEMA_signal_8993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_8996), .Q (new_AGEMA_signal_8997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_9000), .Q (new_AGEMA_signal_9001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_9004), .Q (new_AGEMA_signal_9005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_9008), .Q (new_AGEMA_signal_9009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_9012), .Q (new_AGEMA_signal_9013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_9016), .Q (new_AGEMA_signal_9017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_9020), .Q (new_AGEMA_signal_9021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_9024), .Q (new_AGEMA_signal_9025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_9028), .Q (new_AGEMA_signal_9029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_9032), .Q (new_AGEMA_signal_9033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_9036), .Q (new_AGEMA_signal_9037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_9040), .Q (new_AGEMA_signal_9041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_9044), .Q (new_AGEMA_signal_9045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_9048), .Q (new_AGEMA_signal_9049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_9052), .Q (new_AGEMA_signal_9053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_9056), .Q (new_AGEMA_signal_9057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_9060), .Q (new_AGEMA_signal_9061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_9064), .Q (new_AGEMA_signal_9065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_9068), .Q (new_AGEMA_signal_9069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_9072), .Q (new_AGEMA_signal_9073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_9076), .Q (new_AGEMA_signal_9077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_9080), .Q (new_AGEMA_signal_9081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_9084), .Q (new_AGEMA_signal_9085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_9088), .Q (new_AGEMA_signal_9089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_9092), .Q (new_AGEMA_signal_9093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_9096), .Q (new_AGEMA_signal_9097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_9100), .Q (new_AGEMA_signal_9101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_9104), .Q (new_AGEMA_signal_9105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_9108), .Q (new_AGEMA_signal_9109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_9112), .Q (new_AGEMA_signal_9113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_9116), .Q (new_AGEMA_signal_9117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_9120), .Q (new_AGEMA_signal_9121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_9124), .Q (new_AGEMA_signal_9125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_9128), .Q (new_AGEMA_signal_9129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_9132), .Q (new_AGEMA_signal_9133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_9136), .Q (new_AGEMA_signal_9137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_9140), .Q (new_AGEMA_signal_9141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_9144), .Q (new_AGEMA_signal_9145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_9148), .Q (new_AGEMA_signal_9149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_9152), .Q (new_AGEMA_signal_9153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_9156), .Q (new_AGEMA_signal_9157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_9160), .Q (new_AGEMA_signal_9161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_9164), .Q (new_AGEMA_signal_9165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_9168), .Q (new_AGEMA_signal_9169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_9172), .Q (new_AGEMA_signal_9173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_9176), .Q (new_AGEMA_signal_9177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_9180), .Q (new_AGEMA_signal_9181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_9184), .Q (new_AGEMA_signal_9185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_9188), .Q (new_AGEMA_signal_9189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_9192), .Q (new_AGEMA_signal_9193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_9196), .Q (new_AGEMA_signal_9197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_9200), .Q (new_AGEMA_signal_9201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_9204), .Q (new_AGEMA_signal_9205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_9208), .Q (new_AGEMA_signal_9209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_9212), .Q (new_AGEMA_signal_9213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_9216), .Q (new_AGEMA_signal_9217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_9220), .Q (new_AGEMA_signal_9221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_9224), .Q (new_AGEMA_signal_9225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_9228), .Q (new_AGEMA_signal_9229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_9232), .Q (new_AGEMA_signal_9233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_9236), .Q (new_AGEMA_signal_9237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_9240), .Q (new_AGEMA_signal_9241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_9244), .Q (new_AGEMA_signal_9245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_9248), .Q (new_AGEMA_signal_9249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_9252), .Q (new_AGEMA_signal_9253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_9256), .Q (new_AGEMA_signal_9257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_9260), .Q (new_AGEMA_signal_9261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_9264), .Q (new_AGEMA_signal_9265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_9268), .Q (new_AGEMA_signal_9269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_9272), .Q (new_AGEMA_signal_9273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_9276), .Q (new_AGEMA_signal_9277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_9280), .Q (new_AGEMA_signal_9281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_9284), .Q (new_AGEMA_signal_9285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_9288), .Q (new_AGEMA_signal_9289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_9292), .Q (new_AGEMA_signal_9293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_9296), .Q (new_AGEMA_signal_9297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_9300), .Q (new_AGEMA_signal_9301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_9304), .Q (new_AGEMA_signal_9305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_9308), .Q (new_AGEMA_signal_9309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_9312), .Q (new_AGEMA_signal_9313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_9316), .Q (new_AGEMA_signal_9317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_9320), .Q (new_AGEMA_signal_9321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_9324), .Q (new_AGEMA_signal_9325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_9328), .Q (new_AGEMA_signal_9329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_9332), .Q (new_AGEMA_signal_9333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_9336), .Q (new_AGEMA_signal_9337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_9340), .Q (new_AGEMA_signal_9341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_9344), .Q (new_AGEMA_signal_9345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_9348), .Q (new_AGEMA_signal_9349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_9352), .Q (new_AGEMA_signal_9353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_9356), .Q (new_AGEMA_signal_9357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_9360), .Q (new_AGEMA_signal_9361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_9364), .Q (new_AGEMA_signal_9365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_9368), .Q (new_AGEMA_signal_9369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_9372), .Q (new_AGEMA_signal_9373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_9376), .Q (new_AGEMA_signal_9377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_9380), .Q (new_AGEMA_signal_9381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_9384), .Q (new_AGEMA_signal_9385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_9388), .Q (new_AGEMA_signal_9389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_9392), .Q (new_AGEMA_signal_9393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_9396), .Q (new_AGEMA_signal_9397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_9400), .Q (new_AGEMA_signal_9401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_9404), .Q (new_AGEMA_signal_9405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_9408), .Q (new_AGEMA_signal_9409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_9412), .Q (new_AGEMA_signal_9413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_9416), .Q (new_AGEMA_signal_9417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_9420), .Q (new_AGEMA_signal_9421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_9424), .Q (new_AGEMA_signal_9425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_9428), .Q (new_AGEMA_signal_9429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_9432), .Q (new_AGEMA_signal_9433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_9436), .Q (new_AGEMA_signal_9437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_9440), .Q (new_AGEMA_signal_9441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_9444), .Q (new_AGEMA_signal_9445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_9448), .Q (new_AGEMA_signal_9449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_9452), .Q (new_AGEMA_signal_9453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_9456), .Q (new_AGEMA_signal_9457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_9460), .Q (new_AGEMA_signal_9461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_9464), .Q (new_AGEMA_signal_9465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_9468), .Q (new_AGEMA_signal_9469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_9472), .Q (new_AGEMA_signal_9473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_9476), .Q (new_AGEMA_signal_9477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_9480), .Q (new_AGEMA_signal_9481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_9484), .Q (new_AGEMA_signal_9485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_9488), .Q (new_AGEMA_signal_9489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_9492), .Q (new_AGEMA_signal_9493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_9496), .Q (new_AGEMA_signal_9497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_9500), .Q (new_AGEMA_signal_9501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_9504), .Q (new_AGEMA_signal_9505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_9508), .Q (new_AGEMA_signal_9509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_9512), .Q (new_AGEMA_signal_9513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_9516), .Q (new_AGEMA_signal_9517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_9520), .Q (new_AGEMA_signal_9521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_9524), .Q (new_AGEMA_signal_9525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_9528), .Q (new_AGEMA_signal_9529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_9532), .Q (new_AGEMA_signal_9533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_9536), .Q (new_AGEMA_signal_9537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_9540), .Q (new_AGEMA_signal_9541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_9544), .Q (new_AGEMA_signal_9545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_9548), .Q (new_AGEMA_signal_9549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_9552), .Q (new_AGEMA_signal_9553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_9556), .Q (new_AGEMA_signal_9557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_9560), .Q (new_AGEMA_signal_9561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_9564), .Q (new_AGEMA_signal_9565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_9568), .Q (new_AGEMA_signal_9569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_9572), .Q (new_AGEMA_signal_9573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_9576), .Q (new_AGEMA_signal_9577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_9580), .Q (new_AGEMA_signal_9581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_9584), .Q (new_AGEMA_signal_9585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_9588), .Q (new_AGEMA_signal_9589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_9592), .Q (new_AGEMA_signal_9593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_9596), .Q (new_AGEMA_signal_9597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_9600), .Q (new_AGEMA_signal_9601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_9604), .Q (new_AGEMA_signal_9605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_9608), .Q (new_AGEMA_signal_9609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_9612), .Q (new_AGEMA_signal_9613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_9616), .Q (new_AGEMA_signal_9617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_9620), .Q (new_AGEMA_signal_9621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_9624), .Q (new_AGEMA_signal_9625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_9628), .Q (new_AGEMA_signal_9629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_9632), .Q (new_AGEMA_signal_9633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_9636), .Q (new_AGEMA_signal_9637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_9640), .Q (new_AGEMA_signal_9641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_9644), .Q (new_AGEMA_signal_9645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_9648), .Q (new_AGEMA_signal_9649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_9652), .Q (new_AGEMA_signal_9653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_9656), .Q (new_AGEMA_signal_9657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_9660), .Q (new_AGEMA_signal_9661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_9664), .Q (new_AGEMA_signal_9665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_9668), .Q (new_AGEMA_signal_9669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_9672), .Q (new_AGEMA_signal_9673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_9676), .Q (new_AGEMA_signal_9677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_9680), .Q (new_AGEMA_signal_9681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_9684), .Q (new_AGEMA_signal_9685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_9688), .Q (new_AGEMA_signal_9689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_9692), .Q (new_AGEMA_signal_9693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_9696), .Q (new_AGEMA_signal_9697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_9700), .Q (new_AGEMA_signal_9701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_9704), .Q (new_AGEMA_signal_9705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_9708), .Q (new_AGEMA_signal_9709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_9712), .Q (new_AGEMA_signal_9713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_9716), .Q (new_AGEMA_signal_9717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_9720), .Q (new_AGEMA_signal_9721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_9724), .Q (new_AGEMA_signal_9725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_9728), .Q (new_AGEMA_signal_9729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_9732), .Q (new_AGEMA_signal_9733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_9736), .Q (new_AGEMA_signal_9737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_9740), .Q (new_AGEMA_signal_9741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_9744), .Q (new_AGEMA_signal_9745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_9748), .Q (new_AGEMA_signal_9749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_9752), .Q (new_AGEMA_signal_9753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_9756), .Q (new_AGEMA_signal_9757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_9760), .Q (new_AGEMA_signal_9761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_9764), .Q (new_AGEMA_signal_9765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_9768), .Q (new_AGEMA_signal_9769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_9772), .Q (new_AGEMA_signal_9773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_9776), .Q (new_AGEMA_signal_9777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_9780), .Q (new_AGEMA_signal_9781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_9784), .Q (new_AGEMA_signal_9785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_9788), .Q (new_AGEMA_signal_9789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_9792), .Q (new_AGEMA_signal_9793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_9796), .Q (new_AGEMA_signal_9797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_9800), .Q (new_AGEMA_signal_9801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_9804), .Q (new_AGEMA_signal_9805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_9808), .Q (new_AGEMA_signal_9809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_9812), .Q (new_AGEMA_signal_9813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_9816), .Q (new_AGEMA_signal_9817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_9820), .Q (new_AGEMA_signal_9821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_9824), .Q (new_AGEMA_signal_9825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_9828), .Q (new_AGEMA_signal_9829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_9832), .Q (new_AGEMA_signal_9833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_9836), .Q (new_AGEMA_signal_9837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_9840), .Q (new_AGEMA_signal_9841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_9844), .Q (new_AGEMA_signal_9845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_9848), .Q (new_AGEMA_signal_9849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_9852), .Q (new_AGEMA_signal_9853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_9856), .Q (new_AGEMA_signal_9857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_9860), .Q (new_AGEMA_signal_9861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_9864), .Q (new_AGEMA_signal_9865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_9868), .Q (new_AGEMA_signal_9869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_9872), .Q (new_AGEMA_signal_9873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_9876), .Q (new_AGEMA_signal_9877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_9880), .Q (new_AGEMA_signal_9881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_9884), .Q (new_AGEMA_signal_9885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_9888), .Q (new_AGEMA_signal_9889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_9892), .Q (new_AGEMA_signal_9893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_9896), .Q (new_AGEMA_signal_9897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_9900), .Q (new_AGEMA_signal_9901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_9904), .Q (new_AGEMA_signal_9905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_9908), .Q (new_AGEMA_signal_9909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_9912), .Q (new_AGEMA_signal_9913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_9916), .Q (new_AGEMA_signal_9917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_9920), .Q (new_AGEMA_signal_9921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_9924), .Q (new_AGEMA_signal_9925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_9928), .Q (new_AGEMA_signal_9929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4896 ( .C (clk), .D (new_AGEMA_signal_9932), .Q (new_AGEMA_signal_9933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_9936), .Q (new_AGEMA_signal_9937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_9940), .Q (new_AGEMA_signal_9941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4908 ( .C (clk), .D (new_AGEMA_signal_9944), .Q (new_AGEMA_signal_9945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_9948), .Q (new_AGEMA_signal_9949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_9952), .Q (new_AGEMA_signal_9953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4920 ( .C (clk), .D (new_AGEMA_signal_9956), .Q (new_AGEMA_signal_9957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_9960), .Q (new_AGEMA_signal_9961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_9964), .Q (new_AGEMA_signal_9965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_9968), .Q (new_AGEMA_signal_9969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_9972), .Q (new_AGEMA_signal_9973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_9976), .Q (new_AGEMA_signal_9977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_9980), .Q (new_AGEMA_signal_9981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_9984), .Q (new_AGEMA_signal_9985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_9988), .Q (new_AGEMA_signal_9989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_9992), .Q (new_AGEMA_signal_9993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_9996), .Q (new_AGEMA_signal_9997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_10000), .Q (new_AGEMA_signal_10001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_10004), .Q (new_AGEMA_signal_10005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_10008), .Q (new_AGEMA_signal_10009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_10012), .Q (new_AGEMA_signal_10013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_10016), .Q (new_AGEMA_signal_10017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_10020), .Q (new_AGEMA_signal_10021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_10024), .Q (new_AGEMA_signal_10025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_10028), .Q (new_AGEMA_signal_10029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_10032), .Q (new_AGEMA_signal_10033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_10036), .Q (new_AGEMA_signal_10037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_10040), .Q (new_AGEMA_signal_10041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_10044), .Q (new_AGEMA_signal_10045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_10048), .Q (new_AGEMA_signal_10049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_10052), .Q (new_AGEMA_signal_10053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_10056), .Q (new_AGEMA_signal_10057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_10060), .Q (new_AGEMA_signal_10061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_10064), .Q (new_AGEMA_signal_10065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_10068), .Q (new_AGEMA_signal_10069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_10072), .Q (new_AGEMA_signal_10073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_10076), .Q (new_AGEMA_signal_10077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_10080), .Q (new_AGEMA_signal_10081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_10084), .Q (new_AGEMA_signal_10085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_10088), .Q (new_AGEMA_signal_10089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_10092), .Q (new_AGEMA_signal_10093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_10096), .Q (new_AGEMA_signal_10097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_10100), .Q (new_AGEMA_signal_10101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_10104), .Q (new_AGEMA_signal_10105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_10108), .Q (new_AGEMA_signal_10109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_10112), .Q (new_AGEMA_signal_10113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_10116), .Q (new_AGEMA_signal_10117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_10120), .Q (new_AGEMA_signal_10121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_10124), .Q (new_AGEMA_signal_10125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_10128), .Q (new_AGEMA_signal_10129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_10132), .Q (new_AGEMA_signal_10133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_10136), .Q (new_AGEMA_signal_10137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_10140), .Q (new_AGEMA_signal_10141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_10144), .Q (new_AGEMA_signal_10145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_10148), .Q (new_AGEMA_signal_10149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_10152), .Q (new_AGEMA_signal_10153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_10156), .Q (new_AGEMA_signal_10157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_10160), .Q (new_AGEMA_signal_10161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_10164), .Q (new_AGEMA_signal_10165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_10168), .Q (new_AGEMA_signal_10169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_10172), .Q (new_AGEMA_signal_10173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_10176), .Q (new_AGEMA_signal_10177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_10180), .Q (new_AGEMA_signal_10181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_10184), .Q (new_AGEMA_signal_10185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_10188), .Q (new_AGEMA_signal_10189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_10192), .Q (new_AGEMA_signal_10193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_10196), .Q (new_AGEMA_signal_10197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_10200), .Q (new_AGEMA_signal_10201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_10204), .Q (new_AGEMA_signal_10205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_10208), .Q (new_AGEMA_signal_10209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_10212), .Q (new_AGEMA_signal_10213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_10216), .Q (new_AGEMA_signal_10217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_10220), .Q (new_AGEMA_signal_10221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_10224), .Q (new_AGEMA_signal_10225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_10228), .Q (new_AGEMA_signal_10229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_10232), .Q (new_AGEMA_signal_10233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_10236), .Q (new_AGEMA_signal_10237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_10240), .Q (new_AGEMA_signal_10241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_10244), .Q (new_AGEMA_signal_10245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_10248), .Q (new_AGEMA_signal_10249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_10252), .Q (new_AGEMA_signal_10253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_10256), .Q (new_AGEMA_signal_10257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_10260), .Q (new_AGEMA_signal_10261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_10264), .Q (new_AGEMA_signal_10265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_10268), .Q (new_AGEMA_signal_10269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_10272), .Q (new_AGEMA_signal_10273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_10276), .Q (new_AGEMA_signal_10277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_10280), .Q (new_AGEMA_signal_10281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_10284), .Q (new_AGEMA_signal_10285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_10288), .Q (new_AGEMA_signal_10289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_10292), .Q (new_AGEMA_signal_10293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_10296), .Q (new_AGEMA_signal_10297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_10300), .Q (new_AGEMA_signal_10301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_10304), .Q (new_AGEMA_signal_10305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_10308), .Q (new_AGEMA_signal_10309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_10312), .Q (new_AGEMA_signal_10313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_10316), .Q (new_AGEMA_signal_10317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_10320), .Q (new_AGEMA_signal_10321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_10324), .Q (new_AGEMA_signal_10325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_10328), .Q (new_AGEMA_signal_10329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_10332), .Q (new_AGEMA_signal_10333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_10336), .Q (new_AGEMA_signal_10337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_10340), .Q (new_AGEMA_signal_10341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_10344), .Q (new_AGEMA_signal_10345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_10348), .Q (new_AGEMA_signal_10349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_10352), .Q (new_AGEMA_signal_10353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_10356), .Q (new_AGEMA_signal_10357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_10360), .Q (new_AGEMA_signal_10361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_10364), .Q (new_AGEMA_signal_10365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_10368), .Q (new_AGEMA_signal_10369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_10372), .Q (new_AGEMA_signal_10373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_10376), .Q (new_AGEMA_signal_10377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_10380), .Q (new_AGEMA_signal_10381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_10384), .Q (new_AGEMA_signal_10385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_10388), .Q (new_AGEMA_signal_10389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_10392), .Q (new_AGEMA_signal_10393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_10396), .Q (new_AGEMA_signal_10397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_10400), .Q (new_AGEMA_signal_10401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_10404), .Q (new_AGEMA_signal_10405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_10408), .Q (new_AGEMA_signal_10409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_10412), .Q (new_AGEMA_signal_10413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_10416), .Q (new_AGEMA_signal_10417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_10420), .Q (new_AGEMA_signal_10421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_10424), .Q (new_AGEMA_signal_10425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_10428), .Q (new_AGEMA_signal_10429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_10432), .Q (new_AGEMA_signal_10433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_10436), .Q (new_AGEMA_signal_10437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_10440), .Q (new_AGEMA_signal_10441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_10444), .Q (new_AGEMA_signal_10445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_10448), .Q (new_AGEMA_signal_10449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_10452), .Q (new_AGEMA_signal_10453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_10456), .Q (new_AGEMA_signal_10457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_10460), .Q (new_AGEMA_signal_10461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_10464), .Q (new_AGEMA_signal_10465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_10468), .Q (new_AGEMA_signal_10469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_10472), .Q (new_AGEMA_signal_10473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_10476), .Q (new_AGEMA_signal_10477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_10480), .Q (new_AGEMA_signal_10481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_10484), .Q (new_AGEMA_signal_10485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_10488), .Q (new_AGEMA_signal_10489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_10492), .Q (new_AGEMA_signal_10493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_10496), .Q (new_AGEMA_signal_10497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_10500), .Q (new_AGEMA_signal_10501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_10504), .Q (new_AGEMA_signal_10505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_10508), .Q (new_AGEMA_signal_10509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_10512), .Q (new_AGEMA_signal_10513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_10516), .Q (new_AGEMA_signal_10517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_10520), .Q (new_AGEMA_signal_10521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_10524), .Q (new_AGEMA_signal_10525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_10528), .Q (new_AGEMA_signal_10529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_10532), .Q (new_AGEMA_signal_10533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_10536), .Q (new_AGEMA_signal_10537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_10540), .Q (new_AGEMA_signal_10541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_10544), .Q (new_AGEMA_signal_10545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_10548), .Q (new_AGEMA_signal_10549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_10552), .Q (new_AGEMA_signal_10553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_10556), .Q (new_AGEMA_signal_10557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_10560), .Q (new_AGEMA_signal_10561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_10564), .Q (new_AGEMA_signal_10565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_10568), .Q (new_AGEMA_signal_10569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_10572), .Q (new_AGEMA_signal_10573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_10576), .Q (new_AGEMA_signal_10577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_10580), .Q (new_AGEMA_signal_10581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_10584), .Q (new_AGEMA_signal_10585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_10588), .Q (new_AGEMA_signal_10589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_10592), .Q (new_AGEMA_signal_10593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_10596), .Q (new_AGEMA_signal_10597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_10600), .Q (new_AGEMA_signal_10601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_10604), .Q (new_AGEMA_signal_10605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_10608), .Q (new_AGEMA_signal_10609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_10612), .Q (new_AGEMA_signal_10613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_10616), .Q (new_AGEMA_signal_10617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_10620), .Q (new_AGEMA_signal_10621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_10624), .Q (new_AGEMA_signal_10625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_10628), .Q (new_AGEMA_signal_10629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_10632), .Q (new_AGEMA_signal_10633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_10636), .Q (new_AGEMA_signal_10637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_10640), .Q (new_AGEMA_signal_10641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_10644), .Q (new_AGEMA_signal_10645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_10648), .Q (new_AGEMA_signal_10649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_10652), .Q (new_AGEMA_signal_10653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_10656), .Q (new_AGEMA_signal_10657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_10660), .Q (new_AGEMA_signal_10661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_10664), .Q (new_AGEMA_signal_10665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_10668), .Q (new_AGEMA_signal_10669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_10672), .Q (new_AGEMA_signal_10673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_10676), .Q (new_AGEMA_signal_10677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_10680), .Q (new_AGEMA_signal_10681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_10684), .Q (new_AGEMA_signal_10685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_10688), .Q (new_AGEMA_signal_10689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_10692), .Q (new_AGEMA_signal_10693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_10696), .Q (new_AGEMA_signal_10697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_10700), .Q (new_AGEMA_signal_10701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_10704), .Q (new_AGEMA_signal_10705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_10708), .Q (new_AGEMA_signal_10709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_10712), .Q (new_AGEMA_signal_10713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_10716), .Q (new_AGEMA_signal_10717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_10720), .Q (new_AGEMA_signal_10721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_10724), .Q (new_AGEMA_signal_10725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_10728), .Q (new_AGEMA_signal_10729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_10732), .Q (new_AGEMA_signal_10733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_10736), .Q (new_AGEMA_signal_10737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_10740), .Q (new_AGEMA_signal_10741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_10744), .Q (new_AGEMA_signal_10745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_10748), .Q (new_AGEMA_signal_10749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_10752), .Q (new_AGEMA_signal_10753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_10756), .Q (new_AGEMA_signal_10757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_10760), .Q (new_AGEMA_signal_10761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_10764), .Q (new_AGEMA_signal_10765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_10768), .Q (new_AGEMA_signal_10769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_10772), .Q (new_AGEMA_signal_10773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_10776), .Q (new_AGEMA_signal_10777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_10780), .Q (new_AGEMA_signal_10781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_10784), .Q (new_AGEMA_signal_10785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_10788), .Q (new_AGEMA_signal_10789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_10792), .Q (new_AGEMA_signal_10793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5760 ( .C (clk), .D (new_AGEMA_signal_10796), .Q (new_AGEMA_signal_10797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_10800), .Q (new_AGEMA_signal_10801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_10804), .Q (new_AGEMA_signal_10805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_10808), .Q (new_AGEMA_signal_10809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_10812), .Q (new_AGEMA_signal_10813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_10816), .Q (new_AGEMA_signal_10817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_10820), .Q (new_AGEMA_signal_10821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_10824), .Q (new_AGEMA_signal_10825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_10828), .Q (new_AGEMA_signal_10829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_10832), .Q (new_AGEMA_signal_10833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_10836), .Q (new_AGEMA_signal_10837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_10840), .Q (new_AGEMA_signal_10841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_10844), .Q (new_AGEMA_signal_10845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_10848), .Q (new_AGEMA_signal_10849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_10852), .Q (new_AGEMA_signal_10853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_10856), .Q (new_AGEMA_signal_10857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_10860), .Q (new_AGEMA_signal_10861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_10864), .Q (new_AGEMA_signal_10865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_10868), .Q (new_AGEMA_signal_10869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_10872), .Q (new_AGEMA_signal_10873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_10876), .Q (new_AGEMA_signal_10877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_10880), .Q (new_AGEMA_signal_10881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_10884), .Q (new_AGEMA_signal_10885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_10888), .Q (new_AGEMA_signal_10889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_10892), .Q (new_AGEMA_signal_10893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_10896), .Q (new_AGEMA_signal_10897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_10900), .Q (new_AGEMA_signal_10901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5868 ( .C (clk), .D (new_AGEMA_signal_10904), .Q (new_AGEMA_signal_10905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_10908), .Q (new_AGEMA_signal_10909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_10912), .Q (new_AGEMA_signal_10913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_10916), .Q (new_AGEMA_signal_10917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_10920), .Q (new_AGEMA_signal_10921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_10924), .Q (new_AGEMA_signal_10925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_10928), .Q (new_AGEMA_signal_10929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_10932), .Q (new_AGEMA_signal_10933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_10936), .Q (new_AGEMA_signal_10937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_10940), .Q (new_AGEMA_signal_10941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_10944), .Q (new_AGEMA_signal_10945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_10948), .Q (new_AGEMA_signal_10949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_10952), .Q (new_AGEMA_signal_10953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_10956), .Q (new_AGEMA_signal_10957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_10960), .Q (new_AGEMA_signal_10961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_10964), .Q (new_AGEMA_signal_10965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_10968), .Q (new_AGEMA_signal_10969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_10972), .Q (new_AGEMA_signal_10973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_10976), .Q (new_AGEMA_signal_10977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_10980), .Q (new_AGEMA_signal_10981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_10984), .Q (new_AGEMA_signal_10985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_10988), .Q (new_AGEMA_signal_10989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_10992), .Q (new_AGEMA_signal_10993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_10996), .Q (new_AGEMA_signal_10997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_11000), .Q (new_AGEMA_signal_11001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_11004), .Q (new_AGEMA_signal_11005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_11008), .Q (new_AGEMA_signal_11009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5976 ( .C (clk), .D (new_AGEMA_signal_11012), .Q (new_AGEMA_signal_11013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_11016), .Q (new_AGEMA_signal_11017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_11020), .Q (new_AGEMA_signal_11021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_11024), .Q (new_AGEMA_signal_11025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_11028), .Q (new_AGEMA_signal_11029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_11032), .Q (new_AGEMA_signal_11033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_11036), .Q (new_AGEMA_signal_11037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_11040), .Q (new_AGEMA_signal_11041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_11044), .Q (new_AGEMA_signal_11045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_11048), .Q (new_AGEMA_signal_11049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_11052), .Q (new_AGEMA_signal_11053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_11056), .Q (new_AGEMA_signal_11057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_11060), .Q (new_AGEMA_signal_11061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_11064), .Q (new_AGEMA_signal_11065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_11068), .Q (new_AGEMA_signal_11069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_11072), .Q (new_AGEMA_signal_11073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_11076), .Q (new_AGEMA_signal_11077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_11080), .Q (new_AGEMA_signal_11081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_11084), .Q (new_AGEMA_signal_11085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6052 ( .C (clk), .D (new_AGEMA_signal_11088), .Q (new_AGEMA_signal_11089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6056 ( .C (clk), .D (new_AGEMA_signal_11092), .Q (new_AGEMA_signal_11093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6060 ( .C (clk), .D (new_AGEMA_signal_11096), .Q (new_AGEMA_signal_11097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6064 ( .C (clk), .D (new_AGEMA_signal_11100), .Q (new_AGEMA_signal_11101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6068 ( .C (clk), .D (new_AGEMA_signal_11104), .Q (new_AGEMA_signal_11105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6072 ( .C (clk), .D (new_AGEMA_signal_11108), .Q (new_AGEMA_signal_11109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6076 ( .C (clk), .D (new_AGEMA_signal_11112), .Q (new_AGEMA_signal_11113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6080 ( .C (clk), .D (new_AGEMA_signal_11116), .Q (new_AGEMA_signal_11117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6084 ( .C (clk), .D (new_AGEMA_signal_11120), .Q (new_AGEMA_signal_11121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6088 ( .C (clk), .D (new_AGEMA_signal_11124), .Q (new_AGEMA_signal_11125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6092 ( .C (clk), .D (new_AGEMA_signal_11128), .Q (new_AGEMA_signal_11129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6096 ( .C (clk), .D (new_AGEMA_signal_11132), .Q (new_AGEMA_signal_11133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6100 ( .C (clk), .D (new_AGEMA_signal_11136), .Q (new_AGEMA_signal_11137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6104 ( .C (clk), .D (new_AGEMA_signal_11140), .Q (new_AGEMA_signal_11141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6108 ( .C (clk), .D (new_AGEMA_signal_11144), .Q (new_AGEMA_signal_11145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6112 ( .C (clk), .D (new_AGEMA_signal_11148), .Q (new_AGEMA_signal_11149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6116 ( .C (clk), .D (new_AGEMA_signal_11152), .Q (new_AGEMA_signal_11153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6120 ( .C (clk), .D (new_AGEMA_signal_11156), .Q (new_AGEMA_signal_11157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6124 ( .C (clk), .D (new_AGEMA_signal_11160), .Q (new_AGEMA_signal_11161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6128 ( .C (clk), .D (new_AGEMA_signal_11164), .Q (new_AGEMA_signal_11165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6132 ( .C (clk), .D (new_AGEMA_signal_11168), .Q (new_AGEMA_signal_11169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6136 ( .C (clk), .D (new_AGEMA_signal_11172), .Q (new_AGEMA_signal_11173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6140 ( .C (clk), .D (new_AGEMA_signal_11176), .Q (new_AGEMA_signal_11177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6144 ( .C (clk), .D (new_AGEMA_signal_11180), .Q (new_AGEMA_signal_11181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6148 ( .C (clk), .D (new_AGEMA_signal_11184), .Q (new_AGEMA_signal_11185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6152 ( .C (clk), .D (new_AGEMA_signal_11188), .Q (new_AGEMA_signal_11189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6156 ( .C (clk), .D (new_AGEMA_signal_11192), .Q (new_AGEMA_signal_11193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6160 ( .C (clk), .D (new_AGEMA_signal_11196), .Q (new_AGEMA_signal_11197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6164 ( .C (clk), .D (new_AGEMA_signal_11200), .Q (new_AGEMA_signal_11201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6168 ( .C (clk), .D (new_AGEMA_signal_11204), .Q (new_AGEMA_signal_11205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6172 ( .C (clk), .D (new_AGEMA_signal_11208), .Q (new_AGEMA_signal_11209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6176 ( .C (clk), .D (new_AGEMA_signal_11212), .Q (new_AGEMA_signal_11213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6180 ( .C (clk), .D (new_AGEMA_signal_11216), .Q (new_AGEMA_signal_11217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6184 ( .C (clk), .D (new_AGEMA_signal_11220), .Q (new_AGEMA_signal_11221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6188 ( .C (clk), .D (new_AGEMA_signal_11224), .Q (new_AGEMA_signal_11225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6192 ( .C (clk), .D (new_AGEMA_signal_11228), .Q (new_AGEMA_signal_11229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6196 ( .C (clk), .D (new_AGEMA_signal_11232), .Q (new_AGEMA_signal_11233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6200 ( .C (clk), .D (new_AGEMA_signal_11236), .Q (new_AGEMA_signal_11237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6204 ( .C (clk), .D (new_AGEMA_signal_11240), .Q (new_AGEMA_signal_11241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6208 ( .C (clk), .D (new_AGEMA_signal_11244), .Q (new_AGEMA_signal_11245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6212 ( .C (clk), .D (new_AGEMA_signal_11248), .Q (new_AGEMA_signal_11249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6216 ( .C (clk), .D (new_AGEMA_signal_11252), .Q (new_AGEMA_signal_11253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6220 ( .C (clk), .D (new_AGEMA_signal_11256), .Q (new_AGEMA_signal_11257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6224 ( .C (clk), .D (new_AGEMA_signal_11260), .Q (new_AGEMA_signal_11261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6228 ( .C (clk), .D (new_AGEMA_signal_11264), .Q (new_AGEMA_signal_11265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6232 ( .C (clk), .D (new_AGEMA_signal_11268), .Q (new_AGEMA_signal_11269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6236 ( .C (clk), .D (new_AGEMA_signal_11272), .Q (new_AGEMA_signal_11273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6240 ( .C (clk), .D (new_AGEMA_signal_11276), .Q (new_AGEMA_signal_11277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6244 ( .C (clk), .D (new_AGEMA_signal_11280), .Q (new_AGEMA_signal_11281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6248 ( .C (clk), .D (new_AGEMA_signal_11284), .Q (new_AGEMA_signal_11285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6252 ( .C (clk), .D (new_AGEMA_signal_11288), .Q (new_AGEMA_signal_11289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6256 ( .C (clk), .D (new_AGEMA_signal_11292), .Q (new_AGEMA_signal_11293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6260 ( .C (clk), .D (new_AGEMA_signal_11296), .Q (new_AGEMA_signal_11297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6264 ( .C (clk), .D (new_AGEMA_signal_11300), .Q (new_AGEMA_signal_11301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6268 ( .C (clk), .D (new_AGEMA_signal_11304), .Q (new_AGEMA_signal_11305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6272 ( .C (clk), .D (new_AGEMA_signal_11308), .Q (new_AGEMA_signal_11309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6276 ( .C (clk), .D (new_AGEMA_signal_11312), .Q (new_AGEMA_signal_11313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6280 ( .C (clk), .D (new_AGEMA_signal_11316), .Q (new_AGEMA_signal_11317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6284 ( .C (clk), .D (new_AGEMA_signal_11320), .Q (new_AGEMA_signal_11321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6288 ( .C (clk), .D (new_AGEMA_signal_11324), .Q (new_AGEMA_signal_11325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6292 ( .C (clk), .D (new_AGEMA_signal_11328), .Q (new_AGEMA_signal_11329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6296 ( .C (clk), .D (new_AGEMA_signal_11332), .Q (new_AGEMA_signal_11333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6300 ( .C (clk), .D (new_AGEMA_signal_11336), .Q (new_AGEMA_signal_11337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6304 ( .C (clk), .D (new_AGEMA_signal_11340), .Q (new_AGEMA_signal_11341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6308 ( .C (clk), .D (new_AGEMA_signal_11344), .Q (new_AGEMA_signal_11345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6312 ( .C (clk), .D (new_AGEMA_signal_11348), .Q (new_AGEMA_signal_11349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6316 ( .C (clk), .D (new_AGEMA_signal_11352), .Q (new_AGEMA_signal_11353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6320 ( .C (clk), .D (new_AGEMA_signal_11356), .Q (new_AGEMA_signal_11357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6324 ( .C (clk), .D (new_AGEMA_signal_11360), .Q (new_AGEMA_signal_11361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6328 ( .C (clk), .D (new_AGEMA_signal_11364), .Q (new_AGEMA_signal_11365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6332 ( .C (clk), .D (new_AGEMA_signal_11368), .Q (new_AGEMA_signal_11369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6336 ( .C (clk), .D (new_AGEMA_signal_11372), .Q (new_AGEMA_signal_11373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6340 ( .C (clk), .D (new_AGEMA_signal_11376), .Q (new_AGEMA_signal_11377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6344 ( .C (clk), .D (new_AGEMA_signal_11380), .Q (new_AGEMA_signal_11381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6348 ( .C (clk), .D (new_AGEMA_signal_11384), .Q (new_AGEMA_signal_11385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6352 ( .C (clk), .D (new_AGEMA_signal_11388), .Q (new_AGEMA_signal_11389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6356 ( .C (clk), .D (new_AGEMA_signal_11392), .Q (new_AGEMA_signal_11393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6360 ( .C (clk), .D (new_AGEMA_signal_11396), .Q (new_AGEMA_signal_11397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6364 ( .C (clk), .D (new_AGEMA_signal_11400), .Q (new_AGEMA_signal_11401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6368 ( .C (clk), .D (new_AGEMA_signal_11404), .Q (new_AGEMA_signal_11405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6372 ( .C (clk), .D (new_AGEMA_signal_11408), .Q (new_AGEMA_signal_11409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6376 ( .C (clk), .D (new_AGEMA_signal_11412), .Q (new_AGEMA_signal_11413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6380 ( .C (clk), .D (new_AGEMA_signal_11416), .Q (new_AGEMA_signal_11417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6384 ( .C (clk), .D (new_AGEMA_signal_11420), .Q (new_AGEMA_signal_11421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6388 ( .C (clk), .D (new_AGEMA_signal_11424), .Q (new_AGEMA_signal_11425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6392 ( .C (clk), .D (new_AGEMA_signal_11428), .Q (new_AGEMA_signal_11429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6396 ( .C (clk), .D (new_AGEMA_signal_11432), .Q (new_AGEMA_signal_11433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6400 ( .C (clk), .D (new_AGEMA_signal_11436), .Q (new_AGEMA_signal_11437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6404 ( .C (clk), .D (new_AGEMA_signal_11440), .Q (new_AGEMA_signal_11441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6408 ( .C (clk), .D (new_AGEMA_signal_11444), .Q (new_AGEMA_signal_11445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6412 ( .C (clk), .D (new_AGEMA_signal_11448), .Q (new_AGEMA_signal_11449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6416 ( .C (clk), .D (new_AGEMA_signal_11452), .Q (new_AGEMA_signal_11453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6420 ( .C (clk), .D (new_AGEMA_signal_11456), .Q (new_AGEMA_signal_11457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6424 ( .C (clk), .D (new_AGEMA_signal_11460), .Q (new_AGEMA_signal_11461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6428 ( .C (clk), .D (new_AGEMA_signal_11464), .Q (new_AGEMA_signal_11465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6432 ( .C (clk), .D (new_AGEMA_signal_11468), .Q (new_AGEMA_signal_11469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6436 ( .C (clk), .D (new_AGEMA_signal_11472), .Q (new_AGEMA_signal_11473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6440 ( .C (clk), .D (new_AGEMA_signal_11476), .Q (new_AGEMA_signal_11477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6444 ( .C (clk), .D (new_AGEMA_signal_11480), .Q (new_AGEMA_signal_11481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6448 ( .C (clk), .D (new_AGEMA_signal_11484), .Q (new_AGEMA_signal_11485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6452 ( .C (clk), .D (new_AGEMA_signal_11488), .Q (new_AGEMA_signal_11489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6456 ( .C (clk), .D (new_AGEMA_signal_11492), .Q (new_AGEMA_signal_11493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6460 ( .C (clk), .D (new_AGEMA_signal_11496), .Q (new_AGEMA_signal_11497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6464 ( .C (clk), .D (new_AGEMA_signal_11500), .Q (new_AGEMA_signal_11501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6468 ( .C (clk), .D (new_AGEMA_signal_11504), .Q (new_AGEMA_signal_11505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6472 ( .C (clk), .D (new_AGEMA_signal_11508), .Q (new_AGEMA_signal_11509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6476 ( .C (clk), .D (new_AGEMA_signal_11512), .Q (new_AGEMA_signal_11513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6480 ( .C (clk), .D (new_AGEMA_signal_11516), .Q (new_AGEMA_signal_11517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6484 ( .C (clk), .D (new_AGEMA_signal_11520), .Q (new_AGEMA_signal_11521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6488 ( .C (clk), .D (new_AGEMA_signal_11524), .Q (new_AGEMA_signal_11525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6492 ( .C (clk), .D (new_AGEMA_signal_11528), .Q (new_AGEMA_signal_11529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6496 ( .C (clk), .D (new_AGEMA_signal_11532), .Q (new_AGEMA_signal_11533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6500 ( .C (clk), .D (new_AGEMA_signal_11536), .Q (new_AGEMA_signal_11537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6504 ( .C (clk), .D (new_AGEMA_signal_11540), .Q (new_AGEMA_signal_11541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6508 ( .C (clk), .D (new_AGEMA_signal_11544), .Q (new_AGEMA_signal_11545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6512 ( .C (clk), .D (new_AGEMA_signal_11548), .Q (new_AGEMA_signal_11549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6516 ( .C (clk), .D (new_AGEMA_signal_11552), .Q (new_AGEMA_signal_11553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6520 ( .C (clk), .D (new_AGEMA_signal_11556), .Q (new_AGEMA_signal_11557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6524 ( .C (clk), .D (new_AGEMA_signal_11560), .Q (new_AGEMA_signal_11561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6528 ( .C (clk), .D (new_AGEMA_signal_11564), .Q (new_AGEMA_signal_11565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6532 ( .C (clk), .D (new_AGEMA_signal_11568), .Q (new_AGEMA_signal_11569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6536 ( .C (clk), .D (new_AGEMA_signal_11572), .Q (new_AGEMA_signal_11573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6540 ( .C (clk), .D (new_AGEMA_signal_11576), .Q (new_AGEMA_signal_11577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6544 ( .C (clk), .D (new_AGEMA_signal_11580), .Q (new_AGEMA_signal_11581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6548 ( .C (clk), .D (new_AGEMA_signal_11584), .Q (new_AGEMA_signal_11585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6552 ( .C (clk), .D (new_AGEMA_signal_11588), .Q (new_AGEMA_signal_11589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6556 ( .C (clk), .D (new_AGEMA_signal_11592), .Q (new_AGEMA_signal_11593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6560 ( .C (clk), .D (new_AGEMA_signal_11596), .Q (new_AGEMA_signal_11597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6564 ( .C (clk), .D (new_AGEMA_signal_11600), .Q (new_AGEMA_signal_11601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6568 ( .C (clk), .D (new_AGEMA_signal_11604), .Q (new_AGEMA_signal_11605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6572 ( .C (clk), .D (new_AGEMA_signal_11608), .Q (new_AGEMA_signal_11609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6576 ( .C (clk), .D (new_AGEMA_signal_11612), .Q (new_AGEMA_signal_11613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6580 ( .C (clk), .D (new_AGEMA_signal_11616), .Q (new_AGEMA_signal_11617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6584 ( .C (clk), .D (new_AGEMA_signal_11620), .Q (new_AGEMA_signal_11621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6588 ( .C (clk), .D (new_AGEMA_signal_11624), .Q (new_AGEMA_signal_11625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6592 ( .C (clk), .D (new_AGEMA_signal_11628), .Q (new_AGEMA_signal_11629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6596 ( .C (clk), .D (new_AGEMA_signal_11632), .Q (new_AGEMA_signal_11633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6600 ( .C (clk), .D (new_AGEMA_signal_11636), .Q (new_AGEMA_signal_11637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6604 ( .C (clk), .D (new_AGEMA_signal_11640), .Q (new_AGEMA_signal_11641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6608 ( .C (clk), .D (new_AGEMA_signal_11644), .Q (new_AGEMA_signal_11645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6612 ( .C (clk), .D (new_AGEMA_signal_11648), .Q (new_AGEMA_signal_11649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6616 ( .C (clk), .D (new_AGEMA_signal_11652), .Q (new_AGEMA_signal_11653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6620 ( .C (clk), .D (new_AGEMA_signal_11656), .Q (new_AGEMA_signal_11657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6624 ( .C (clk), .D (new_AGEMA_signal_11660), .Q (new_AGEMA_signal_11661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6628 ( .C (clk), .D (new_AGEMA_signal_11664), .Q (new_AGEMA_signal_11665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6632 ( .C (clk), .D (new_AGEMA_signal_11668), .Q (new_AGEMA_signal_11669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6636 ( .C (clk), .D (new_AGEMA_signal_11672), .Q (new_AGEMA_signal_11673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6640 ( .C (clk), .D (new_AGEMA_signal_11676), .Q (new_AGEMA_signal_11677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6644 ( .C (clk), .D (new_AGEMA_signal_11680), .Q (new_AGEMA_signal_11681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6648 ( .C (clk), .D (new_AGEMA_signal_11684), .Q (new_AGEMA_signal_11685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6652 ( .C (clk), .D (new_AGEMA_signal_11688), .Q (new_AGEMA_signal_11689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6656 ( .C (clk), .D (new_AGEMA_signal_11692), .Q (new_AGEMA_signal_11693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6660 ( .C (clk), .D (new_AGEMA_signal_11696), .Q (new_AGEMA_signal_11697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6664 ( .C (clk), .D (new_AGEMA_signal_11700), .Q (new_AGEMA_signal_11701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6668 ( .C (clk), .D (new_AGEMA_signal_11704), .Q (new_AGEMA_signal_11705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6672 ( .C (clk), .D (new_AGEMA_signal_11708), .Q (new_AGEMA_signal_11709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6676 ( .C (clk), .D (new_AGEMA_signal_11712), .Q (new_AGEMA_signal_11713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6680 ( .C (clk), .D (new_AGEMA_signal_11716), .Q (new_AGEMA_signal_11717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6684 ( .C (clk), .D (new_AGEMA_signal_11720), .Q (new_AGEMA_signal_11721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6688 ( .C (clk), .D (new_AGEMA_signal_11724), .Q (new_AGEMA_signal_11725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6692 ( .C (clk), .D (new_AGEMA_signal_11728), .Q (new_AGEMA_signal_11729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6696 ( .C (clk), .D (new_AGEMA_signal_11732), .Q (new_AGEMA_signal_11733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6700 ( .C (clk), .D (new_AGEMA_signal_11736), .Q (new_AGEMA_signal_11737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6704 ( .C (clk), .D (new_AGEMA_signal_11740), .Q (new_AGEMA_signal_11741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6708 ( .C (clk), .D (new_AGEMA_signal_11744), .Q (new_AGEMA_signal_11745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6712 ( .C (clk), .D (new_AGEMA_signal_11748), .Q (new_AGEMA_signal_11749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6716 ( .C (clk), .D (new_AGEMA_signal_11752), .Q (new_AGEMA_signal_11753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6720 ( .C (clk), .D (new_AGEMA_signal_11756), .Q (new_AGEMA_signal_11757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6724 ( .C (clk), .D (new_AGEMA_signal_11760), .Q (new_AGEMA_signal_11761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6728 ( .C (clk), .D (new_AGEMA_signal_11764), .Q (new_AGEMA_signal_11765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6732 ( .C (clk), .D (new_AGEMA_signal_11768), .Q (new_AGEMA_signal_11769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6736 ( .C (clk), .D (new_AGEMA_signal_11772), .Q (new_AGEMA_signal_11773) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C (clk), .D (new_AGEMA_signal_11776), .Q (new_AGEMA_signal_11777) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C (clk), .D (new_AGEMA_signal_11780), .Q (new_AGEMA_signal_11781) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C (clk), .D (new_AGEMA_signal_11784), .Q (new_AGEMA_signal_11785) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C (clk), .D (new_AGEMA_signal_11788), .Q (new_AGEMA_signal_11789) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C (clk), .D (new_AGEMA_signal_11792), .Q (new_AGEMA_signal_11793) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C (clk), .D (new_AGEMA_signal_11796), .Q (new_AGEMA_signal_11797) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C (clk), .D (new_AGEMA_signal_11800), .Q (new_AGEMA_signal_11801) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C (clk), .D (new_AGEMA_signal_11804), .Q (new_AGEMA_signal_11805) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C (clk), .D (new_AGEMA_signal_11808), .Q (new_AGEMA_signal_11809) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C (clk), .D (new_AGEMA_signal_11812), .Q (new_AGEMA_signal_11813) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C (clk), .D (new_AGEMA_signal_11816), .Q (new_AGEMA_signal_11817) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C (clk), .D (new_AGEMA_signal_11820), .Q (new_AGEMA_signal_11821) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C (clk), .D (new_AGEMA_signal_11824), .Q (new_AGEMA_signal_11825) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C (clk), .D (new_AGEMA_signal_11828), .Q (new_AGEMA_signal_11829) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C (clk), .D (new_AGEMA_signal_11832), .Q (new_AGEMA_signal_11833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6800 ( .C (clk), .D (new_AGEMA_signal_11836), .Q (new_AGEMA_signal_11837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6804 ( .C (clk), .D (new_AGEMA_signal_11840), .Q (new_AGEMA_signal_11841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6808 ( .C (clk), .D (new_AGEMA_signal_11844), .Q (new_AGEMA_signal_11845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6812 ( .C (clk), .D (new_AGEMA_signal_11848), .Q (new_AGEMA_signal_11849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6816 ( .C (clk), .D (new_AGEMA_signal_11852), .Q (new_AGEMA_signal_11853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6820 ( .C (clk), .D (new_AGEMA_signal_11856), .Q (new_AGEMA_signal_11857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6824 ( .C (clk), .D (new_AGEMA_signal_11860), .Q (new_AGEMA_signal_11861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6828 ( .C (clk), .D (new_AGEMA_signal_11864), .Q (new_AGEMA_signal_11865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6832 ( .C (clk), .D (new_AGEMA_signal_11868), .Q (new_AGEMA_signal_11869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6836 ( .C (clk), .D (new_AGEMA_signal_11872), .Q (new_AGEMA_signal_11873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6840 ( .C (clk), .D (new_AGEMA_signal_11876), .Q (new_AGEMA_signal_11877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6844 ( .C (clk), .D (new_AGEMA_signal_11880), .Q (new_AGEMA_signal_11881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6848 ( .C (clk), .D (new_AGEMA_signal_11884), .Q (new_AGEMA_signal_11885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6852 ( .C (clk), .D (new_AGEMA_signal_11888), .Q (new_AGEMA_signal_11889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6856 ( .C (clk), .D (new_AGEMA_signal_11892), .Q (new_AGEMA_signal_11893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6860 ( .C (clk), .D (new_AGEMA_signal_11896), .Q (new_AGEMA_signal_11897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6864 ( .C (clk), .D (new_AGEMA_signal_11900), .Q (new_AGEMA_signal_11901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6868 ( .C (clk), .D (new_AGEMA_signal_11904), .Q (new_AGEMA_signal_11905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6872 ( .C (clk), .D (new_AGEMA_signal_11908), .Q (new_AGEMA_signal_11909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6876 ( .C (clk), .D (new_AGEMA_signal_11912), .Q (new_AGEMA_signal_11913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6880 ( .C (clk), .D (new_AGEMA_signal_11916), .Q (new_AGEMA_signal_11917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6884 ( .C (clk), .D (new_AGEMA_signal_11920), .Q (new_AGEMA_signal_11921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6888 ( .C (clk), .D (new_AGEMA_signal_11924), .Q (new_AGEMA_signal_11925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6892 ( .C (clk), .D (new_AGEMA_signal_11928), .Q (new_AGEMA_signal_11929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6896 ( .C (clk), .D (new_AGEMA_signal_11932), .Q (new_AGEMA_signal_11933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6900 ( .C (clk), .D (new_AGEMA_signal_11936), .Q (new_AGEMA_signal_11937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6904 ( .C (clk), .D (new_AGEMA_signal_11940), .Q (new_AGEMA_signal_11941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6908 ( .C (clk), .D (new_AGEMA_signal_11944), .Q (new_AGEMA_signal_11945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6912 ( .C (clk), .D (new_AGEMA_signal_11948), .Q (new_AGEMA_signal_11949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6916 ( .C (clk), .D (new_AGEMA_signal_11952), .Q (new_AGEMA_signal_11953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6920 ( .C (clk), .D (new_AGEMA_signal_11956), .Q (new_AGEMA_signal_11957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6924 ( .C (clk), .D (new_AGEMA_signal_11960), .Q (new_AGEMA_signal_11961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6928 ( .C (clk), .D (new_AGEMA_signal_11964), .Q (new_AGEMA_signal_11965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6932 ( .C (clk), .D (new_AGEMA_signal_11968), .Q (new_AGEMA_signal_11969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6936 ( .C (clk), .D (new_AGEMA_signal_11972), .Q (new_AGEMA_signal_11973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6940 ( .C (clk), .D (new_AGEMA_signal_11976), .Q (new_AGEMA_signal_11977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6944 ( .C (clk), .D (new_AGEMA_signal_11980), .Q (new_AGEMA_signal_11981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6948 ( .C (clk), .D (new_AGEMA_signal_11984), .Q (new_AGEMA_signal_11985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6952 ( .C (clk), .D (new_AGEMA_signal_11988), .Q (new_AGEMA_signal_11989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6956 ( .C (clk), .D (new_AGEMA_signal_11992), .Q (new_AGEMA_signal_11993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6960 ( .C (clk), .D (new_AGEMA_signal_11996), .Q (new_AGEMA_signal_11997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6964 ( .C (clk), .D (new_AGEMA_signal_12000), .Q (new_AGEMA_signal_12001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6968 ( .C (clk), .D (new_AGEMA_signal_12004), .Q (new_AGEMA_signal_12005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6972 ( .C (clk), .D (new_AGEMA_signal_12008), .Q (new_AGEMA_signal_12009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6976 ( .C (clk), .D (new_AGEMA_signal_12012), .Q (new_AGEMA_signal_12013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6980 ( .C (clk), .D (new_AGEMA_signal_12016), .Q (new_AGEMA_signal_12017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6984 ( .C (clk), .D (new_AGEMA_signal_12020), .Q (new_AGEMA_signal_12021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6988 ( .C (clk), .D (new_AGEMA_signal_12024), .Q (new_AGEMA_signal_12025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6992 ( .C (clk), .D (new_AGEMA_signal_12028), .Q (new_AGEMA_signal_12029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6996 ( .C (clk), .D (new_AGEMA_signal_12032), .Q (new_AGEMA_signal_12033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7000 ( .C (clk), .D (new_AGEMA_signal_12036), .Q (new_AGEMA_signal_12037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7004 ( .C (clk), .D (new_AGEMA_signal_12040), .Q (new_AGEMA_signal_12041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7008 ( .C (clk), .D (new_AGEMA_signal_12044), .Q (new_AGEMA_signal_12045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7012 ( .C (clk), .D (new_AGEMA_signal_12048), .Q (new_AGEMA_signal_12049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7016 ( .C (clk), .D (new_AGEMA_signal_12052), .Q (new_AGEMA_signal_12053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7020 ( .C (clk), .D (new_AGEMA_signal_12056), .Q (new_AGEMA_signal_12057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7024 ( .C (clk), .D (new_AGEMA_signal_12060), .Q (new_AGEMA_signal_12061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7028 ( .C (clk), .D (new_AGEMA_signal_12064), .Q (new_AGEMA_signal_12065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7032 ( .C (clk), .D (new_AGEMA_signal_12068), .Q (new_AGEMA_signal_12069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7036 ( .C (clk), .D (new_AGEMA_signal_12072), .Q (new_AGEMA_signal_12073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7040 ( .C (clk), .D (new_AGEMA_signal_12076), .Q (new_AGEMA_signal_12077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7044 ( .C (clk), .D (new_AGEMA_signal_12080), .Q (new_AGEMA_signal_12081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7048 ( .C (clk), .D (new_AGEMA_signal_12084), .Q (new_AGEMA_signal_12085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7052 ( .C (clk), .D (new_AGEMA_signal_12088), .Q (new_AGEMA_signal_12089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7056 ( .C (clk), .D (new_AGEMA_signal_12092), .Q (new_AGEMA_signal_12093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7060 ( .C (clk), .D (new_AGEMA_signal_12096), .Q (new_AGEMA_signal_12097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7064 ( .C (clk), .D (new_AGEMA_signal_12100), .Q (new_AGEMA_signal_12101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7068 ( .C (clk), .D (new_AGEMA_signal_12104), .Q (new_AGEMA_signal_12105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7072 ( .C (clk), .D (new_AGEMA_signal_12108), .Q (new_AGEMA_signal_12109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7076 ( .C (clk), .D (new_AGEMA_signal_12112), .Q (new_AGEMA_signal_12113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7080 ( .C (clk), .D (new_AGEMA_signal_12116), .Q (new_AGEMA_signal_12117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7084 ( .C (clk), .D (new_AGEMA_signal_12120), .Q (new_AGEMA_signal_12121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7088 ( .C (clk), .D (new_AGEMA_signal_12124), .Q (new_AGEMA_signal_12125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7092 ( .C (clk), .D (new_AGEMA_signal_12128), .Q (new_AGEMA_signal_12129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7096 ( .C (clk), .D (new_AGEMA_signal_12132), .Q (new_AGEMA_signal_12133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7100 ( .C (clk), .D (new_AGEMA_signal_12136), .Q (new_AGEMA_signal_12137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7104 ( .C (clk), .D (new_AGEMA_signal_12140), .Q (new_AGEMA_signal_12141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7108 ( .C (clk), .D (new_AGEMA_signal_12144), .Q (new_AGEMA_signal_12145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7112 ( .C (clk), .D (new_AGEMA_signal_12148), .Q (new_AGEMA_signal_12149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7116 ( .C (clk), .D (new_AGEMA_signal_12152), .Q (new_AGEMA_signal_12153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7120 ( .C (clk), .D (new_AGEMA_signal_12156), .Q (new_AGEMA_signal_12157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7124 ( .C (clk), .D (new_AGEMA_signal_12160), .Q (new_AGEMA_signal_12161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7128 ( .C (clk), .D (new_AGEMA_signal_12164), .Q (new_AGEMA_signal_12165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7132 ( .C (clk), .D (new_AGEMA_signal_12168), .Q (new_AGEMA_signal_12169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7136 ( .C (clk), .D (new_AGEMA_signal_12172), .Q (new_AGEMA_signal_12173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7140 ( .C (clk), .D (new_AGEMA_signal_12176), .Q (new_AGEMA_signal_12177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7144 ( .C (clk), .D (new_AGEMA_signal_12180), .Q (new_AGEMA_signal_12181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7148 ( .C (clk), .D (new_AGEMA_signal_12184), .Q (new_AGEMA_signal_12185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7152 ( .C (clk), .D (new_AGEMA_signal_12188), .Q (new_AGEMA_signal_12189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7156 ( .C (clk), .D (new_AGEMA_signal_12192), .Q (new_AGEMA_signal_12193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7160 ( .C (clk), .D (new_AGEMA_signal_12196), .Q (new_AGEMA_signal_12197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7164 ( .C (clk), .D (new_AGEMA_signal_12200), .Q (new_AGEMA_signal_12201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7168 ( .C (clk), .D (new_AGEMA_signal_12204), .Q (new_AGEMA_signal_12205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7172 ( .C (clk), .D (new_AGEMA_signal_12208), .Q (new_AGEMA_signal_12209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7176 ( .C (clk), .D (new_AGEMA_signal_12212), .Q (new_AGEMA_signal_12213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7180 ( .C (clk), .D (new_AGEMA_signal_12216), .Q (new_AGEMA_signal_12217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7184 ( .C (clk), .D (new_AGEMA_signal_12220), .Q (new_AGEMA_signal_12221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7188 ( .C (clk), .D (new_AGEMA_signal_12224), .Q (new_AGEMA_signal_12225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7192 ( .C (clk), .D (new_AGEMA_signal_12228), .Q (new_AGEMA_signal_12229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7196 ( .C (clk), .D (new_AGEMA_signal_12232), .Q (new_AGEMA_signal_12233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7200 ( .C (clk), .D (new_AGEMA_signal_12236), .Q (new_AGEMA_signal_12237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7204 ( .C (clk), .D (new_AGEMA_signal_12240), .Q (new_AGEMA_signal_12241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7208 ( .C (clk), .D (new_AGEMA_signal_12244), .Q (new_AGEMA_signal_12245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7212 ( .C (clk), .D (new_AGEMA_signal_12248), .Q (new_AGEMA_signal_12249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7216 ( .C (clk), .D (new_AGEMA_signal_12252), .Q (new_AGEMA_signal_12253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7220 ( .C (clk), .D (new_AGEMA_signal_12256), .Q (new_AGEMA_signal_12257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7224 ( .C (clk), .D (new_AGEMA_signal_12260), .Q (new_AGEMA_signal_12261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7228 ( .C (clk), .D (new_AGEMA_signal_12264), .Q (new_AGEMA_signal_12265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7232 ( .C (clk), .D (new_AGEMA_signal_12268), .Q (new_AGEMA_signal_12269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7236 ( .C (clk), .D (new_AGEMA_signal_12272), .Q (new_AGEMA_signal_12273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7240 ( .C (clk), .D (new_AGEMA_signal_12276), .Q (new_AGEMA_signal_12277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7244 ( .C (clk), .D (new_AGEMA_signal_12280), .Q (new_AGEMA_signal_12281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7248 ( .C (clk), .D (new_AGEMA_signal_12284), .Q (new_AGEMA_signal_12285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7252 ( .C (clk), .D (new_AGEMA_signal_12288), .Q (new_AGEMA_signal_12289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7256 ( .C (clk), .D (new_AGEMA_signal_12292), .Q (new_AGEMA_signal_12293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7260 ( .C (clk), .D (new_AGEMA_signal_12296), .Q (new_AGEMA_signal_12297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7264 ( .C (clk), .D (new_AGEMA_signal_12300), .Q (new_AGEMA_signal_12301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7268 ( .C (clk), .D (new_AGEMA_signal_12304), .Q (new_AGEMA_signal_12305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7272 ( .C (clk), .D (new_AGEMA_signal_12308), .Q (new_AGEMA_signal_12309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7276 ( .C (clk), .D (new_AGEMA_signal_12312), .Q (new_AGEMA_signal_12313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7280 ( .C (clk), .D (new_AGEMA_signal_12316), .Q (new_AGEMA_signal_12317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7284 ( .C (clk), .D (new_AGEMA_signal_12320), .Q (new_AGEMA_signal_12321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7288 ( .C (clk), .D (new_AGEMA_signal_12324), .Q (new_AGEMA_signal_12325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7292 ( .C (clk), .D (new_AGEMA_signal_12328), .Q (new_AGEMA_signal_12329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7296 ( .C (clk), .D (new_AGEMA_signal_12332), .Q (new_AGEMA_signal_12333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7300 ( .C (clk), .D (new_AGEMA_signal_12336), .Q (new_AGEMA_signal_12337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7304 ( .C (clk), .D (new_AGEMA_signal_12340), .Q (new_AGEMA_signal_12341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7308 ( .C (clk), .D (new_AGEMA_signal_12344), .Q (new_AGEMA_signal_12345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7312 ( .C (clk), .D (new_AGEMA_signal_12348), .Q (new_AGEMA_signal_12349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7316 ( .C (clk), .D (new_AGEMA_signal_12352), .Q (new_AGEMA_signal_12353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7320 ( .C (clk), .D (new_AGEMA_signal_12356), .Q (new_AGEMA_signal_12357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7324 ( .C (clk), .D (new_AGEMA_signal_12360), .Q (new_AGEMA_signal_12361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7328 ( .C (clk), .D (new_AGEMA_signal_12364), .Q (new_AGEMA_signal_12365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7332 ( .C (clk), .D (new_AGEMA_signal_12368), .Q (new_AGEMA_signal_12369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7336 ( .C (clk), .D (new_AGEMA_signal_12372), .Q (new_AGEMA_signal_12373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7340 ( .C (clk), .D (new_AGEMA_signal_12376), .Q (new_AGEMA_signal_12377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7344 ( .C (clk), .D (new_AGEMA_signal_12380), .Q (new_AGEMA_signal_12381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7348 ( .C (clk), .D (new_AGEMA_signal_12384), .Q (new_AGEMA_signal_12385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7352 ( .C (clk), .D (new_AGEMA_signal_12388), .Q (new_AGEMA_signal_12389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7356 ( .C (clk), .D (new_AGEMA_signal_12392), .Q (new_AGEMA_signal_12393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7360 ( .C (clk), .D (new_AGEMA_signal_12396), .Q (new_AGEMA_signal_12397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7364 ( .C (clk), .D (new_AGEMA_signal_12400), .Q (new_AGEMA_signal_12401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7368 ( .C (clk), .D (new_AGEMA_signal_12404), .Q (new_AGEMA_signal_12405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7372 ( .C (clk), .D (new_AGEMA_signal_12408), .Q (new_AGEMA_signal_12409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7376 ( .C (clk), .D (new_AGEMA_signal_12412), .Q (new_AGEMA_signal_12413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7380 ( .C (clk), .D (new_AGEMA_signal_12416), .Q (new_AGEMA_signal_12417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7384 ( .C (clk), .D (new_AGEMA_signal_12420), .Q (new_AGEMA_signal_12421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7388 ( .C (clk), .D (new_AGEMA_signal_12424), .Q (new_AGEMA_signal_12425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7392 ( .C (clk), .D (new_AGEMA_signal_12428), .Q (new_AGEMA_signal_12429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7396 ( .C (clk), .D (new_AGEMA_signal_12432), .Q (new_AGEMA_signal_12433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7400 ( .C (clk), .D (new_AGEMA_signal_12436), .Q (new_AGEMA_signal_12437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7404 ( .C (clk), .D (new_AGEMA_signal_12440), .Q (new_AGEMA_signal_12441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7408 ( .C (clk), .D (new_AGEMA_signal_12444), .Q (new_AGEMA_signal_12445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7412 ( .C (clk), .D (new_AGEMA_signal_12448), .Q (new_AGEMA_signal_12449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7416 ( .C (clk), .D (new_AGEMA_signal_12452), .Q (new_AGEMA_signal_12453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7420 ( .C (clk), .D (new_AGEMA_signal_12456), .Q (new_AGEMA_signal_12457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7424 ( .C (clk), .D (new_AGEMA_signal_12460), .Q (new_AGEMA_signal_12461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7428 ( .C (clk), .D (new_AGEMA_signal_12464), .Q (new_AGEMA_signal_12465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7432 ( .C (clk), .D (new_AGEMA_signal_12468), .Q (new_AGEMA_signal_12469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7436 ( .C (clk), .D (new_AGEMA_signal_12472), .Q (new_AGEMA_signal_12473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7440 ( .C (clk), .D (new_AGEMA_signal_12476), .Q (new_AGEMA_signal_12477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7444 ( .C (clk), .D (new_AGEMA_signal_12480), .Q (new_AGEMA_signal_12481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7448 ( .C (clk), .D (new_AGEMA_signal_12484), .Q (new_AGEMA_signal_12485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7452 ( .C (clk), .D (new_AGEMA_signal_12488), .Q (new_AGEMA_signal_12489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7456 ( .C (clk), .D (new_AGEMA_signal_12492), .Q (new_AGEMA_signal_12493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7460 ( .C (clk), .D (new_AGEMA_signal_12496), .Q (new_AGEMA_signal_12497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7464 ( .C (clk), .D (new_AGEMA_signal_12500), .Q (new_AGEMA_signal_12501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7468 ( .C (clk), .D (new_AGEMA_signal_12504), .Q (new_AGEMA_signal_12505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7472 ( .C (clk), .D (new_AGEMA_signal_12508), .Q (new_AGEMA_signal_12509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7476 ( .C (clk), .D (new_AGEMA_signal_12512), .Q (new_AGEMA_signal_12513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7480 ( .C (clk), .D (new_AGEMA_signal_12516), .Q (new_AGEMA_signal_12517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7484 ( .C (clk), .D (new_AGEMA_signal_12520), .Q (new_AGEMA_signal_12521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7488 ( .C (clk), .D (new_AGEMA_signal_12524), .Q (new_AGEMA_signal_12525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7492 ( .C (clk), .D (new_AGEMA_signal_12528), .Q (new_AGEMA_signal_12529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7496 ( .C (clk), .D (new_AGEMA_signal_12532), .Q (new_AGEMA_signal_12533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7500 ( .C (clk), .D (new_AGEMA_signal_12536), .Q (new_AGEMA_signal_12537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7504 ( .C (clk), .D (new_AGEMA_signal_12540), .Q (new_AGEMA_signal_12541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7508 ( .C (clk), .D (new_AGEMA_signal_12544), .Q (new_AGEMA_signal_12545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7512 ( .C (clk), .D (new_AGEMA_signal_12548), .Q (new_AGEMA_signal_12549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7516 ( .C (clk), .D (new_AGEMA_signal_12552), .Q (new_AGEMA_signal_12553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7520 ( .C (clk), .D (new_AGEMA_signal_12556), .Q (new_AGEMA_signal_12557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7524 ( .C (clk), .D (new_AGEMA_signal_12560), .Q (new_AGEMA_signal_12561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7528 ( .C (clk), .D (new_AGEMA_signal_12564), .Q (new_AGEMA_signal_12565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7532 ( .C (clk), .D (new_AGEMA_signal_12568), .Q (new_AGEMA_signal_12569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7536 ( .C (clk), .D (new_AGEMA_signal_12572), .Q (new_AGEMA_signal_12573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7540 ( .C (clk), .D (new_AGEMA_signal_12576), .Q (new_AGEMA_signal_12577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7544 ( .C (clk), .D (new_AGEMA_signal_12580), .Q (new_AGEMA_signal_12581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7548 ( .C (clk), .D (new_AGEMA_signal_12584), .Q (new_AGEMA_signal_12585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7552 ( .C (clk), .D (new_AGEMA_signal_12588), .Q (new_AGEMA_signal_12589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7556 ( .C (clk), .D (new_AGEMA_signal_12592), .Q (new_AGEMA_signal_12593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7560 ( .C (clk), .D (new_AGEMA_signal_12596), .Q (new_AGEMA_signal_12597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7564 ( .C (clk), .D (new_AGEMA_signal_12600), .Q (new_AGEMA_signal_12601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7568 ( .C (clk), .D (new_AGEMA_signal_12604), .Q (new_AGEMA_signal_12605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7572 ( .C (clk), .D (new_AGEMA_signal_12608), .Q (new_AGEMA_signal_12609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7576 ( .C (clk), .D (new_AGEMA_signal_12612), .Q (new_AGEMA_signal_12613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7580 ( .C (clk), .D (new_AGEMA_signal_12616), .Q (new_AGEMA_signal_12617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7584 ( .C (clk), .D (new_AGEMA_signal_12620), .Q (new_AGEMA_signal_12621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7588 ( .C (clk), .D (new_AGEMA_signal_12624), .Q (new_AGEMA_signal_12625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7592 ( .C (clk), .D (new_AGEMA_signal_12628), .Q (new_AGEMA_signal_12629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7596 ( .C (clk), .D (new_AGEMA_signal_12632), .Q (new_AGEMA_signal_12633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7600 ( .C (clk), .D (new_AGEMA_signal_12636), .Q (new_AGEMA_signal_12637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7604 ( .C (clk), .D (new_AGEMA_signal_12640), .Q (new_AGEMA_signal_12641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7608 ( .C (clk), .D (new_AGEMA_signal_12644), .Q (new_AGEMA_signal_12645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7612 ( .C (clk), .D (new_AGEMA_signal_12648), .Q (new_AGEMA_signal_12649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7616 ( .C (clk), .D (new_AGEMA_signal_12652), .Q (new_AGEMA_signal_12653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7620 ( .C (clk), .D (new_AGEMA_signal_12656), .Q (new_AGEMA_signal_12657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7624 ( .C (clk), .D (new_AGEMA_signal_12660), .Q (new_AGEMA_signal_12661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7628 ( .C (clk), .D (new_AGEMA_signal_12664), .Q (new_AGEMA_signal_12665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7632 ( .C (clk), .D (new_AGEMA_signal_12668), .Q (new_AGEMA_signal_12669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7636 ( .C (clk), .D (new_AGEMA_signal_12672), .Q (new_AGEMA_signal_12673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7640 ( .C (clk), .D (new_AGEMA_signal_12676), .Q (new_AGEMA_signal_12677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7644 ( .C (clk), .D (new_AGEMA_signal_12680), .Q (new_AGEMA_signal_12681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7648 ( .C (clk), .D (new_AGEMA_signal_12684), .Q (new_AGEMA_signal_12685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7652 ( .C (clk), .D (new_AGEMA_signal_12688), .Q (new_AGEMA_signal_12689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7656 ( .C (clk), .D (new_AGEMA_signal_12692), .Q (new_AGEMA_signal_12693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7660 ( .C (clk), .D (new_AGEMA_signal_12696), .Q (new_AGEMA_signal_12697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7664 ( .C (clk), .D (new_AGEMA_signal_12700), .Q (new_AGEMA_signal_12701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7668 ( .C (clk), .D (new_AGEMA_signal_12704), .Q (new_AGEMA_signal_12705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7672 ( .C (clk), .D (new_AGEMA_signal_12708), .Q (new_AGEMA_signal_12709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7676 ( .C (clk), .D (new_AGEMA_signal_12712), .Q (new_AGEMA_signal_12713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7680 ( .C (clk), .D (new_AGEMA_signal_12716), .Q (new_AGEMA_signal_12717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7684 ( .C (clk), .D (new_AGEMA_signal_12720), .Q (new_AGEMA_signal_12721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7688 ( .C (clk), .D (new_AGEMA_signal_12724), .Q (new_AGEMA_signal_12725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7692 ( .C (clk), .D (new_AGEMA_signal_12728), .Q (new_AGEMA_signal_12729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7696 ( .C (clk), .D (new_AGEMA_signal_12732), .Q (new_AGEMA_signal_12733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7700 ( .C (clk), .D (new_AGEMA_signal_12736), .Q (new_AGEMA_signal_12737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7704 ( .C (clk), .D (new_AGEMA_signal_12740), .Q (new_AGEMA_signal_12741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7708 ( .C (clk), .D (new_AGEMA_signal_12744), .Q (new_AGEMA_signal_12745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7712 ( .C (clk), .D (new_AGEMA_signal_12748), .Q (new_AGEMA_signal_12749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7716 ( .C (clk), .D (new_AGEMA_signal_12752), .Q (new_AGEMA_signal_12753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7720 ( .C (clk), .D (new_AGEMA_signal_12756), .Q (new_AGEMA_signal_12757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7724 ( .C (clk), .D (new_AGEMA_signal_12760), .Q (new_AGEMA_signal_12761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7728 ( .C (clk), .D (new_AGEMA_signal_12764), .Q (new_AGEMA_signal_12765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7732 ( .C (clk), .D (new_AGEMA_signal_12768), .Q (new_AGEMA_signal_12769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7736 ( .C (clk), .D (new_AGEMA_signal_12772), .Q (new_AGEMA_signal_12773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7740 ( .C (clk), .D (new_AGEMA_signal_12776), .Q (new_AGEMA_signal_12777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7744 ( .C (clk), .D (new_AGEMA_signal_12780), .Q (new_AGEMA_signal_12781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7748 ( .C (clk), .D (new_AGEMA_signal_12784), .Q (new_AGEMA_signal_12785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7752 ( .C (clk), .D (new_AGEMA_signal_12788), .Q (new_AGEMA_signal_12789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7756 ( .C (clk), .D (new_AGEMA_signal_12792), .Q (new_AGEMA_signal_12793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7760 ( .C (clk), .D (new_AGEMA_signal_12796), .Q (new_AGEMA_signal_12797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7764 ( .C (clk), .D (new_AGEMA_signal_12800), .Q (new_AGEMA_signal_12801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7768 ( .C (clk), .D (new_AGEMA_signal_12804), .Q (new_AGEMA_signal_12805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7772 ( .C (clk), .D (new_AGEMA_signal_12808), .Q (new_AGEMA_signal_12809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7776 ( .C (clk), .D (new_AGEMA_signal_12812), .Q (new_AGEMA_signal_12813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7780 ( .C (clk), .D (new_AGEMA_signal_12816), .Q (new_AGEMA_signal_12817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7784 ( .C (clk), .D (new_AGEMA_signal_12820), .Q (new_AGEMA_signal_12821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7788 ( .C (clk), .D (new_AGEMA_signal_12824), .Q (new_AGEMA_signal_12825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7792 ( .C (clk), .D (new_AGEMA_signal_12828), .Q (new_AGEMA_signal_12829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7796 ( .C (clk), .D (new_AGEMA_signal_12832), .Q (new_AGEMA_signal_12833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7800 ( .C (clk), .D (new_AGEMA_signal_12836), .Q (new_AGEMA_signal_12837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7804 ( .C (clk), .D (new_AGEMA_signal_12840), .Q (new_AGEMA_signal_12841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7808 ( .C (clk), .D (new_AGEMA_signal_12844), .Q (new_AGEMA_signal_12845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7812 ( .C (clk), .D (new_AGEMA_signal_12848), .Q (new_AGEMA_signal_12849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7816 ( .C (clk), .D (new_AGEMA_signal_12852), .Q (new_AGEMA_signal_12853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7820 ( .C (clk), .D (new_AGEMA_signal_12856), .Q (new_AGEMA_signal_12857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7824 ( .C (clk), .D (new_AGEMA_signal_12860), .Q (new_AGEMA_signal_12861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7828 ( .C (clk), .D (new_AGEMA_signal_12864), .Q (new_AGEMA_signal_12865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7832 ( .C (clk), .D (new_AGEMA_signal_12868), .Q (new_AGEMA_signal_12869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7836 ( .C (clk), .D (new_AGEMA_signal_12872), .Q (new_AGEMA_signal_12873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7840 ( .C (clk), .D (new_AGEMA_signal_12876), .Q (new_AGEMA_signal_12877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7844 ( .C (clk), .D (new_AGEMA_signal_12880), .Q (new_AGEMA_signal_12881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7848 ( .C (clk), .D (new_AGEMA_signal_12884), .Q (new_AGEMA_signal_12885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7852 ( .C (clk), .D (new_AGEMA_signal_12888), .Q (new_AGEMA_signal_12889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7856 ( .C (clk), .D (new_AGEMA_signal_12892), .Q (new_AGEMA_signal_12893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7860 ( .C (clk), .D (new_AGEMA_signal_12896), .Q (new_AGEMA_signal_12897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7864 ( .C (clk), .D (new_AGEMA_signal_12900), .Q (new_AGEMA_signal_12901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7868 ( .C (clk), .D (new_AGEMA_signal_12904), .Q (new_AGEMA_signal_12905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7872 ( .C (clk), .D (new_AGEMA_signal_12908), .Q (new_AGEMA_signal_12909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7876 ( .C (clk), .D (new_AGEMA_signal_12912), .Q (new_AGEMA_signal_12913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7880 ( .C (clk), .D (new_AGEMA_signal_12916), .Q (new_AGEMA_signal_12917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7884 ( .C (clk), .D (new_AGEMA_signal_12920), .Q (new_AGEMA_signal_12921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7888 ( .C (clk), .D (new_AGEMA_signal_12924), .Q (new_AGEMA_signal_12925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7892 ( .C (clk), .D (new_AGEMA_signal_12928), .Q (new_AGEMA_signal_12929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7896 ( .C (clk), .D (new_AGEMA_signal_12932), .Q (new_AGEMA_signal_12933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7900 ( .C (clk), .D (new_AGEMA_signal_12936), .Q (new_AGEMA_signal_12937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7904 ( .C (clk), .D (new_AGEMA_signal_12940), .Q (new_AGEMA_signal_12941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7908 ( .C (clk), .D (new_AGEMA_signal_12944), .Q (new_AGEMA_signal_12945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7912 ( .C (clk), .D (new_AGEMA_signal_12948), .Q (new_AGEMA_signal_12949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7916 ( .C (clk), .D (new_AGEMA_signal_12952), .Q (new_AGEMA_signal_12953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7920 ( .C (clk), .D (new_AGEMA_signal_12956), .Q (new_AGEMA_signal_12957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7924 ( .C (clk), .D (new_AGEMA_signal_12960), .Q (new_AGEMA_signal_12961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7928 ( .C (clk), .D (new_AGEMA_signal_12964), .Q (new_AGEMA_signal_12965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7932 ( .C (clk), .D (new_AGEMA_signal_12968), .Q (new_AGEMA_signal_12969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7936 ( .C (clk), .D (new_AGEMA_signal_12972), .Q (new_AGEMA_signal_12973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7940 ( .C (clk), .D (new_AGEMA_signal_12976), .Q (new_AGEMA_signal_12977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7944 ( .C (clk), .D (new_AGEMA_signal_12980), .Q (new_AGEMA_signal_12981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_7948 ( .C (clk), .D (new_AGEMA_signal_12984), .Q (new_AGEMA_signal_12985) ) ;
    buf_clk new_AGEMA_reg_buffer_7952 ( .C (clk), .D (new_AGEMA_signal_12988), .Q (new_AGEMA_signal_12989) ) ;
    buf_clk new_AGEMA_reg_buffer_7956 ( .C (clk), .D (new_AGEMA_signal_12992), .Q (new_AGEMA_signal_12993) ) ;
    buf_clk new_AGEMA_reg_buffer_7960 ( .C (clk), .D (new_AGEMA_signal_12996), .Q (new_AGEMA_signal_12997) ) ;
    buf_clk new_AGEMA_reg_buffer_7964 ( .C (clk), .D (new_AGEMA_signal_13000), .Q (new_AGEMA_signal_13001) ) ;
    buf_clk new_AGEMA_reg_buffer_7968 ( .C (clk), .D (new_AGEMA_signal_13004), .Q (new_AGEMA_signal_13005) ) ;
    buf_clk new_AGEMA_reg_buffer_7972 ( .C (clk), .D (new_AGEMA_signal_13008), .Q (new_AGEMA_signal_13009) ) ;
    buf_clk new_AGEMA_reg_buffer_7976 ( .C (clk), .D (new_AGEMA_signal_13012), .Q (new_AGEMA_signal_13013) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5975, new_AGEMA_signal_5974, RoundReg_Inst_ff_SDE_0_next_state}), .clk (clk), .Q ({ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6209, new_AGEMA_signal_6208, RoundReg_Inst_ff_SDE_1_next_state}), .clk (clk), .Q ({ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, RoundReg_Inst_ff_SDE_2_next_state}), .clk (clk), .Q ({ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, RoundReg_Inst_ff_SDE_3_next_state}), .clk (clk), .Q ({ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6217, new_AGEMA_signal_6216, RoundReg_Inst_ff_SDE_4_next_state}), .clk (clk), .Q ({ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5983, new_AGEMA_signal_5982, RoundReg_Inst_ff_SDE_5_next_state}), .clk (clk), .Q ({ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5987, new_AGEMA_signal_5986, RoundReg_Inst_ff_SDE_6_next_state}), .clk (clk), .Q ({ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, RoundReg_Inst_ff_SDE_7_next_state}), .clk (clk), .Q ({ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5995, new_AGEMA_signal_5994, RoundReg_Inst_ff_SDE_8_next_state}), .clk (clk), .Q ({ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6221, new_AGEMA_signal_6220, RoundReg_Inst_ff_SDE_9_next_state}), .clk (clk), .Q ({ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5999, new_AGEMA_signal_5998, RoundReg_Inst_ff_SDE_10_next_state}), .clk (clk), .Q ({ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, RoundReg_Inst_ff_SDE_11_next_state}), .clk (clk), .Q ({ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6229, new_AGEMA_signal_6228, RoundReg_Inst_ff_SDE_12_next_state}), .clk (clk), .Q ({ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, RoundReg_Inst_ff_SDE_13_next_state}), .clk (clk), .Q ({ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6007, new_AGEMA_signal_6006, RoundReg_Inst_ff_SDE_14_next_state}), .clk (clk), .Q ({ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6011, new_AGEMA_signal_6010, RoundReg_Inst_ff_SDE_15_next_state}), .clk (clk), .Q ({ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, RoundReg_Inst_ff_SDE_16_next_state}), .clk (clk), .Q ({ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6233, new_AGEMA_signal_6232, RoundReg_Inst_ff_SDE_17_next_state}), .clk (clk), .Q ({ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6019, new_AGEMA_signal_6018, RoundReg_Inst_ff_SDE_18_next_state}), .clk (clk), .Q ({ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, RoundReg_Inst_ff_SDE_19_next_state}), .clk (clk), .Q ({ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6241, new_AGEMA_signal_6240, RoundReg_Inst_ff_SDE_20_next_state}), .clk (clk), .Q ({ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6023, new_AGEMA_signal_6022, RoundReg_Inst_ff_SDE_21_next_state}), .clk (clk), .Q ({ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, RoundReg_Inst_ff_SDE_22_next_state}), .clk (clk), .Q ({ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6031, new_AGEMA_signal_6030, RoundReg_Inst_ff_SDE_23_next_state}), .clk (clk), .Q ({ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6035, new_AGEMA_signal_6034, RoundReg_Inst_ff_SDE_24_next_state}), .clk (clk), .Q ({ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6245, new_AGEMA_signal_6244, RoundReg_Inst_ff_SDE_25_next_state}), .clk (clk), .Q ({ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, RoundReg_Inst_ff_SDE_26_next_state}), .clk (clk), .Q ({ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, RoundReg_Inst_ff_SDE_27_next_state}), .clk (clk), .Q ({ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6253, new_AGEMA_signal_6252, RoundReg_Inst_ff_SDE_28_next_state}), .clk (clk), .Q ({ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6043, new_AGEMA_signal_6042, RoundReg_Inst_ff_SDE_29_next_state}), .clk (clk), .Q ({ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6047, new_AGEMA_signal_6046, RoundReg_Inst_ff_SDE_30_next_state}), .clk (clk), .Q ({ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, RoundReg_Inst_ff_SDE_31_next_state}), .clk (clk), .Q ({ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11845, new_AGEMA_signal_11841, new_AGEMA_signal_11837}), .clk (clk), .Q ({ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11857, new_AGEMA_signal_11853, new_AGEMA_signal_11849}), .clk (clk), .Q ({ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11869, new_AGEMA_signal_11865, new_AGEMA_signal_11861}), .clk (clk), .Q ({ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11881, new_AGEMA_signal_11877, new_AGEMA_signal_11873}), .clk (clk), .Q ({ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11893, new_AGEMA_signal_11889, new_AGEMA_signal_11885}), .clk (clk), .Q ({ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11905, new_AGEMA_signal_11901, new_AGEMA_signal_11897}), .clk (clk), .Q ({ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11917, new_AGEMA_signal_11913, new_AGEMA_signal_11909}), .clk (clk), .Q ({ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11929, new_AGEMA_signal_11925, new_AGEMA_signal_11921}), .clk (clk), .Q ({ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11941, new_AGEMA_signal_11937, new_AGEMA_signal_11933}), .clk (clk), .Q ({ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11953, new_AGEMA_signal_11949, new_AGEMA_signal_11945}), .clk (clk), .Q ({ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11965, new_AGEMA_signal_11961, new_AGEMA_signal_11957}), .clk (clk), .Q ({ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11977, new_AGEMA_signal_11973, new_AGEMA_signal_11969}), .clk (clk), .Q ({ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_11989, new_AGEMA_signal_11985, new_AGEMA_signal_11981}), .clk (clk), .Q ({ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12001, new_AGEMA_signal_11997, new_AGEMA_signal_11993}), .clk (clk), .Q ({ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12013, new_AGEMA_signal_12009, new_AGEMA_signal_12005}), .clk (clk), .Q ({ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12025, new_AGEMA_signal_12021, new_AGEMA_signal_12017}), .clk (clk), .Q ({ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12037, new_AGEMA_signal_12033, new_AGEMA_signal_12029}), .clk (clk), .Q ({ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12049, new_AGEMA_signal_12045, new_AGEMA_signal_12041}), .clk (clk), .Q ({ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12061, new_AGEMA_signal_12057, new_AGEMA_signal_12053}), .clk (clk), .Q ({ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12073, new_AGEMA_signal_12069, new_AGEMA_signal_12065}), .clk (clk), .Q ({ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12085, new_AGEMA_signal_12081, new_AGEMA_signal_12077}), .clk (clk), .Q ({ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12097, new_AGEMA_signal_12093, new_AGEMA_signal_12089}), .clk (clk), .Q ({ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12109, new_AGEMA_signal_12105, new_AGEMA_signal_12101}), .clk (clk), .Q ({ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12121, new_AGEMA_signal_12117, new_AGEMA_signal_12113}), .clk (clk), .Q ({ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12133, new_AGEMA_signal_12129, new_AGEMA_signal_12125}), .clk (clk), .Q ({ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12145, new_AGEMA_signal_12141, new_AGEMA_signal_12137}), .clk (clk), .Q ({ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12157, new_AGEMA_signal_12153, new_AGEMA_signal_12149}), .clk (clk), .Q ({ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12169, new_AGEMA_signal_12165, new_AGEMA_signal_12161}), .clk (clk), .Q ({ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12181, new_AGEMA_signal_12177, new_AGEMA_signal_12173}), .clk (clk), .Q ({ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12193, new_AGEMA_signal_12189, new_AGEMA_signal_12185}), .clk (clk), .Q ({ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12205, new_AGEMA_signal_12201, new_AGEMA_signal_12197}), .clk (clk), .Q ({ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12217, new_AGEMA_signal_12213, new_AGEMA_signal_12209}), .clk (clk), .Q ({ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12229, new_AGEMA_signal_12225, new_AGEMA_signal_12221}), .clk (clk), .Q ({ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12241, new_AGEMA_signal_12237, new_AGEMA_signal_12233}), .clk (clk), .Q ({ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12253, new_AGEMA_signal_12249, new_AGEMA_signal_12245}), .clk (clk), .Q ({ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12265, new_AGEMA_signal_12261, new_AGEMA_signal_12257}), .clk (clk), .Q ({ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12277, new_AGEMA_signal_12273, new_AGEMA_signal_12269}), .clk (clk), .Q ({ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12289, new_AGEMA_signal_12285, new_AGEMA_signal_12281}), .clk (clk), .Q ({ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12301, new_AGEMA_signal_12297, new_AGEMA_signal_12293}), .clk (clk), .Q ({ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12313, new_AGEMA_signal_12309, new_AGEMA_signal_12305}), .clk (clk), .Q ({ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12325, new_AGEMA_signal_12321, new_AGEMA_signal_12317}), .clk (clk), .Q ({ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12337, new_AGEMA_signal_12333, new_AGEMA_signal_12329}), .clk (clk), .Q ({ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12349, new_AGEMA_signal_12345, new_AGEMA_signal_12341}), .clk (clk), .Q ({ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12361, new_AGEMA_signal_12357, new_AGEMA_signal_12353}), .clk (clk), .Q ({ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12373, new_AGEMA_signal_12369, new_AGEMA_signal_12365}), .clk (clk), .Q ({ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12385, new_AGEMA_signal_12381, new_AGEMA_signal_12377}), .clk (clk), .Q ({ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12397, new_AGEMA_signal_12393, new_AGEMA_signal_12389}), .clk (clk), .Q ({ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12409, new_AGEMA_signal_12405, new_AGEMA_signal_12401}), .clk (clk), .Q ({ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12421, new_AGEMA_signal_12417, new_AGEMA_signal_12413}), .clk (clk), .Q ({ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12433, new_AGEMA_signal_12429, new_AGEMA_signal_12425}), .clk (clk), .Q ({ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12445, new_AGEMA_signal_12441, new_AGEMA_signal_12437}), .clk (clk), .Q ({ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12457, new_AGEMA_signal_12453, new_AGEMA_signal_12449}), .clk (clk), .Q ({ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12469, new_AGEMA_signal_12465, new_AGEMA_signal_12461}), .clk (clk), .Q ({ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12481, new_AGEMA_signal_12477, new_AGEMA_signal_12473}), .clk (clk), .Q ({ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12493, new_AGEMA_signal_12489, new_AGEMA_signal_12485}), .clk (clk), .Q ({ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12505, new_AGEMA_signal_12501, new_AGEMA_signal_12497}), .clk (clk), .Q ({ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12517, new_AGEMA_signal_12513, new_AGEMA_signal_12509}), .clk (clk), .Q ({ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12529, new_AGEMA_signal_12525, new_AGEMA_signal_12521}), .clk (clk), .Q ({ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12541, new_AGEMA_signal_12537, new_AGEMA_signal_12533}), .clk (clk), .Q ({ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12553, new_AGEMA_signal_12549, new_AGEMA_signal_12545}), .clk (clk), .Q ({ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12565, new_AGEMA_signal_12561, new_AGEMA_signal_12557}), .clk (clk), .Q ({ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12577, new_AGEMA_signal_12573, new_AGEMA_signal_12569}), .clk (clk), .Q ({ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12589, new_AGEMA_signal_12585, new_AGEMA_signal_12581}), .clk (clk), .Q ({ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12601, new_AGEMA_signal_12597, new_AGEMA_signal_12593}), .clk (clk), .Q ({ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12613, new_AGEMA_signal_12609, new_AGEMA_signal_12605}), .clk (clk), .Q ({ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12625, new_AGEMA_signal_12621, new_AGEMA_signal_12617}), .clk (clk), .Q ({ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12637, new_AGEMA_signal_12633, new_AGEMA_signal_12629}), .clk (clk), .Q ({ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12649, new_AGEMA_signal_12645, new_AGEMA_signal_12641}), .clk (clk), .Q ({ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12661, new_AGEMA_signal_12657, new_AGEMA_signal_12653}), .clk (clk), .Q ({ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12673, new_AGEMA_signal_12669, new_AGEMA_signal_12665}), .clk (clk), .Q ({ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12685, new_AGEMA_signal_12681, new_AGEMA_signal_12677}), .clk (clk), .Q ({ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12697, new_AGEMA_signal_12693, new_AGEMA_signal_12689}), .clk (clk), .Q ({ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12709, new_AGEMA_signal_12705, new_AGEMA_signal_12701}), .clk (clk), .Q ({ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12721, new_AGEMA_signal_12717, new_AGEMA_signal_12713}), .clk (clk), .Q ({ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12733, new_AGEMA_signal_12729, new_AGEMA_signal_12725}), .clk (clk), .Q ({ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12745, new_AGEMA_signal_12741, new_AGEMA_signal_12737}), .clk (clk), .Q ({ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12757, new_AGEMA_signal_12753, new_AGEMA_signal_12749}), .clk (clk), .Q ({ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12769, new_AGEMA_signal_12765, new_AGEMA_signal_12761}), .clk (clk), .Q ({ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12781, new_AGEMA_signal_12777, new_AGEMA_signal_12773}), .clk (clk), .Q ({ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12793, new_AGEMA_signal_12789, new_AGEMA_signal_12785}), .clk (clk), .Q ({ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12805, new_AGEMA_signal_12801, new_AGEMA_signal_12797}), .clk (clk), .Q ({ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12817, new_AGEMA_signal_12813, new_AGEMA_signal_12809}), .clk (clk), .Q ({ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12829, new_AGEMA_signal_12825, new_AGEMA_signal_12821}), .clk (clk), .Q ({ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12841, new_AGEMA_signal_12837, new_AGEMA_signal_12833}), .clk (clk), .Q ({ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12853, new_AGEMA_signal_12849, new_AGEMA_signal_12845}), .clk (clk), .Q ({ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12865, new_AGEMA_signal_12861, new_AGEMA_signal_12857}), .clk (clk), .Q ({ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12877, new_AGEMA_signal_12873, new_AGEMA_signal_12869}), .clk (clk), .Q ({ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12889, new_AGEMA_signal_12885, new_AGEMA_signal_12881}), .clk (clk), .Q ({ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12901, new_AGEMA_signal_12897, new_AGEMA_signal_12893}), .clk (clk), .Q ({ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12913, new_AGEMA_signal_12909, new_AGEMA_signal_12905}), .clk (clk), .Q ({ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12925, new_AGEMA_signal_12921, new_AGEMA_signal_12917}), .clk (clk), .Q ({ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12937, new_AGEMA_signal_12933, new_AGEMA_signal_12929}), .clk (clk), .Q ({ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12949, new_AGEMA_signal_12945, new_AGEMA_signal_12941}), .clk (clk), .Q ({ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12961, new_AGEMA_signal_12957, new_AGEMA_signal_12953}), .clk (clk), .Q ({ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12973, new_AGEMA_signal_12969, new_AGEMA_signal_12965}), .clk (clk), .Q ({ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_12985, new_AGEMA_signal_12981, new_AGEMA_signal_12977}), .clk (clk), .Q ({ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, KeyReg_Inst_ff_SDE_0_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, KSSubBytesInput[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6079, new_AGEMA_signal_6078, KeyReg_Inst_ff_SDE_1_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, KSSubBytesInput[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6083, new_AGEMA_signal_6082, KeyReg_Inst_ff_SDE_2_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, KSSubBytesInput[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, KeyReg_Inst_ff_SDE_3_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, KSSubBytesInput[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6091, new_AGEMA_signal_6090, KeyReg_Inst_ff_SDE_4_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, KSSubBytesInput[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6095, new_AGEMA_signal_6094, KeyReg_Inst_ff_SDE_5_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, KSSubBytesInput[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, KeyReg_Inst_ff_SDE_6_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, KSSubBytesInput[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6103, new_AGEMA_signal_6102, KeyReg_Inst_ff_SDE_7_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KSSubBytesInput[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, KeyReg_Inst_ff_SDE_8_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KSSubBytesInput[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6107, new_AGEMA_signal_6106, KeyReg_Inst_ff_SDE_9_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, KSSubBytesInput[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, KeyReg_Inst_ff_SDE_10_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, KSSubBytesInput[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6115, new_AGEMA_signal_6114, KeyReg_Inst_ff_SDE_11_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, KSSubBytesInput[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6119, new_AGEMA_signal_6118, KeyReg_Inst_ff_SDE_12_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, KSSubBytesInput[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, KeyReg_Inst_ff_SDE_13_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, KSSubBytesInput[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6127, new_AGEMA_signal_6126, KeyReg_Inst_ff_SDE_14_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, KSSubBytesInput[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6131, new_AGEMA_signal_6130, KeyReg_Inst_ff_SDE_15_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, KSSubBytesInput[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyReg_Inst_ff_SDE_16_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, KSSubBytesInput[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, KeyReg_Inst_ff_SDE_17_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, KSSubBytesInput[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6139, new_AGEMA_signal_6138, KeyReg_Inst_ff_SDE_18_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, KSSubBytesInput[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6143, new_AGEMA_signal_6142, KeyReg_Inst_ff_SDE_19_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, KSSubBytesInput[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, KeyReg_Inst_ff_SDE_20_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, KSSubBytesInput[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6151, new_AGEMA_signal_6150, KeyReg_Inst_ff_SDE_21_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, KSSubBytesInput[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6155, new_AGEMA_signal_6154, KeyReg_Inst_ff_SDE_22_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, KSSubBytesInput[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, KeyReg_Inst_ff_SDE_23_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, KSSubBytesInput[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6163, new_AGEMA_signal_6162, KeyReg_Inst_ff_SDE_24_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, KSSubBytesInput[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6257, new_AGEMA_signal_6256, KeyReg_Inst_ff_SDE_25_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, KSSubBytesInput[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, KeyReg_Inst_ff_SDE_26_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, KSSubBytesInput[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6265, new_AGEMA_signal_6264, KeyReg_Inst_ff_SDE_27_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, KSSubBytesInput[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6269, new_AGEMA_signal_6268, KeyReg_Inst_ff_SDE_28_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, KSSubBytesInput[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, KeyReg_Inst_ff_SDE_29_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, KSSubBytesInput[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6277, new_AGEMA_signal_6276, KeyReg_Inst_ff_SDE_30_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, KSSubBytesInput[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6281, new_AGEMA_signal_6280, KeyReg_Inst_ff_SDE_31_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, KSSubBytesInput[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5461, new_AGEMA_signal_5460, KeyReg_Inst_ff_SDE_32_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, RoundKey[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, KeyReg_Inst_ff_SDE_33_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, RoundKey[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5791, new_AGEMA_signal_5790, KeyReg_Inst_ff_SDE_34_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, RoundKey[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyReg_Inst_ff_SDE_35_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, RoundKey[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, KeyReg_Inst_ff_SDE_36_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, RoundKey[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5803, new_AGEMA_signal_5802, KeyReg_Inst_ff_SDE_37_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, RoundKey[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyReg_Inst_ff_SDE_38_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, RoundKey[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, KeyReg_Inst_ff_SDE_39_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, RoundKey[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5465, new_AGEMA_signal_5464, KeyReg_Inst_ff_SDE_40_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, RoundKey[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5815, new_AGEMA_signal_5814, KeyReg_Inst_ff_SDE_41_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, RoundKey[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyReg_Inst_ff_SDE_42_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, RoundKey[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, KeyReg_Inst_ff_SDE_43_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, RoundKey[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5827, new_AGEMA_signal_5826, KeyReg_Inst_ff_SDE_44_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, RoundKey[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5831, new_AGEMA_signal_5830, KeyReg_Inst_ff_SDE_45_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, RoundKey[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, KeyReg_Inst_ff_SDE_46_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, RoundKey[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5839, new_AGEMA_signal_5838, KeyReg_Inst_ff_SDE_47_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, RoundKey[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, KeyReg_Inst_ff_SDE_48_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, RoundKey[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5843, new_AGEMA_signal_5842, KeyReg_Inst_ff_SDE_49_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, RoundKey[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, KeyReg_Inst_ff_SDE_50_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, RoundKey[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5851, new_AGEMA_signal_5850, KeyReg_Inst_ff_SDE_51_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, RoundKey[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5855, new_AGEMA_signal_5854, KeyReg_Inst_ff_SDE_52_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, RoundKey[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, KeyReg_Inst_ff_SDE_53_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, RoundKey[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5863, new_AGEMA_signal_5862, KeyReg_Inst_ff_SDE_54_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, RoundKey[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5867, new_AGEMA_signal_5866, KeyReg_Inst_ff_SDE_55_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, RoundKey[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, KeyReg_Inst_ff_SDE_56_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, RoundKey[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6167, new_AGEMA_signal_6166, KeyReg_Inst_ff_SDE_57_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, RoundKey[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, KeyReg_Inst_ff_SDE_58_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, RoundKey[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6175, new_AGEMA_signal_6174, KeyReg_Inst_ff_SDE_59_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, RoundKey[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6179, new_AGEMA_signal_6178, KeyReg_Inst_ff_SDE_60_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, RoundKey[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, KeyReg_Inst_ff_SDE_61_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, RoundKey[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6187, new_AGEMA_signal_6186, KeyReg_Inst_ff_SDE_62_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, RoundKey[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_6191, new_AGEMA_signal_6190, KeyReg_Inst_ff_SDE_63_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, RoundKey[63]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, KeyReg_Inst_ff_SDE_64_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, RoundKey[64]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5473, new_AGEMA_signal_5472, KeyReg_Inst_ff_SDE_65_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, RoundKey[65]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5477, new_AGEMA_signal_5476, KeyReg_Inst_ff_SDE_66_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, RoundKey[66]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, KeyReg_Inst_ff_SDE_67_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, RoundKey[67]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5485, new_AGEMA_signal_5484, KeyReg_Inst_ff_SDE_68_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, RoundKey[68]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5489, new_AGEMA_signal_5488, KeyReg_Inst_ff_SDE_69_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, RoundKey[69]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5493, new_AGEMA_signal_5492, KeyReg_Inst_ff_SDE_70_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, RoundKey[70]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5497, new_AGEMA_signal_5496, KeyReg_Inst_ff_SDE_71_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, RoundKey[71]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5173, new_AGEMA_signal_5172, KeyReg_Inst_ff_SDE_72_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, RoundKey[72]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5501, new_AGEMA_signal_5500, KeyReg_Inst_ff_SDE_73_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, RoundKey[73]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, KeyReg_Inst_ff_SDE_74_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, RoundKey[74]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5509, new_AGEMA_signal_5508, KeyReg_Inst_ff_SDE_75_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, RoundKey[75]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5513, new_AGEMA_signal_5512, KeyReg_Inst_ff_SDE_76_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, RoundKey[76]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, KeyReg_Inst_ff_SDE_77_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, RoundKey[77]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5521, new_AGEMA_signal_5520, KeyReg_Inst_ff_SDE_78_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, RoundKey[78]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5525, new_AGEMA_signal_5524, KeyReg_Inst_ff_SDE_79_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, RoundKey[79]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5177, new_AGEMA_signal_5176, KeyReg_Inst_ff_SDE_80_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, RoundKey[80]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, KeyReg_Inst_ff_SDE_81_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, RoundKey[81]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, KeyReg_Inst_ff_SDE_82_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, RoundKey[82]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5537, new_AGEMA_signal_5536, KeyReg_Inst_ff_SDE_83_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, RoundKey[83]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, KeyReg_Inst_ff_SDE_84_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, RoundKey[84]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, KeyReg_Inst_ff_SDE_85_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, RoundKey[85]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5549, new_AGEMA_signal_5548, KeyReg_Inst_ff_SDE_86_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, RoundKey[86]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, KeyReg_Inst_ff_SDE_87_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, RoundKey[87]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, KeyReg_Inst_ff_SDE_88_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, RoundKey[88]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5875, new_AGEMA_signal_5874, KeyReg_Inst_ff_SDE_89_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, RoundKey[89]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5879, new_AGEMA_signal_5878, KeyReg_Inst_ff_SDE_90_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, RoundKey[90]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, KeyReg_Inst_ff_SDE_91_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, RoundKey[91]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5887, new_AGEMA_signal_5886, KeyReg_Inst_ff_SDE_92_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, RoundKey[92]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5891, new_AGEMA_signal_5890, KeyReg_Inst_ff_SDE_93_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, RoundKey[93]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, KeyReg_Inst_ff_SDE_94_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, RoundKey[94]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5899, new_AGEMA_signal_5898, KeyReg_Inst_ff_SDE_95_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, RoundKey[95]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4979, new_AGEMA_signal_4978, KeyReg_Inst_ff_SDE_96_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, RoundKey[96]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, KeyReg_Inst_ff_SDE_97_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, RoundKey[97]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5185, new_AGEMA_signal_5184, KeyReg_Inst_ff_SDE_98_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, RoundKey[98]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5189, new_AGEMA_signal_5188, KeyReg_Inst_ff_SDE_99_next_state}), .clk (clk), .Q ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, RoundKey[99]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, KeyReg_Inst_ff_SDE_100_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, RoundKey[100]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5197, new_AGEMA_signal_5196, KeyReg_Inst_ff_SDE_101_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, RoundKey[101]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5201, new_AGEMA_signal_5200, KeyReg_Inst_ff_SDE_102_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2359, new_AGEMA_signal_2358, RoundKey[102]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5205, new_AGEMA_signal_5204, KeyReg_Inst_ff_SDE_103_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, RoundKey[103]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, KeyReg_Inst_ff_SDE_104_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2371, new_AGEMA_signal_2370, RoundKey[104]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5209, new_AGEMA_signal_5208, KeyReg_Inst_ff_SDE_105_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, RoundKey[105]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5213, new_AGEMA_signal_5212, KeyReg_Inst_ff_SDE_106_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, RoundKey[106]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, KeyReg_Inst_ff_SDE_107_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, RoundKey[107]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5221, new_AGEMA_signal_5220, KeyReg_Inst_ff_SDE_108_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, RoundKey[108]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5225, new_AGEMA_signal_5224, KeyReg_Inst_ff_SDE_109_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, RoundKey[109]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, KeyReg_Inst_ff_SDE_110_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, RoundKey[110]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5233, new_AGEMA_signal_5232, KeyReg_Inst_ff_SDE_111_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, RoundKey[111]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, KeyReg_Inst_ff_SDE_112_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, RoundKey[112]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5237, new_AGEMA_signal_5236, KeyReg_Inst_ff_SDE_113_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, RoundKey[113]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5241, new_AGEMA_signal_5240, KeyReg_Inst_ff_SDE_114_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, RoundKey[114]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5245, new_AGEMA_signal_5244, KeyReg_Inst_ff_SDE_115_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, RoundKey[115]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5249, new_AGEMA_signal_5248, KeyReg_Inst_ff_SDE_116_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, RoundKey[116]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, KeyReg_Inst_ff_SDE_117_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, RoundKey[117]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5257, new_AGEMA_signal_5256, KeyReg_Inst_ff_SDE_118_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, RoundKey[118]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5261, new_AGEMA_signal_5260, KeyReg_Inst_ff_SDE_119_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, RoundKey[119]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, KeyReg_Inst_ff_SDE_120_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, RoundKey[120]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5561, new_AGEMA_signal_5560, KeyReg_Inst_ff_SDE_121_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, RoundKey[121]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, KeyReg_Inst_ff_SDE_122_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, RoundKey[122]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, KeyReg_Inst_ff_SDE_123_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, RoundKey[123]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5573, new_AGEMA_signal_5572, KeyReg_Inst_ff_SDE_124_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, RoundKey[124]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, KeyReg_Inst_ff_SDE_125_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, RoundKey[125]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, KeyReg_Inst_ff_SDE_126_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, RoundKey[126]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_5585, new_AGEMA_signal_5584, KeyReg_Inst_ff_SDE_127_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D (new_AGEMA_signal_12989), .CK (clk), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D (new_AGEMA_signal_12993), .CK (clk), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D (new_AGEMA_signal_12997), .CK (clk), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D (new_AGEMA_signal_13001), .CK (clk), .Q (RoundCounter[3]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_0__FF_FF ( .D (new_AGEMA_signal_13005), .CK (clk), .Q (InRoundCounter[0]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_1__FF_FF ( .D (new_AGEMA_signal_13009), .CK (clk), .Q (InRoundCounter[1]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_2__FF_FF ( .D (new_AGEMA_signal_13013), .CK (clk), .Q (InRoundCounter[2]), .QN () ) ;
endmodule
