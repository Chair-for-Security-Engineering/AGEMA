////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module Midori64 in file /AGEMA/Designs/Midori_round_based/AGEMA/Midori64.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module Midori64_HPC3_Pipeline_d2 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, key_s2, DataIn_s1, DataIn_s2, Fresh, DataOut_s0, done, DataOut_s1, DataOut_s2);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [63:0] DataIn_s1 ;
    input [63:0] DataIn_s2 ;
    input [1535:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    output [63:0] DataOut_s2 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n12 ;
    wire controller_roundCounter_n11 ;
    wire controller_roundCounter_n10 ;
    wire controller_roundCounter_n9 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n7 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n3 ;
    wire controller_roundCounter_n2 ;
    wire controller_roundCounter_n1 ;
    wire controller_roundCounter_N10 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N8 ;
    wire controller_roundCounter_N7 ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_SelectedKey_0_ ;
    wire Midori_rounds_SelectedKey_1_ ;
    wire Midori_rounds_SelectedKey_2_ ;
    wire Midori_rounds_SelectedKey_3_ ;
    wire Midori_rounds_SelectedKey_4_ ;
    wire Midori_rounds_SelectedKey_5_ ;
    wire Midori_rounds_SelectedKey_6_ ;
    wire Midori_rounds_SelectedKey_7_ ;
    wire Midori_rounds_SelectedKey_8_ ;
    wire Midori_rounds_SelectedKey_9_ ;
    wire Midori_rounds_SelectedKey_10_ ;
    wire Midori_rounds_SelectedKey_11_ ;
    wire Midori_rounds_SelectedKey_12_ ;
    wire Midori_rounds_SelectedKey_13_ ;
    wire Midori_rounds_SelectedKey_14_ ;
    wire Midori_rounds_SelectedKey_15_ ;
    wire Midori_rounds_SelectedKey_16_ ;
    wire Midori_rounds_SelectedKey_17_ ;
    wire Midori_rounds_SelectedKey_18_ ;
    wire Midori_rounds_SelectedKey_19_ ;
    wire Midori_rounds_SelectedKey_20_ ;
    wire Midori_rounds_SelectedKey_21_ ;
    wire Midori_rounds_SelectedKey_22_ ;
    wire Midori_rounds_SelectedKey_23_ ;
    wire Midori_rounds_SelectedKey_24_ ;
    wire Midori_rounds_SelectedKey_25_ ;
    wire Midori_rounds_SelectedKey_26_ ;
    wire Midori_rounds_SelectedKey_27_ ;
    wire Midori_rounds_SelectedKey_28_ ;
    wire Midori_rounds_SelectedKey_29_ ;
    wire Midori_rounds_SelectedKey_30_ ;
    wire Midori_rounds_SelectedKey_31_ ;
    wire Midori_rounds_SelectedKey_32_ ;
    wire Midori_rounds_SelectedKey_33_ ;
    wire Midori_rounds_SelectedKey_34_ ;
    wire Midori_rounds_SelectedKey_35_ ;
    wire Midori_rounds_SelectedKey_36_ ;
    wire Midori_rounds_SelectedKey_37_ ;
    wire Midori_rounds_SelectedKey_38_ ;
    wire Midori_rounds_SelectedKey_39_ ;
    wire Midori_rounds_SelectedKey_40_ ;
    wire Midori_rounds_SelectedKey_41_ ;
    wire Midori_rounds_SelectedKey_42_ ;
    wire Midori_rounds_SelectedKey_43_ ;
    wire Midori_rounds_SelectedKey_44_ ;
    wire Midori_rounds_SelectedKey_45_ ;
    wire Midori_rounds_SelectedKey_46_ ;
    wire Midori_rounds_SelectedKey_47_ ;
    wire Midori_rounds_SelectedKey_48_ ;
    wire Midori_rounds_SelectedKey_49_ ;
    wire Midori_rounds_SelectedKey_50_ ;
    wire Midori_rounds_SelectedKey_51_ ;
    wire Midori_rounds_SelectedKey_52_ ;
    wire Midori_rounds_SelectedKey_53_ ;
    wire Midori_rounds_SelectedKey_54_ ;
    wire Midori_rounds_SelectedKey_55_ ;
    wire Midori_rounds_SelectedKey_56_ ;
    wire Midori_rounds_SelectedKey_57_ ;
    wire Midori_rounds_SelectedKey_58_ ;
    wire Midori_rounds_SelectedKey_59_ ;
    wire Midori_rounds_SelectedKey_60_ ;
    wire Midori_rounds_SelectedKey_61_ ;
    wire Midori_rounds_SelectedKey_62_ ;
    wire Midori_rounds_SelectedKey_63_ ;
    wire Midori_rounds_constant_MUX_n217 ;
    wire Midori_rounds_constant_MUX_n216 ;
    wire Midori_rounds_constant_MUX_n215 ;
    wire Midori_rounds_constant_MUX_n214 ;
    wire Midori_rounds_constant_MUX_n213 ;
    wire Midori_rounds_constant_MUX_n212 ;
    wire Midori_rounds_constant_MUX_n211 ;
    wire Midori_rounds_constant_MUX_n210 ;
    wire Midori_rounds_constant_MUX_n209 ;
    wire Midori_rounds_constant_MUX_n208 ;
    wire Midori_rounds_constant_MUX_n207 ;
    wire Midori_rounds_constant_MUX_n206 ;
    wire Midori_rounds_constant_MUX_n205 ;
    wire Midori_rounds_constant_MUX_n204 ;
    wire Midori_rounds_constant_MUX_n203 ;
    wire Midori_rounds_constant_MUX_n202 ;
    wire Midori_rounds_constant_MUX_n201 ;
    wire Midori_rounds_constant_MUX_n200 ;
    wire Midori_rounds_constant_MUX_n199 ;
    wire Midori_rounds_constant_MUX_n198 ;
    wire Midori_rounds_constant_MUX_n197 ;
    wire Midori_rounds_constant_MUX_n196 ;
    wire Midori_rounds_constant_MUX_n195 ;
    wire Midori_rounds_constant_MUX_n194 ;
    wire Midori_rounds_constant_MUX_n193 ;
    wire Midori_rounds_constant_MUX_n192 ;
    wire Midori_rounds_constant_MUX_n191 ;
    wire Midori_rounds_constant_MUX_n190 ;
    wire Midori_rounds_constant_MUX_n189 ;
    wire Midori_rounds_constant_MUX_n188 ;
    wire Midori_rounds_constant_MUX_n187 ;
    wire Midori_rounds_constant_MUX_n186 ;
    wire Midori_rounds_constant_MUX_n185 ;
    wire Midori_rounds_constant_MUX_n184 ;
    wire Midori_rounds_constant_MUX_n183 ;
    wire Midori_rounds_constant_MUX_n182 ;
    wire Midori_rounds_constant_MUX_n181 ;
    wire Midori_rounds_constant_MUX_n180 ;
    wire Midori_rounds_constant_MUX_n179 ;
    wire Midori_rounds_constant_MUX_n178 ;
    wire Midori_rounds_constant_MUX_n177 ;
    wire Midori_rounds_constant_MUX_n176 ;
    wire Midori_rounds_constant_MUX_n175 ;
    wire Midori_rounds_constant_MUX_n174 ;
    wire Midori_rounds_constant_MUX_n173 ;
    wire Midori_rounds_constant_MUX_n172 ;
    wire Midori_rounds_constant_MUX_n171 ;
    wire Midori_rounds_constant_MUX_n170 ;
    wire Midori_rounds_constant_MUX_n169 ;
    wire Midori_rounds_constant_MUX_n168 ;
    wire Midori_rounds_constant_MUX_n167 ;
    wire Midori_rounds_constant_MUX_n166 ;
    wire Midori_rounds_constant_MUX_n165 ;
    wire Midori_rounds_constant_MUX_n164 ;
    wire Midori_rounds_constant_MUX_n163 ;
    wire Midori_rounds_constant_MUX_n162 ;
    wire Midori_rounds_constant_MUX_n161 ;
    wire Midori_rounds_constant_MUX_n160 ;
    wire Midori_rounds_constant_MUX_n159 ;
    wire Midori_rounds_constant_MUX_n158 ;
    wire Midori_rounds_constant_MUX_n157 ;
    wire Midori_rounds_constant_MUX_n156 ;
    wire Midori_rounds_constant_MUX_n155 ;
    wire Midori_rounds_constant_MUX_n154 ;
    wire Midori_rounds_constant_MUX_n153 ;
    wire Midori_rounds_constant_MUX_n152 ;
    wire Midori_rounds_constant_MUX_n151 ;
    wire Midori_rounds_constant_MUX_n150 ;
    wire Midori_rounds_constant_MUX_n149 ;
    wire Midori_rounds_constant_MUX_n148 ;
    wire Midori_rounds_constant_MUX_n147 ;
    wire Midori_rounds_constant_MUX_n146 ;
    wire Midori_rounds_constant_MUX_n145 ;
    wire Midori_rounds_constant_MUX_n144 ;
    wire Midori_rounds_constant_MUX_n143 ;
    wire Midori_rounds_constant_MUX_n142 ;
    wire Midori_rounds_constant_MUX_n141 ;
    wire Midori_rounds_constant_MUX_n140 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n135 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_MUXInst_n11 ;
    wire Midori_rounds_MUXInst_n10 ;
    wire Midori_rounds_MUXInst_n9 ;
    wire Midori_rounds_MUXInst_n8 ;
    wire Midori_rounds_roundResult_Reg_SFF_0_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_1_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_2_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_3_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_4_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_5_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_6_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_7_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_8_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_9_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_10_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_11_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_12_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_13_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_14_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_15_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_16_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_17_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_18_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_19_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_20_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_21_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_22_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_23_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_24_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_25_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_26_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_27_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_28_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_29_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_30_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_31_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_32_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_33_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_34_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_35_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_36_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_37_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_38_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_39_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_40_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_41_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_42_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_43_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_44_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_45_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_46_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_47_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_48_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_49_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_50_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_51_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_52_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_53_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_54_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_55_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_56_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_57_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_58_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_59_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_60_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_61_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_62_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_63_DQ ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [15:0] Midori_rounds_round_Constant ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;

    /* cells in depth 0 */
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U64 ( .a ({key_s2[73], key_s1[73], key_s0[73]}), .b ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U63 ( .a ({key_s2[72], key_s1[72], key_s0[72]}), .b ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U62 ( .a ({key_s2[71], key_s1[71], key_s0[71]}), .b ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U61 ( .a ({key_s2[6], key_s1[6], key_s0[6]}), .b ({key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U60 ( .a ({key_s2[127], key_s1[127], key_s0[127]}), .b ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U59 ( .a ({key_s2[126], key_s1[126], key_s0[126]}), .b ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U58 ( .a ({key_s2[125], key_s1[125], key_s0[125]}), .b ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U57 ( .a ({key_s2[124], key_s1[124], key_s0[124]}), .b ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U56 ( .a ({key_s2[5], key_s1[5], key_s0[5]}), .b ({key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U55 ( .a ({key_s2[123], key_s1[123], key_s0[123]}), .b ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U54 ( .a ({key_s2[122], key_s1[122], key_s0[122]}), .b ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U53 ( .a ({key_s2[121], key_s1[121], key_s0[121]}), .b ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U52 ( .a ({key_s2[120], key_s1[120], key_s0[120]}), .b ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U51 ( .a ({key_s2[119], key_s1[119], key_s0[119]}), .b ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U50 ( .a ({key_s2[118], key_s1[118], key_s0[118]}), .b ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U49 ( .a ({key_s2[117], key_s1[117], key_s0[117]}), .b ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U48 ( .a ({key_s2[116], key_s1[116], key_s0[116]}), .b ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U47 ( .a ({key_s2[115], key_s1[115], key_s0[115]}), .b ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U46 ( .a ({key_s2[114], key_s1[114], key_s0[114]}), .b ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U45 ( .a ({key_s2[4], key_s1[4], key_s0[4]}), .b ({key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U44 ( .a ({key_s2[113], key_s1[113], key_s0[113]}), .b ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U43 ( .a ({key_s2[112], key_s1[112], key_s0[112]}), .b ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U42 ( .a ({key_s2[111], key_s1[111], key_s0[111]}), .b ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U41 ( .a ({key_s2[110], key_s1[110], key_s0[110]}), .b ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U40 ( .a ({key_s2[109], key_s1[109], key_s0[109]}), .b ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U39 ( .a ({key_s2[108], key_s1[108], key_s0[108]}), .b ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U38 ( .a ({key_s2[107], key_s1[107], key_s0[107]}), .b ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U37 ( .a ({key_s2[106], key_s1[106], key_s0[106]}), .b ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U36 ( .a ({key_s2[105], key_s1[105], key_s0[105]}), .b ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U35 ( .a ({key_s2[104], key_s1[104], key_s0[104]}), .b ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U34 ( .a ({key_s2[3], key_s1[3], key_s0[3]}), .b ({key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U33 ( .a ({key_s2[103], key_s1[103], key_s0[103]}), .b ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U32 ( .a ({key_s2[102], key_s1[102], key_s0[102]}), .b ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U31 ( .a ({key_s2[101], key_s1[101], key_s0[101]}), .b ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U30 ( .a ({key_s2[100], key_s1[100], key_s0[100]}), .b ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U29 ( .a ({key_s2[35], key_s1[35], key_s0[35]}), .b ({key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U28 ( .a ({key_s2[34], key_s1[34], key_s0[34]}), .b ({key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U27 ( .a ({key_s2[33], key_s1[33], key_s0[33]}), .b ({key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U26 ( .a ({key_s2[32], key_s1[32], key_s0[32]}), .b ({key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U25 ( .a ({key_s2[31], key_s1[31], key_s0[31]}), .b ({key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U24 ( .a ({key_s2[30], key_s1[30], key_s0[30]}), .b ({key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U23 ( .a ({key_s2[2], key_s1[2], key_s0[2]}), .b ({key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U22 ( .a ({key_s2[29], key_s1[29], key_s0[29]}), .b ({key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U21 ( .a ({key_s2[28], key_s1[28], key_s0[28]}), .b ({key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U20 ( .a ({key_s2[27], key_s1[27], key_s0[27]}), .b ({key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U19 ( .a ({key_s2[26], key_s1[26], key_s0[26]}), .b ({key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U18 ( .a ({key_s2[25], key_s1[25], key_s0[25]}), .b ({key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U17 ( .a ({key_s2[24], key_s1[24], key_s0[24]}), .b ({key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U16 ( .a ({key_s2[23], key_s1[23], key_s0[23]}), .b ({key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U15 ( .a ({key_s2[22], key_s1[22], key_s0[22]}), .b ({key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U14 ( .a ({key_s2[21], key_s1[21], key_s0[21]}), .b ({key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U13 ( .a ({key_s2[20], key_s1[20], key_s0[20]}), .b ({key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U12 ( .a ({key_s2[1], key_s1[1], key_s0[1]}), .b ({key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U11 ( .a ({key_s2[19], key_s1[19], key_s0[19]}), .b ({key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U10 ( .a ({key_s2[18], key_s1[18], key_s0[18]}), .b ({key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U9 ( .a ({key_s2[17], key_s1[17], key_s0[17]}), .b ({key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U8 ( .a ({key_s2[16], key_s1[16], key_s0[16]}), .b ({key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U7 ( .a ({key_s2[15], key_s1[15], key_s0[15]}), .b ({key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U6 ( .a ({key_s2[14], key_s1[14], key_s0[14]}), .b ({key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U5 ( .a ({key_s2[13], key_s1[13], key_s0[13]}), .b ({key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U4 ( .a ({key_s2[12], key_s1[12], key_s0[12]}), .b ({key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U3 ( .a ({key_s2[11], key_s1[11], key_s0[11]}), .b ({key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U2 ( .a ({key_s2[10], key_s1[10], key_s0[10]}), .b ({key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) keys_U1 ( .a ({key_s2[0], key_s1[0], key_s0[0]}), .b ({key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}) ) ;
    NOR2_X1 controller_U3 ( .A1 (controller_n2), .A2 (controller_n1), .ZN (new_AGEMA_signal_5520) ) ;
    NAND2_X1 controller_U2 ( .A1 (round_Signal[0]), .A2 (round_Signal[1]), .ZN (controller_n1) ) ;
    NAND2_X1 controller_U1 ( .A1 (round_Signal[2]), .A2 (round_Signal[3]), .ZN (controller_n2) ) ;
    INV_X1 controller_roundCounter_U14 ( .A (controller_roundCounter_n13), .ZN (controller_roundCounter_n2) ) ;
    MUX2_X1 controller_roundCounter_U13 ( .S (controller_roundCounter_n6), .A (controller_roundCounter_n12), .B (controller_roundCounter_n11), .Z (controller_roundCounter_n13) ) ;
    NOR2_X1 controller_roundCounter_U12 ( .A1 (reset), .A2 (controller_roundCounter_n10), .ZN (controller_roundCounter_N8) ) ;
    XNOR2_X1 controller_roundCounter_U11 ( .A (round_Signal[0]), .B (round_Signal[1]), .ZN (controller_roundCounter_n10) ) ;
    MUX2_X1 controller_roundCounter_U10 ( .S (round_Signal[3]), .A (controller_roundCounter_n9), .B (controller_roundCounter_n8), .Z (controller_roundCounter_N10) ) ;
    NAND2_X1 controller_roundCounter_U9 ( .A1 (controller_roundCounter_n12), .A2 (controller_roundCounter_n7), .ZN (controller_roundCounter_n8) ) ;
    NAND2_X1 controller_roundCounter_U8 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n3), .ZN (controller_roundCounter_n7) ) ;
    NOR2_X1 controller_roundCounter_U7 ( .A1 (controller_roundCounter_n5), .A2 (controller_roundCounter_N7), .ZN (controller_roundCounter_n12) ) ;
    NOR2_X1 controller_roundCounter_U6 ( .A1 (round_Signal[1]), .A2 (reset), .ZN (controller_roundCounter_n5) ) ;
    NOR2_X1 controller_roundCounter_U5 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n11), .ZN (controller_roundCounter_n9) ) ;
    NAND2_X1 controller_roundCounter_U4 ( .A1 (round_Signal[1]), .A2 (controller_roundCounter_n4), .ZN (controller_roundCounter_n11) ) ;
    NOR2_X1 controller_roundCounter_U3 ( .A1 (reset), .A2 (controller_roundCounter_n1), .ZN (controller_roundCounter_n4) ) ;
    NOR2_X1 controller_roundCounter_U2 ( .A1 (reset), .A2 (round_Signal[0]), .ZN (controller_roundCounter_N7) ) ;
    INV_X1 controller_roundCounter_U1 ( .A (reset), .ZN (controller_roundCounter_n3) ) ;
    INV_X1 controller_roundCounter_count_reg_0__U1 ( .A (round_Signal[0]), .ZN (controller_roundCounter_n1) ) ;
    INV_X1 controller_roundCounter_count_reg_2__U1 ( .A (round_Signal[2]), .ZN (controller_roundCounter_n6) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U64 ( .a ({new_AGEMA_signal_1461, new_AGEMA_signal_1460, wk[9]}), .b ({DataIn_s2[9], DataIn_s1[9], DataIn_s0[9]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, Midori_add_Result_Start[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U63 ( .a ({new_AGEMA_signal_1467, new_AGEMA_signal_1466, wk[8]}), .b ({DataIn_s2[8], DataIn_s1[8], DataIn_s0[8]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, Midori_add_Result_Start[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U62 ( .a ({new_AGEMA_signal_1473, new_AGEMA_signal_1472, wk[7]}), .b ({DataIn_s2[7], DataIn_s1[7], DataIn_s0[7]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, Midori_add_Result_Start[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U61 ( .a ({new_AGEMA_signal_1479, new_AGEMA_signal_1478, wk[6]}), .b ({DataIn_s2[6], DataIn_s1[6], DataIn_s0[6]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, Midori_add_Result_Start[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U60 ( .a ({new_AGEMA_signal_1485, new_AGEMA_signal_1484, wk[63]}), .b ({DataIn_s2[63], DataIn_s1[63], DataIn_s0[63]}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, Midori_add_Result_Start[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U59 ( .a ({new_AGEMA_signal_1491, new_AGEMA_signal_1490, wk[62]}), .b ({DataIn_s2[62], DataIn_s1[62], DataIn_s0[62]}), .c ({new_AGEMA_signal_2145, new_AGEMA_signal_2144, Midori_add_Result_Start[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U58 ( .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496, wk[61]}), .b ({DataIn_s2[61], DataIn_s1[61], DataIn_s0[61]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, Midori_add_Result_Start[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U57 ( .a ({new_AGEMA_signal_1503, new_AGEMA_signal_1502, wk[60]}), .b ({DataIn_s2[60], DataIn_s1[60], DataIn_s0[60]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, Midori_add_Result_Start[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U56 ( .a ({new_AGEMA_signal_1509, new_AGEMA_signal_1508, wk[5]}), .b ({DataIn_s2[5], DataIn_s1[5], DataIn_s0[5]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, Midori_add_Result_Start[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U55 ( .a ({new_AGEMA_signal_1515, new_AGEMA_signal_1514, wk[59]}), .b ({DataIn_s2[59], DataIn_s1[59], DataIn_s0[59]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, Midori_add_Result_Start[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U54 ( .a ({new_AGEMA_signal_1521, new_AGEMA_signal_1520, wk[58]}), .b ({DataIn_s2[58], DataIn_s1[58], DataIn_s0[58]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, Midori_add_Result_Start[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U53 ( .a ({new_AGEMA_signal_1527, new_AGEMA_signal_1526, wk[57]}), .b ({DataIn_s2[57], DataIn_s1[57], DataIn_s0[57]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, Midori_add_Result_Start[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U52 ( .a ({new_AGEMA_signal_1533, new_AGEMA_signal_1532, wk[56]}), .b ({DataIn_s2[56], DataIn_s1[56], DataIn_s0[56]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, Midori_add_Result_Start[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U51 ( .a ({new_AGEMA_signal_1539, new_AGEMA_signal_1538, wk[55]}), .b ({DataIn_s2[55], DataIn_s1[55], DataIn_s0[55]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, Midori_add_Result_Start[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U50 ( .a ({new_AGEMA_signal_1545, new_AGEMA_signal_1544, wk[54]}), .b ({DataIn_s2[54], DataIn_s1[54], DataIn_s0[54]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, Midori_add_Result_Start[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U49 ( .a ({new_AGEMA_signal_1551, new_AGEMA_signal_1550, wk[53]}), .b ({DataIn_s2[53], DataIn_s1[53], DataIn_s0[53]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, Midori_add_Result_Start[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U48 ( .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1556, wk[52]}), .b ({DataIn_s2[52], DataIn_s1[52], DataIn_s0[52]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, Midori_add_Result_Start[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U47 ( .a ({new_AGEMA_signal_1563, new_AGEMA_signal_1562, wk[51]}), .b ({DataIn_s2[51], DataIn_s1[51], DataIn_s0[51]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, Midori_add_Result_Start[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U46 ( .a ({new_AGEMA_signal_1569, new_AGEMA_signal_1568, wk[50]}), .b ({DataIn_s2[50], DataIn_s1[50], DataIn_s0[50]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, Midori_add_Result_Start[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U45 ( .a ({new_AGEMA_signal_1575, new_AGEMA_signal_1574, wk[4]}), .b ({DataIn_s2[4], DataIn_s1[4], DataIn_s0[4]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, Midori_add_Result_Start[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U44 ( .a ({new_AGEMA_signal_1581, new_AGEMA_signal_1580, wk[49]}), .b ({DataIn_s2[49], DataIn_s1[49], DataIn_s0[49]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, Midori_add_Result_Start[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U43 ( .a ({new_AGEMA_signal_1587, new_AGEMA_signal_1586, wk[48]}), .b ({DataIn_s2[48], DataIn_s1[48], DataIn_s0[48]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, Midori_add_Result_Start[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U42 ( .a ({new_AGEMA_signal_1593, new_AGEMA_signal_1592, wk[47]}), .b ({DataIn_s2[47], DataIn_s1[47], DataIn_s0[47]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, Midori_add_Result_Start[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U41 ( .a ({new_AGEMA_signal_1599, new_AGEMA_signal_1598, wk[46]}), .b ({DataIn_s2[46], DataIn_s1[46], DataIn_s0[46]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, Midori_add_Result_Start[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U40 ( .a ({new_AGEMA_signal_1605, new_AGEMA_signal_1604, wk[45]}), .b ({DataIn_s2[45], DataIn_s1[45], DataIn_s0[45]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, Midori_add_Result_Start[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U39 ( .a ({new_AGEMA_signal_1611, new_AGEMA_signal_1610, wk[44]}), .b ({DataIn_s2[44], DataIn_s1[44], DataIn_s0[44]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, Midori_add_Result_Start[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U38 ( .a ({new_AGEMA_signal_1617, new_AGEMA_signal_1616, wk[43]}), .b ({DataIn_s2[43], DataIn_s1[43], DataIn_s0[43]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, Midori_add_Result_Start[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U37 ( .a ({new_AGEMA_signal_1623, new_AGEMA_signal_1622, wk[42]}), .b ({DataIn_s2[42], DataIn_s1[42], DataIn_s0[42]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, Midori_add_Result_Start[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U36 ( .a ({new_AGEMA_signal_1629, new_AGEMA_signal_1628, wk[41]}), .b ({DataIn_s2[41], DataIn_s1[41], DataIn_s0[41]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, Midori_add_Result_Start[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U35 ( .a ({new_AGEMA_signal_1635, new_AGEMA_signal_1634, wk[40]}), .b ({DataIn_s2[40], DataIn_s1[40], DataIn_s0[40]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, Midori_add_Result_Start[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U34 ( .a ({new_AGEMA_signal_1641, new_AGEMA_signal_1640, wk[3]}), .b ({DataIn_s2[3], DataIn_s1[3], DataIn_s0[3]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, Midori_add_Result_Start[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U33 ( .a ({new_AGEMA_signal_1647, new_AGEMA_signal_1646, wk[39]}), .b ({DataIn_s2[39], DataIn_s1[39], DataIn_s0[39]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, Midori_add_Result_Start[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U32 ( .a ({new_AGEMA_signal_1653, new_AGEMA_signal_1652, wk[38]}), .b ({DataIn_s2[38], DataIn_s1[38], DataIn_s0[38]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, Midori_add_Result_Start[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U31 ( .a ({new_AGEMA_signal_1659, new_AGEMA_signal_1658, wk[37]}), .b ({DataIn_s2[37], DataIn_s1[37], DataIn_s0[37]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, Midori_add_Result_Start[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U30 ( .a ({new_AGEMA_signal_1665, new_AGEMA_signal_1664, wk[36]}), .b ({DataIn_s2[36], DataIn_s1[36], DataIn_s0[36]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, Midori_add_Result_Start[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U29 ( .a ({new_AGEMA_signal_1671, new_AGEMA_signal_1670, wk[35]}), .b ({DataIn_s2[35], DataIn_s1[35], DataIn_s0[35]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, Midori_add_Result_Start[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U28 ( .a ({new_AGEMA_signal_1677, new_AGEMA_signal_1676, wk[34]}), .b ({DataIn_s2[34], DataIn_s1[34], DataIn_s0[34]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, Midori_add_Result_Start[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U27 ( .a ({new_AGEMA_signal_1683, new_AGEMA_signal_1682, wk[33]}), .b ({DataIn_s2[33], DataIn_s1[33], DataIn_s0[33]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, Midori_add_Result_Start[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U26 ( .a ({new_AGEMA_signal_1689, new_AGEMA_signal_1688, wk[32]}), .b ({DataIn_s2[32], DataIn_s1[32], DataIn_s0[32]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, Midori_add_Result_Start[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U25 ( .a ({new_AGEMA_signal_1695, new_AGEMA_signal_1694, wk[31]}), .b ({DataIn_s2[31], DataIn_s1[31], DataIn_s0[31]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, Midori_add_Result_Start[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U24 ( .a ({new_AGEMA_signal_1701, new_AGEMA_signal_1700, wk[30]}), .b ({DataIn_s2[30], DataIn_s1[30], DataIn_s0[30]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, Midori_add_Result_Start[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U23 ( .a ({new_AGEMA_signal_1707, new_AGEMA_signal_1706, wk[2]}), .b ({DataIn_s2[2], DataIn_s1[2], DataIn_s0[2]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, Midori_add_Result_Start[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U22 ( .a ({new_AGEMA_signal_1713, new_AGEMA_signal_1712, wk[29]}), .b ({DataIn_s2[29], DataIn_s1[29], DataIn_s0[29]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, Midori_add_Result_Start[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U21 ( .a ({new_AGEMA_signal_1719, new_AGEMA_signal_1718, wk[28]}), .b ({DataIn_s2[28], DataIn_s1[28], DataIn_s0[28]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, Midori_add_Result_Start[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U20 ( .a ({new_AGEMA_signal_1725, new_AGEMA_signal_1724, wk[27]}), .b ({DataIn_s2[27], DataIn_s1[27], DataIn_s0[27]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, Midori_add_Result_Start[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U19 ( .a ({new_AGEMA_signal_1731, new_AGEMA_signal_1730, wk[26]}), .b ({DataIn_s2[26], DataIn_s1[26], DataIn_s0[26]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, Midori_add_Result_Start[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U18 ( .a ({new_AGEMA_signal_1737, new_AGEMA_signal_1736, wk[25]}), .b ({DataIn_s2[25], DataIn_s1[25], DataIn_s0[25]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, Midori_add_Result_Start[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U17 ( .a ({new_AGEMA_signal_1743, new_AGEMA_signal_1742, wk[24]}), .b ({DataIn_s2[24], DataIn_s1[24], DataIn_s0[24]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, Midori_add_Result_Start[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U16 ( .a ({new_AGEMA_signal_1749, new_AGEMA_signal_1748, wk[23]}), .b ({DataIn_s2[23], DataIn_s1[23], DataIn_s0[23]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, Midori_add_Result_Start[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U15 ( .a ({new_AGEMA_signal_1755, new_AGEMA_signal_1754, wk[22]}), .b ({DataIn_s2[22], DataIn_s1[22], DataIn_s0[22]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, Midori_add_Result_Start[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U14 ( .a ({new_AGEMA_signal_1761, new_AGEMA_signal_1760, wk[21]}), .b ({DataIn_s2[21], DataIn_s1[21], DataIn_s0[21]}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, Midori_add_Result_Start[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U13 ( .a ({new_AGEMA_signal_1767, new_AGEMA_signal_1766, wk[20]}), .b ({DataIn_s2[20], DataIn_s1[20], DataIn_s0[20]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, Midori_add_Result_Start[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U12 ( .a ({new_AGEMA_signal_1773, new_AGEMA_signal_1772, wk[1]}), .b ({DataIn_s2[1], DataIn_s1[1], DataIn_s0[1]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, Midori_add_Result_Start[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U11 ( .a ({new_AGEMA_signal_1779, new_AGEMA_signal_1778, wk[19]}), .b ({DataIn_s2[19], DataIn_s1[19], DataIn_s0[19]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, Midori_add_Result_Start[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U10 ( .a ({new_AGEMA_signal_1785, new_AGEMA_signal_1784, wk[18]}), .b ({DataIn_s2[18], DataIn_s1[18], DataIn_s0[18]}), .c ({new_AGEMA_signal_2341, new_AGEMA_signal_2340, Midori_add_Result_Start[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U9 ( .a ({new_AGEMA_signal_1791, new_AGEMA_signal_1790, wk[17]}), .b ({DataIn_s2[17], DataIn_s1[17], DataIn_s0[17]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, Midori_add_Result_Start[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U8 ( .a ({new_AGEMA_signal_1797, new_AGEMA_signal_1796, wk[16]}), .b ({DataIn_s2[16], DataIn_s1[16], DataIn_s0[16]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, Midori_add_Result_Start[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U7 ( .a ({new_AGEMA_signal_1803, new_AGEMA_signal_1802, wk[15]}), .b ({DataIn_s2[15], DataIn_s1[15], DataIn_s0[15]}), .c ({new_AGEMA_signal_2353, new_AGEMA_signal_2352, Midori_add_Result_Start[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U6 ( .a ({new_AGEMA_signal_1809, new_AGEMA_signal_1808, wk[14]}), .b ({DataIn_s2[14], DataIn_s1[14], DataIn_s0[14]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, Midori_add_Result_Start[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U5 ( .a ({new_AGEMA_signal_1815, new_AGEMA_signal_1814, wk[13]}), .b ({DataIn_s2[13], DataIn_s1[13], DataIn_s0[13]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, Midori_add_Result_Start[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U4 ( .a ({new_AGEMA_signal_1821, new_AGEMA_signal_1820, wk[12]}), .b ({DataIn_s2[12], DataIn_s1[12], DataIn_s0[12]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, Midori_add_Result_Start[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U3 ( .a ({new_AGEMA_signal_1827, new_AGEMA_signal_1826, wk[11]}), .b ({DataIn_s2[11], DataIn_s1[11], DataIn_s0[11]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, Midori_add_Result_Start[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U2 ( .a ({new_AGEMA_signal_1833, new_AGEMA_signal_1832, wk[10]}), .b ({DataIn_s2[10], DataIn_s1[10], DataIn_s0[10]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, Midori_add_Result_Start[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U1 ( .a ({new_AGEMA_signal_1839, new_AGEMA_signal_1838, wk[0]}), .b ({DataIn_s2[0], DataIn_s1[0], DataIn_s0[0]}), .c ({new_AGEMA_signal_2377, new_AGEMA_signal_2376, Midori_add_Result_Start[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U78 ( .a ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, Midori_rounds_SelectedKey_8_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[2]}), .c ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, Midori_rounds_n16}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U71 ( .a ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, Midori_rounds_SelectedKey_60_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[15]}), .c ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, Midori_rounds_n15}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U65 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_rounds_SelectedKey_56_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[14]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, Midori_rounds_n14}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U60 ( .a ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, Midori_rounds_SelectedKey_52_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[13]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, Midori_rounds_n13}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U56 ( .a ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, Midori_rounds_SelectedKey_4_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[1]}), .c ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, Midori_rounds_n12}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U53 ( .a ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, Midori_rounds_SelectedKey_48_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[12]}), .c ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, Midori_rounds_n11}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U48 ( .a ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_rounds_SelectedKey_44_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[11]}), .c ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, Midori_rounds_n10}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U43 ( .a ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, Midori_rounds_SelectedKey_40_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[10]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, Midori_rounds_n9}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U37 ( .a ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, Midori_rounds_SelectedKey_36_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[9]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, Midori_rounds_n8}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U32 ( .a ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_rounds_SelectedKey_32_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[8]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, Midori_rounds_n7}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U26 ( .a ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, Midori_rounds_SelectedKey_28_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[7]}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, Midori_rounds_n6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U21 ( .a ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, Midori_rounds_SelectedKey_24_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[6]}), .c ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, Midori_rounds_n5}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U16 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, Midori_rounds_SelectedKey_20_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[5]}), .c ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, Midori_rounds_n4}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U10 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_rounds_SelectedKey_16_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[4]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, Midori_rounds_n3}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U5 ( .a ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, Midori_rounds_SelectedKey_12_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[3]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, Midori_rounds_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U1 ( .a ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, Midori_rounds_SelectedKey_0_}), .b ({1'b0, 1'b0, Midori_rounds_round_Constant[0]}), .c ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, Midori_rounds_n1}) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U106 ( .A1 (Midori_rounds_constant_MUX_n217), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_round_Constant[9]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U105 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n214), .ZN (Midori_rounds_constant_MUX_n217) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U104 ( .A1 (Midori_rounds_constant_MUX_n213), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n214) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U103 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_round_Constant[8]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U102 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n208), .ZN (Midori_rounds_round_Constant[7]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U101 ( .A1 (Midori_rounds_round_Constant[11]), .A2 (Midori_rounds_constant_MUX_n207), .ZN (Midori_rounds_constant_MUX_n208) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U100 ( .A1 (Midori_rounds_constant_MUX_n206), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n207) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U99 ( .A1 (Midori_rounds_constant_MUX_n204), .A2 (Midori_rounds_constant_MUX_n203), .ZN (Midori_rounds_constant_MUX_n206) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U98 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n201), .ZN (Midori_rounds_round_Constant[6]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U97 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n199), .ZN (Midori_rounds_constant_MUX_n201) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U96 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n197), .ZN (Midori_rounds_round_Constant[5]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U95 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n196), .ZN (Midori_rounds_constant_MUX_n197) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U94 ( .A1 (Midori_rounds_constant_MUX_n195), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n196) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U93 ( .A1 (Midori_rounds_constant_MUX_n194), .A2 (Midori_rounds_constant_MUX_n195), .ZN (Midori_rounds_round_Constant[4]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U92 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n195) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U91 ( .A1 (Midori_rounds_constant_MUX_n191), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[3]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U90 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n189), .ZN (Midori_rounds_constant_MUX_n191) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U89 ( .A1 (Midori_rounds_constant_MUX_n188), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n189) ) ;
    INV_X1 Midori_rounds_constant_MUX_U88 ( .A (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n188) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U87 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n186), .ZN (Midori_rounds_round_Constant[2]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U86 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n185), .ZN (Midori_rounds_constant_MUX_n186) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U85 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n202) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U84 ( .A1 (Midori_rounds_constant_MUX_n183), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n215) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U83 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n181), .ZN (Midori_rounds_round_Constant[1]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U82 ( .A1 (Midori_rounds_constant_MUX_n187), .A2 (Midori_rounds_constant_MUX_n180), .ZN (Midori_rounds_constant_MUX_n181) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U81 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n204), .ZN (Midori_rounds_constant_MUX_n180) ) ;
    INV_X1 Midori_rounds_constant_MUX_U80 ( .A (Midori_rounds_constant_MUX_n183), .ZN (Midori_rounds_constant_MUX_n204) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U79 ( .A1 (Midori_rounds_constant_MUX_n179), .A2 (Midori_rounds_constant_MUX_n178), .ZN (Midori_rounds_constant_MUX_n183) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U78 ( .A1 (Midori_rounds_constant_MUX_n177), .A2 (Midori_rounds_constant_MUX_n176), .ZN (Midori_rounds_constant_MUX_n178) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U77 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n175), .ZN (Midori_rounds_constant_MUX_n212) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U76 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n173), .Z (Midori_rounds_constant_MUX_n175) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U75 ( .A1 (Midori_rounds_constant_MUX_n172), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[15]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U74 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n172) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U73 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n194), .ZN (Midori_rounds_round_Constant[14]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U72 ( .A1 (Midori_rounds_constant_MUX_n169), .A2 (Midori_rounds_constant_MUX_n168), .ZN (Midori_rounds_constant_MUX_n194) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U71 ( .A1 (Midori_rounds_constant_MUX_n216), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n168) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U70 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n167), .ZN (Midori_rounds_constant_MUX_n205) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U69 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n167) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U68 ( .A1 (Midori_rounds_constant_MUX_n185), .A2 (Midori_rounds_constant_MUX_n164), .ZN (Midori_rounds_round_Constant[13]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U67 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n162), .ZN (Midori_rounds_constant_MUX_n164) ) ;
    INV_X1 Midori_rounds_constant_MUX_U66 ( .A (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n162) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U65 ( .A1 (Midori_rounds_constant_MUX_n161), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n185) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U64 ( .A1 (Midori_rounds_constant_MUX_n160), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[12]) ) ;
    INV_X1 Midori_rounds_constant_MUX_U63 ( .A (Midori_rounds_constant_MUX_n184), .ZN (Midori_rounds_constant_MUX_n190) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U62 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n159), .ZN (Midori_rounds_constant_MUX_n160) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U61 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n159) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U60 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n169), .ZN (Midori_rounds_constant_MUX_n211) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U59 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n158), .ZN (Midori_rounds_constant_MUX_n169) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U58 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n157), .ZN (Midori_rounds_constant_MUX_n158) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U57 ( .A1 (Midori_rounds_constant_MUX_n165), .A2 (Midori_rounds_constant_MUX_n177), .ZN (Midori_rounds_constant_MUX_n157) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U56 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n156), .ZN (Midori_rounds_constant_MUX_n198) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U55 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n155), .ZN (Midori_rounds_constant_MUX_n156) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U54 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n176), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n155) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U53 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n154), .ZN (Midori_rounds_constant_MUX_n200) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U52 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n154) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U51 ( .A1 (Midori_rounds_constant_MUX_n199), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_round_Constant[11]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U50 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n199) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U49 ( .A1 (Midori_rounds_constant_MUX_n152), .A2 (Midori_rounds_constant_MUX_n151), .ZN (Midori_rounds_constant_MUX_n210) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U48 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n151) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U47 ( .A1 (Midori_rounds_constant_MUX_n150), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n170) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U46 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n149), .ZN (Midori_rounds_constant_MUX_n187) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U45 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n149) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U44 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n148), .ZN (Midori_rounds_constant_MUX_n150) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U43 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n148) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U42 ( .A1 (Midori_rounds_constant_MUX_n147), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[10]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U41 ( .A1 (Midori_rounds_constant_MUX_n146), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_constant_MUX_n171) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U40 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n145), .ZN (Midori_rounds_constant_MUX_n213) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U39 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n177), .Z (Midori_rounds_constant_MUX_n145) ) ;
    INV_X1 Midori_rounds_constant_MUX_U38 ( .A (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_constant_MUX_n146) ) ;
    INV_X1 Midori_rounds_constant_MUX_U37 ( .A (Midori_rounds_constant_MUX_n193), .ZN (Midori_rounds_constant_MUX_n147) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U36 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_round_Constant[0]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U35 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n144) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U34 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n143), .ZN (Midori_rounds_constant_MUX_n192) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U33 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n173), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n143) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U32 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n174) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U31 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n173) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U30 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n139), .ZN (Midori_rounds_constant_MUX_n203) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U29 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n176), .Z (Midori_rounds_constant_MUX_n139) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U28 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n152), .ZN (Midori_rounds_constant_MUX_n176) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U27 ( .A1 (round_Signal[3]), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n152) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U26 ( .A1 (Midori_rounds_constant_MUX_n138), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n166) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U25 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n137), .ZN (Midori_rounds_constant_MUX_n182) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U24 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_constant_MUX_n137) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U23 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n136), .ZN (Midori_rounds_constant_MUX_n216) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U22 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n142), .ZN (Midori_rounds_constant_MUX_n136) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U21 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n179), .ZN (Midori_rounds_constant_MUX_n163) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U20 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n179) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U19 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n161), .ZN (Midori_rounds_constant_MUX_n209) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U18 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n135), .ZN (Midori_rounds_constant_MUX_n161) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U17 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n177), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n135) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U16 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n134), .ZN (Midori_rounds_constant_MUX_n165) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U15 ( .A1 (round_Signal[3]), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n134) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U14 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n138), .ZN (Midori_rounds_constant_MUX_n177) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U13 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n133), .ZN (Midori_rounds_constant_MUX_n138) ) ;
    INV_X1 Midori_rounds_constant_MUX_U12 ( .A (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n133) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U11 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n132), .ZN (Midori_rounds_constant_MUX_n193) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U10 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n131), .Z (Midori_rounds_constant_MUX_n132) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U9 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n130), .ZN (Midori_rounds_constant_MUX_n184) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U8 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n131), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n130) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U7 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n153) ) ;
    INV_X1 Midori_rounds_constant_MUX_U6 ( .A (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n141) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U5 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n140) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U4 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n131) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U3 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n142) ) ;
    INV_X1 Midori_rounds_constant_MUX_U2 ( .A (Midori_rounds_constant_MUX_n129), .ZN (Midori_rounds_constant_MUX_n128) ) ;
    INV_X1 Midori_rounds_constant_MUX_U1 ( .A (round_Signal[0]), .ZN (Midori_rounds_constant_MUX_n129) ) ;
    INV_X1 Midori_rounds_MUXInst_U4 ( .A (round_Signal[0]), .ZN (Midori_rounds_MUXInst_n11) ) ;
    INV_X1 Midori_rounds_MUXInst_U3 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n8) ) ;
    INV_X1 Midori_rounds_MUXInst_U2 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n9) ) ;
    INV_X1 Midori_rounds_MUXInst_U1 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n10) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_0_U1 ( .s (round_Signal[0]), .b ({key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, Midori_rounds_SelectedKey_0_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_1_U1 ( .s (round_Signal[0]), .b ({key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, Midori_rounds_SelectedKey_1_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_2_U1 ( .s (round_Signal[0]), .b ({key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1845, new_AGEMA_signal_1844, Midori_rounds_SelectedKey_2_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_3_U1 ( .s (round_Signal[0]), .b ({key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, Midori_rounds_SelectedKey_3_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_4_U1 ( .s (round_Signal[0]), .b ({key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, Midori_rounds_SelectedKey_4_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_5_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, Midori_rounds_SelectedKey_5_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_6_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, Midori_rounds_SelectedKey_6_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_7_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, Midori_rounds_SelectedKey_7_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_8_U1 ( .s (round_Signal[0]), .b ({key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1851, new_AGEMA_signal_1850, Midori_rounds_SelectedKey_8_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_9_U1 ( .s (round_Signal[0]), .b ({key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, Midori_rounds_SelectedKey_9_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_10_U1 ( .s (round_Signal[0]), .b ({key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, Midori_rounds_SelectedKey_10_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_11_U1 ( .s (round_Signal[0]), .b ({key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1857, new_AGEMA_signal_1856, Midori_rounds_SelectedKey_11_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_12_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, Midori_rounds_SelectedKey_12_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_13_U1 ( .s (round_Signal[0]), .b ({key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, Midori_rounds_SelectedKey_13_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_14_U1 ( .s (round_Signal[0]), .b ({key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, Midori_rounds_SelectedKey_14_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_15_U1 ( .s (round_Signal[0]), .b ({key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1863, new_AGEMA_signal_1862, Midori_rounds_SelectedKey_15_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_16_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, Midori_rounds_SelectedKey_16_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_17_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, Midori_rounds_SelectedKey_17_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_18_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, Midori_rounds_SelectedKey_18_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_19_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, Midori_rounds_SelectedKey_19_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_20_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_2587, new_AGEMA_signal_2586, Midori_rounds_SelectedKey_20_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_21_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, Midori_rounds_SelectedKey_21_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_22_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, Midori_rounds_SelectedKey_22_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_23_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_2593, new_AGEMA_signal_2592, Midori_rounds_SelectedKey_23_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_24_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, Midori_rounds_SelectedKey_24_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_25_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, Midori_rounds_SelectedKey_25_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_26_U1 ( .s (round_Signal[0]), .b ({key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, Midori_rounds_SelectedKey_26_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_27_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, Midori_rounds_SelectedKey_27_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_28_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, Midori_rounds_SelectedKey_28_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_29_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, Midori_rounds_SelectedKey_29_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_30_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_2605, new_AGEMA_signal_2604, Midori_rounds_SelectedKey_30_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_31_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, Midori_rounds_SelectedKey_31_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_32_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, Midori_rounds_SelectedKey_32_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_33_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_2611, new_AGEMA_signal_2610, Midori_rounds_SelectedKey_33_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_34_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, Midori_rounds_SelectedKey_34_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_35_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, Midori_rounds_SelectedKey_35_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_36_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, Midori_rounds_SelectedKey_36_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_37_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, Midori_rounds_SelectedKey_37_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_38_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, Midori_rounds_SelectedKey_38_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_39_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_2623, new_AGEMA_signal_2622, Midori_rounds_SelectedKey_39_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_40_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, Midori_rounds_SelectedKey_40_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_41_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, Midori_rounds_SelectedKey_41_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_42_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, Midori_rounds_SelectedKey_42_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_43_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2631, new_AGEMA_signal_2630, Midori_rounds_SelectedKey_43_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_44_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, Midori_rounds_SelectedKey_44_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_45_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, Midori_rounds_SelectedKey_45_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_46_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2637, new_AGEMA_signal_2636, Midori_rounds_SelectedKey_46_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_47_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, Midori_rounds_SelectedKey_47_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_48_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, Midori_rounds_SelectedKey_48_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_49_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2643, new_AGEMA_signal_2642, Midori_rounds_SelectedKey_49_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_50_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, Midori_rounds_SelectedKey_50_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_51_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, Midori_rounds_SelectedKey_51_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_52_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2649, new_AGEMA_signal_2648, Midori_rounds_SelectedKey_52_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_53_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, Midori_rounds_SelectedKey_53_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_54_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, Midori_rounds_SelectedKey_54_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_55_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2655, new_AGEMA_signal_2654, Midori_rounds_SelectedKey_55_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_56_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, Midori_rounds_SelectedKey_56_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_57_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, Midori_rounds_SelectedKey_57_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_58_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2661, new_AGEMA_signal_2660, Midori_rounds_SelectedKey_58_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_59_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, Midori_rounds_SelectedKey_59_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_60_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, Midori_rounds_SelectedKey_60_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_61_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2667, new_AGEMA_signal_2666, Midori_rounds_SelectedKey_61_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_62_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, Midori_rounds_SelectedKey_62_}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_63_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, Midori_rounds_SelectedKey_63_}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U4 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U2 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U1 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U2 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U2 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U2 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U2 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U2 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U2 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U4 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U2 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U1 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U4 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U2 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U1 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U4 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U2 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U1 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U2 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U2 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U2 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U4 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U2 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U1 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U4 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U2 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U1 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U2 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}) ) ;

    /* cells in depth 1 */
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .a ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, Midori_rounds_sub_sBox_PRINCE_0_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .a ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, Midori_rounds_sub_sBox_PRINCE_0_n7}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, Midori_rounds_sub_sBox_PRINCE_0_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .a ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, Midori_rounds_sub_sBox_PRINCE_0_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, Midori_rounds_sub_sBox_PRINCE_0_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .a ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, Midori_rounds_sub_sBox_PRINCE_0_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .a ({new_AGEMA_signal_1881, new_AGEMA_signal_1880, Midori_rounds_sub_sBox_PRINCE_0_n9}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, Midori_rounds_sub_sBox_PRINCE_1_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .a ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .b ({new_AGEMA_signal_1893, new_AGEMA_signal_1892, Midori_rounds_sub_sBox_PRINCE_1_n7}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, Midori_rounds_sub_sBox_PRINCE_1_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .a ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, Midori_rounds_sub_sBox_PRINCE_1_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, Midori_rounds_sub_sBox_PRINCE_1_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U5 ( .a ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, Midori_rounds_sub_sBox_PRINCE_1_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U3 ( .a ({new_AGEMA_signal_1897, new_AGEMA_signal_1896, Midori_rounds_sub_sBox_PRINCE_1_n9}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .a ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, Midori_rounds_sub_sBox_PRINCE_2_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .a ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, Midori_rounds_sub_sBox_PRINCE_2_n7}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, Midori_rounds_sub_sBox_PRINCE_2_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .a ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, Midori_rounds_sub_sBox_PRINCE_2_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, Midori_rounds_sub_sBox_PRINCE_2_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U5 ( .a ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, Midori_rounds_sub_sBox_PRINCE_2_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U3 ( .a ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, Midori_rounds_sub_sBox_PRINCE_2_n9}), .b ({new_AGEMA_signal_1911, new_AGEMA_signal_1910, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .a ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_3_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .a ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .b ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_3_n7}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, Midori_rounds_sub_sBox_PRINCE_3_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .a ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, Midori_rounds_sub_sBox_PRINCE_3_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, Midori_rounds_sub_sBox_PRINCE_3_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U5 ( .a ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_3_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U3 ( .a ({new_AGEMA_signal_1929, new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_3_n9}), .b ({new_AGEMA_signal_1927, new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .a ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_4_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .a ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .b ({new_AGEMA_signal_1941, new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_4_n7}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, Midori_rounds_sub_sBox_PRINCE_4_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .a ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, Midori_rounds_sub_sBox_PRINCE_4_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_2433, new_AGEMA_signal_2432, Midori_rounds_sub_sBox_PRINCE_4_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U5 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_4_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U3 ( .a ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n9}), .b ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .a ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .a ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .b ({new_AGEMA_signal_1957, new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_5_n7}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, Midori_rounds_sub_sBox_PRINCE_5_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .a ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, Midori_rounds_sub_sBox_PRINCE_5_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_2445, new_AGEMA_signal_2444, Midori_rounds_sub_sBox_PRINCE_5_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U5 ( .a ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_5_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U3 ( .a ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_5_n9}), .b ({new_AGEMA_signal_1959, new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .a ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_6_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .a ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_6_n7}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, Midori_rounds_sub_sBox_PRINCE_6_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .a ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, Midori_rounds_sub_sBox_PRINCE_6_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_2457, new_AGEMA_signal_2456, Midori_rounds_sub_sBox_PRINCE_6_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U5 ( .a ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_6_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U3 ( .a ({new_AGEMA_signal_1977, new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_6_n9}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_7_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_7_n7}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, Midori_rounds_sub_sBox_PRINCE_7_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .a ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, Midori_rounds_sub_sBox_PRINCE_7_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_2469, new_AGEMA_signal_2468, Midori_rounds_sub_sBox_PRINCE_7_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .a ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_7_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .a ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_7_n9}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_8_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_8_n7}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, Midori_rounds_sub_sBox_PRINCE_8_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, Midori_rounds_sub_sBox_PRINCE_8_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, Midori_rounds_sub_sBox_PRINCE_8_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_8_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_8_n9}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .a ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, Midori_rounds_sub_sBox_PRINCE_9_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .a ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, Midori_rounds_sub_sBox_PRINCE_9_n7}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, Midori_rounds_sub_sBox_PRINCE_9_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, Midori_rounds_sub_sBox_PRINCE_9_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, Midori_rounds_sub_sBox_PRINCE_9_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .a ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, Midori_rounds_sub_sBox_PRINCE_9_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, Midori_rounds_sub_sBox_PRINCE_9_n9}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, Midori_rounds_sub_sBox_PRINCE_10_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .b ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, Midori_rounds_sub_sBox_PRINCE_10_n7}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, Midori_rounds_sub_sBox_PRINCE_10_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .a ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, Midori_rounds_sub_sBox_PRINCE_10_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, Midori_rounds_sub_sBox_PRINCE_10_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U5 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, Midori_rounds_sub_sBox_PRINCE_10_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U3 ( .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, Midori_rounds_sub_sBox_PRINCE_10_n9}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, Midori_rounds_sub_sBox_PRINCE_11_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, Midori_rounds_sub_sBox_PRINCE_11_n7}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, Midori_rounds_sub_sBox_PRINCE_11_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, Midori_rounds_sub_sBox_PRINCE_11_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, Midori_rounds_sub_sBox_PRINCE_11_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U5 ( .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_sub_sBox_PRINCE_11_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U3 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, Midori_rounds_sub_sBox_PRINCE_11_n9}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_sub_sBox_PRINCE_12_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .a ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .b ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_12_n7}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, Midori_rounds_sub_sBox_PRINCE_12_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, Midori_rounds_sub_sBox_PRINCE_12_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, Midori_rounds_sub_sBox_PRINCE_12_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U5 ( .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_12_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U3 ( .a ({new_AGEMA_signal_2073, new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_12_n9}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .a ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_13_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .b ({new_AGEMA_signal_2085, new_AGEMA_signal_2084, Midori_rounds_sub_sBox_PRINCE_13_n7}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, Midori_rounds_sub_sBox_PRINCE_13_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .a ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, Midori_rounds_sub_sBox_PRINCE_13_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, Midori_rounds_sub_sBox_PRINCE_13_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .a ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_13_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .a ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_13_n9}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .a ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, Midori_rounds_sub_sBox_PRINCE_14_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .a ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_14_n7}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, Midori_rounds_sub_sBox_PRINCE_14_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, Midori_rounds_sub_sBox_PRINCE_14_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, Midori_rounds_sub_sBox_PRINCE_14_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .a ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_14_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, Midori_rounds_sub_sBox_PRINCE_14_n9}), .b ({new_AGEMA_signal_2103, new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .a ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_15_n10}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_15_n7}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, Midori_rounds_sub_sBox_PRINCE_15_n15}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .a ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, Midori_rounds_sub_sBox_PRINCE_15_n4}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, Midori_rounds_sub_sBox_PRINCE_15_n6}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U5 ( .a ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, Midori_rounds_sub_sBox_PRINCE_15_n1}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U3 ( .a ({new_AGEMA_signal_2121, new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_15_n9}), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (Midori_rounds_roundReg_out[1]), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_2673), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n9), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_1880), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_1881), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (Midori_rounds_roundReg_out[0]), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (new_AGEMA_signal_1866), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_1867), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n7), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_1876), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_1877), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (Midori_rounds_roundReg_out[5]), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (new_AGEMA_signal_2682), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n9), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_1897), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (Midori_rounds_roundReg_out[4]), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_1883), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n7), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (new_AGEMA_signal_1893), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (Midori_rounds_roundReg_out[9]), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n9), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_1913), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (Midori_rounds_roundReg_out[8]), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_1899), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n7), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_1909), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (Midori_rounds_roundReg_out[13]), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_2703), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n9), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_1929), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (Midori_rounds_roundReg_out[12]), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (new_AGEMA_signal_1914), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (new_AGEMA_signal_1915), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n7), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_1924), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (new_AGEMA_signal_1925), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (Midori_rounds_roundReg_out[17]), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (new_AGEMA_signal_2712), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_2713), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n9), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (new_AGEMA_signal_1944), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_1945), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (Midori_rounds_roundReg_out[16]), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (new_AGEMA_signal_1930), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (new_AGEMA_signal_1931), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n7), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_1940), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_1941), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (Midori_rounds_roundReg_out[21]), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (new_AGEMA_signal_2722), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n9), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (new_AGEMA_signal_1960), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_1961), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (Midori_rounds_roundReg_out[20]), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (new_AGEMA_signal_1947), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n7), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_1956), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (new_AGEMA_signal_1957), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (Midori_rounds_roundReg_out[25]), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (new_AGEMA_signal_2732), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_2733), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n9), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (new_AGEMA_signal_1976), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_1977), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (Midori_rounds_roundReg_out[24]), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (new_AGEMA_signal_1962), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (new_AGEMA_signal_1963), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n7), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_1972), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_1973), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (Midori_rounds_roundReg_out[29]), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_2742), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_2743), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n9), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (new_AGEMA_signal_1992), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_1993), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (Midori_rounds_roundReg_out[28]), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_1978), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (new_AGEMA_signal_1979), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n7), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (Midori_rounds_roundReg_out[33]), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_2752), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_2753), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n9), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_2009), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (Midori_rounds_roundReg_out[32]), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (new_AGEMA_signal_1994), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (new_AGEMA_signal_1995), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n7), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (new_AGEMA_signal_2004), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_2005), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (Midori_rounds_roundReg_out[37]), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_2762), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_2763), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n9), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_2025), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (Midori_rounds_roundReg_out[36]), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_2010), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (new_AGEMA_signal_2011), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n7), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (new_AGEMA_signal_2020), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (new_AGEMA_signal_2021), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (Midori_rounds_roundReg_out[41]), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_2772), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n9), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (new_AGEMA_signal_2040), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_2041), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (Midori_rounds_roundReg_out[40]), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (new_AGEMA_signal_2027), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n7), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (new_AGEMA_signal_2036), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_2037), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (Midori_rounds_roundReg_out[45]), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_2783), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n9), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (new_AGEMA_signal_2056), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_2057), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (Midori_rounds_roundReg_out[44]), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_2042), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (new_AGEMA_signal_2043), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n7), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (new_AGEMA_signal_2052), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (new_AGEMA_signal_2053), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (Midori_rounds_roundReg_out[49]), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_2792), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n9), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (new_AGEMA_signal_2072), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_2073), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (Midori_rounds_roundReg_out[48]), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (new_AGEMA_signal_2058), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (new_AGEMA_signal_2059), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n7), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (new_AGEMA_signal_2068), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_2069), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (Midori_rounds_roundReg_out[53]), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_2803), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n9), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (new_AGEMA_signal_2088), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_2089), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (Midori_rounds_roundReg_out[52]), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_2074), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (new_AGEMA_signal_2075), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n7), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (new_AGEMA_signal_2084), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (new_AGEMA_signal_2085), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (Midori_rounds_roundReg_out[57]), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_2812), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n9), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (new_AGEMA_signal_2104), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_2105), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (Midori_rounds_roundReg_out[56]), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (new_AGEMA_signal_2090), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (new_AGEMA_signal_2091), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n7), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (new_AGEMA_signal_2100), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_2101), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (Midori_rounds_roundReg_out[61]), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_2823), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n9), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (new_AGEMA_signal_2120), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_2121), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (Midori_rounds_roundReg_out[60]), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_2106), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (new_AGEMA_signal_2107), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n7), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (new_AGEMA_signal_2116), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_2117), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (wk[9]), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_1460), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (wk[7]), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (new_AGEMA_signal_1472), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_1473), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (wk[63]), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_1484), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (wk[61]), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_1496), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (wk[5]), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (new_AGEMA_signal_1508), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (wk[59]), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (new_AGEMA_signal_1514), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (wk[57]), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_1526), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (new_AGEMA_signal_1527), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (wk[55]), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_1538), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_1539), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (wk[53]), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_1550), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (wk[51]), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (new_AGEMA_signal_1562), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_1563), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (wk[49]), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_1580), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (new_AGEMA_signal_1581), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (wk[47]), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_1592), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_1593), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (wk[45]), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (new_AGEMA_signal_1604), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_1605), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (wk[43]), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (new_AGEMA_signal_1616), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_1617), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (wk[41]), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_1628), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (new_AGEMA_signal_1629), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (wk[3]), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_1640), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_1641), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (wk[39]), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_1646), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_1647), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (wk[37]), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_1659), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (wk[35]), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_1670), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_1671), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (wk[33]), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_1682), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_1683), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (wk[31]), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_1694), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_1695), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (wk[29]), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (wk[27]), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_1725), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (wk[25]), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_1736), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_1737), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (wk[23]), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_1748), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_1749), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (wk[21]), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_1760), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_1761), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (wk[1]), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (wk[19]), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_1778), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_1779), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (wk[17]), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_1790), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_1791), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (wk[15]), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_1803), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (wk[13]), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_1814), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_1815), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (wk[11]), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_1826), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_1827), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (Midori_rounds_SelectedKey_9_), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_1853), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (Midori_rounds_SelectedKey_7_), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_2574), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_2575), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (Midori_rounds_SelectedKey_63_), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_2670), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_2671), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (Midori_rounds_SelectedKey_61_), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_2667), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (Midori_rounds_SelectedKey_5_), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_2571), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (Midori_rounds_SelectedKey_59_), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_2662), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_2663), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (Midori_rounds_SelectedKey_57_), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_2659), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (Midori_rounds_SelectedKey_55_), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_2655), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (Midori_rounds_SelectedKey_53_), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_2650), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_2651), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (Midori_rounds_SelectedKey_51_), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (Midori_rounds_SelectedKey_49_), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_2643), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (Midori_rounds_SelectedKey_47_), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (Midori_rounds_SelectedKey_45_), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (Midori_rounds_SelectedKey_43_), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_2631), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (Midori_rounds_SelectedKey_41_), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_2626), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_2627), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (Midori_rounds_SelectedKey_3_), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_1847), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (Midori_rounds_SelectedKey_39_), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (Midori_rounds_SelectedKey_37_), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_2619), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (Midori_rounds_SelectedKey_35_), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_2614), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_2615), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (Midori_rounds_SelectedKey_33_), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_2610), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (Midori_rounds_SelectedKey_31_), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_2607), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (Midori_rounds_SelectedKey_29_), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_2602), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (Midori_rounds_SelectedKey_27_), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (Midori_rounds_SelectedKey_25_), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_2596), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (Midori_rounds_SelectedKey_23_), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_2593), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (Midori_rounds_SelectedKey_21_), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_6296) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_2589), .Q (new_AGEMA_signal_6299) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (Midori_rounds_SelectedKey_1_), .Q (new_AGEMA_signal_6302) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_1842), .Q (new_AGEMA_signal_6305) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_1843), .Q (new_AGEMA_signal_6308) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (Midori_rounds_SelectedKey_19_), .Q (new_AGEMA_signal_6311) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_2584), .Q (new_AGEMA_signal_6314) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_6317) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (Midori_rounds_SelectedKey_17_), .Q (new_AGEMA_signal_6320) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_2580), .Q (new_AGEMA_signal_6323) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_2581), .Q (new_AGEMA_signal_6326) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (Midori_rounds_SelectedKey_15_), .Q (new_AGEMA_signal_6329) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_1862), .Q (new_AGEMA_signal_6332) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_1863), .Q (new_AGEMA_signal_6335) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (Midori_rounds_SelectedKey_13_), .Q (new_AGEMA_signal_6338) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_6341) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_1859), .Q (new_AGEMA_signal_6344) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (Midori_rounds_SelectedKey_11_), .Q (new_AGEMA_signal_6347) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_6350) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_1857), .Q (new_AGEMA_signal_6353) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_6356) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (Midori_add_Result_Start[1]), .Q (new_AGEMA_signal_6359) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_2332), .Q (new_AGEMA_signal_6362) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_2333), .Q (new_AGEMA_signal_6365) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (Midori_add_Result_Start[3]), .Q (new_AGEMA_signal_6368) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_2244), .Q (new_AGEMA_signal_6371) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_2245), .Q (new_AGEMA_signal_6374) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (Midori_add_Result_Start[5]), .Q (new_AGEMA_signal_6377) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_2156), .Q (new_AGEMA_signal_6380) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_2157), .Q (new_AGEMA_signal_6383) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (Midori_add_Result_Start[7]), .Q (new_AGEMA_signal_6386) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_2132), .Q (new_AGEMA_signal_6389) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_2133), .Q (new_AGEMA_signal_6392) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (Midori_add_Result_Start[9]), .Q (new_AGEMA_signal_6395) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_2124), .Q (new_AGEMA_signal_6398) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_2125), .Q (new_AGEMA_signal_6401) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (Midori_add_Result_Start[11]), .Q (new_AGEMA_signal_6404) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_2368), .Q (new_AGEMA_signal_6407) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_6410) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (Midori_add_Result_Start[13]), .Q (new_AGEMA_signal_6413) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_2360), .Q (new_AGEMA_signal_6416) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_2361), .Q (new_AGEMA_signal_6419) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (Midori_add_Result_Start[15]), .Q (new_AGEMA_signal_6422) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_2352), .Q (new_AGEMA_signal_6425) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_2353), .Q (new_AGEMA_signal_6428) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (Midori_add_Result_Start[17]), .Q (new_AGEMA_signal_6431) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_2344), .Q (new_AGEMA_signal_6434) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_2345), .Q (new_AGEMA_signal_6437) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (Midori_add_Result_Start[19]), .Q (new_AGEMA_signal_6440) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_2336), .Q (new_AGEMA_signal_6443) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_2337), .Q (new_AGEMA_signal_6446) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (Midori_add_Result_Start[21]), .Q (new_AGEMA_signal_6449) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_2324), .Q (new_AGEMA_signal_6452) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_2325), .Q (new_AGEMA_signal_6455) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (Midori_add_Result_Start[23]), .Q (new_AGEMA_signal_6458) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_2316), .Q (new_AGEMA_signal_6461) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_2317), .Q (new_AGEMA_signal_6464) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (Midori_add_Result_Start[25]), .Q (new_AGEMA_signal_6467) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_2308), .Q (new_AGEMA_signal_6470) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_2309), .Q (new_AGEMA_signal_6473) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (Midori_add_Result_Start[27]), .Q (new_AGEMA_signal_6476) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_2300), .Q (new_AGEMA_signal_6479) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_2301), .Q (new_AGEMA_signal_6482) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (Midori_add_Result_Start[29]), .Q (new_AGEMA_signal_6485) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_2292), .Q (new_AGEMA_signal_6488) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_2293), .Q (new_AGEMA_signal_6491) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (Midori_add_Result_Start[31]), .Q (new_AGEMA_signal_6494) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_2280), .Q (new_AGEMA_signal_6497) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_2281), .Q (new_AGEMA_signal_6500) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (Midori_add_Result_Start[33]), .Q (new_AGEMA_signal_6503) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_2272), .Q (new_AGEMA_signal_6506) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_2273), .Q (new_AGEMA_signal_6509) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (Midori_add_Result_Start[35]), .Q (new_AGEMA_signal_6512) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_2264), .Q (new_AGEMA_signal_6515) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_2265), .Q (new_AGEMA_signal_6518) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (Midori_add_Result_Start[37]), .Q (new_AGEMA_signal_6521) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_2256), .Q (new_AGEMA_signal_6524) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_2257), .Q (new_AGEMA_signal_6527) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (Midori_add_Result_Start[39]), .Q (new_AGEMA_signal_6530) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_2248), .Q (new_AGEMA_signal_6533) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_2249), .Q (new_AGEMA_signal_6536) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (Midori_add_Result_Start[41]), .Q (new_AGEMA_signal_6539) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_2236), .Q (new_AGEMA_signal_6542) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_2237), .Q (new_AGEMA_signal_6545) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (Midori_add_Result_Start[43]), .Q (new_AGEMA_signal_6548) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_2228), .Q (new_AGEMA_signal_6551) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_2229), .Q (new_AGEMA_signal_6554) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (Midori_add_Result_Start[45]), .Q (new_AGEMA_signal_6557) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_2220), .Q (new_AGEMA_signal_6560) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_2221), .Q (new_AGEMA_signal_6563) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (Midori_add_Result_Start[47]), .Q (new_AGEMA_signal_6566) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_2212), .Q (new_AGEMA_signal_6569) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_2213), .Q (new_AGEMA_signal_6572) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (Midori_add_Result_Start[49]), .Q (new_AGEMA_signal_6575) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_2204), .Q (new_AGEMA_signal_6578) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_2205), .Q (new_AGEMA_signal_6581) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (Midori_add_Result_Start[51]), .Q (new_AGEMA_signal_6584) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_2192), .Q (new_AGEMA_signal_6587) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_2193), .Q (new_AGEMA_signal_6590) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (Midori_add_Result_Start[53]), .Q (new_AGEMA_signal_6593) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_2184), .Q (new_AGEMA_signal_6596) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_2185), .Q (new_AGEMA_signal_6599) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (Midori_add_Result_Start[55]), .Q (new_AGEMA_signal_6602) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_2176), .Q (new_AGEMA_signal_6605) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_2177), .Q (new_AGEMA_signal_6608) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (Midori_add_Result_Start[57]), .Q (new_AGEMA_signal_6611) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_2168), .Q (new_AGEMA_signal_6614) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_2169), .Q (new_AGEMA_signal_6617) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (Midori_add_Result_Start[59]), .Q (new_AGEMA_signal_6620) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_2160), .Q (new_AGEMA_signal_6623) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_2161), .Q (new_AGEMA_signal_6626) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (Midori_add_Result_Start[61]), .Q (new_AGEMA_signal_6629) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_2148), .Q (new_AGEMA_signal_6632) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_2149), .Q (new_AGEMA_signal_6635) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (Midori_add_Result_Start[63]), .Q (new_AGEMA_signal_6638) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_2140), .Q (new_AGEMA_signal_6641) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_2141), .Q (new_AGEMA_signal_6644) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (enc_dec), .Q (new_AGEMA_signal_6791) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (wk[8]), .Q (new_AGEMA_signal_6794) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_1466), .Q (new_AGEMA_signal_6798) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_6802) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (wk[6]), .Q (new_AGEMA_signal_6806) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (new_AGEMA_signal_1478), .Q (new_AGEMA_signal_6810) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_6814) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (wk[62]), .Q (new_AGEMA_signal_6818) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (new_AGEMA_signal_1490), .Q (new_AGEMA_signal_6822) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_6826) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (wk[60]), .Q (new_AGEMA_signal_6830) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_1502), .Q (new_AGEMA_signal_6834) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_6838) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (wk[58]), .Q (new_AGEMA_signal_6842) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (new_AGEMA_signal_1520), .Q (new_AGEMA_signal_6846) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_6850) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (wk[56]), .Q (new_AGEMA_signal_6854) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_1532), .Q (new_AGEMA_signal_6858) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_1533), .Q (new_AGEMA_signal_6862) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (wk[54]), .Q (new_AGEMA_signal_6866) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_1544), .Q (new_AGEMA_signal_6870) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_1545), .Q (new_AGEMA_signal_6874) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (wk[52]), .Q (new_AGEMA_signal_6878) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_1556), .Q (new_AGEMA_signal_6882) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_6886) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (wk[50]), .Q (new_AGEMA_signal_6890) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_1568), .Q (new_AGEMA_signal_6894) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_6898) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (wk[4]), .Q (new_AGEMA_signal_6902) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_1574), .Q (new_AGEMA_signal_6906) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_6910) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (wk[48]), .Q (new_AGEMA_signal_6914) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_1586), .Q (new_AGEMA_signal_6918) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_1587), .Q (new_AGEMA_signal_6922) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (wk[46]), .Q (new_AGEMA_signal_6926) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_1598), .Q (new_AGEMA_signal_6930) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_1599), .Q (new_AGEMA_signal_6934) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (wk[44]), .Q (new_AGEMA_signal_6938) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_1610), .Q (new_AGEMA_signal_6942) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_1611), .Q (new_AGEMA_signal_6946) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (wk[42]), .Q (new_AGEMA_signal_6950) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_1622), .Q (new_AGEMA_signal_6954) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_1623), .Q (new_AGEMA_signal_6958) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (wk[40]), .Q (new_AGEMA_signal_6962) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_1634), .Q (new_AGEMA_signal_6966) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_1635), .Q (new_AGEMA_signal_6970) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (wk[38]), .Q (new_AGEMA_signal_6974) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_1652), .Q (new_AGEMA_signal_6978) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_1653), .Q (new_AGEMA_signal_6982) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (wk[36]), .Q (new_AGEMA_signal_6986) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_1664), .Q (new_AGEMA_signal_6990) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_1665), .Q (new_AGEMA_signal_6994) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (wk[34]), .Q (new_AGEMA_signal_6998) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_7002) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_1677), .Q (new_AGEMA_signal_7006) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (wk[32]), .Q (new_AGEMA_signal_7010) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_1688), .Q (new_AGEMA_signal_7014) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_1689), .Q (new_AGEMA_signal_7018) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (wk[30]), .Q (new_AGEMA_signal_7022) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_1700), .Q (new_AGEMA_signal_7026) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_1701), .Q (new_AGEMA_signal_7030) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (wk[2]), .Q (new_AGEMA_signal_7034) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_7038) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_1707), .Q (new_AGEMA_signal_7042) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (wk[28]), .Q (new_AGEMA_signal_7046) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_1718), .Q (new_AGEMA_signal_7050) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_1719), .Q (new_AGEMA_signal_7054) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (wk[26]), .Q (new_AGEMA_signal_7058) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_1730), .Q (new_AGEMA_signal_7062) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_1731), .Q (new_AGEMA_signal_7066) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (wk[24]), .Q (new_AGEMA_signal_7070) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_1742), .Q (new_AGEMA_signal_7074) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_1743), .Q (new_AGEMA_signal_7078) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (wk[22]), .Q (new_AGEMA_signal_7082) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (new_AGEMA_signal_1754), .Q (new_AGEMA_signal_7086) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_1755), .Q (new_AGEMA_signal_7090) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (wk[20]), .Q (new_AGEMA_signal_7094) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (new_AGEMA_signal_1766), .Q (new_AGEMA_signal_7098) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_1767), .Q (new_AGEMA_signal_7102) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (wk[18]), .Q (new_AGEMA_signal_7106) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (new_AGEMA_signal_1784), .Q (new_AGEMA_signal_7110) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_1785), .Q (new_AGEMA_signal_7114) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (wk[16]), .Q (new_AGEMA_signal_7118) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (new_AGEMA_signal_1796), .Q (new_AGEMA_signal_7122) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_1797), .Q (new_AGEMA_signal_7126) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (wk[14]), .Q (new_AGEMA_signal_7130) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (new_AGEMA_signal_1808), .Q (new_AGEMA_signal_7134) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_1809), .Q (new_AGEMA_signal_7138) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (wk[12]), .Q (new_AGEMA_signal_7142) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_7146) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_1821), .Q (new_AGEMA_signal_7150) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (wk[10]), .Q (new_AGEMA_signal_7154) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_7158) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_1833), .Q (new_AGEMA_signal_7162) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (wk[0]), .Q (new_AGEMA_signal_7166) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_7170) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_1839), .Q (new_AGEMA_signal_7174) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (Midori_rounds_n16), .Q (new_AGEMA_signal_7178) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_3426), .Q (new_AGEMA_signal_7182) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_3427), .Q (new_AGEMA_signal_7186) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (Midori_rounds_SelectedKey_6_), .Q (new_AGEMA_signal_7190) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (new_AGEMA_signal_2572), .Q (new_AGEMA_signal_7194) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_2573), .Q (new_AGEMA_signal_7198) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (Midori_rounds_SelectedKey_62_), .Q (new_AGEMA_signal_7202) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_2668), .Q (new_AGEMA_signal_7206) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_7210) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (Midori_rounds_n15), .Q (new_AGEMA_signal_7214) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_7218) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_3537), .Q (new_AGEMA_signal_7222) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (Midori_rounds_SelectedKey_58_), .Q (new_AGEMA_signal_7226) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_7230) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_2661), .Q (new_AGEMA_signal_7234) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (Midori_rounds_n14), .Q (new_AGEMA_signal_7238) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_3538), .Q (new_AGEMA_signal_7242) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_3539), .Q (new_AGEMA_signal_7246) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (Midori_rounds_SelectedKey_54_), .Q (new_AGEMA_signal_7250) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_2652), .Q (new_AGEMA_signal_7254) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_2653), .Q (new_AGEMA_signal_7258) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (Midori_rounds_n13), .Q (new_AGEMA_signal_7262) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_7266) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_7270) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (Midori_rounds_SelectedKey_50_), .Q (new_AGEMA_signal_7274) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_2644), .Q (new_AGEMA_signal_7278) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_7282) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (Midori_rounds_n12), .Q (new_AGEMA_signal_7286) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_3542), .Q (new_AGEMA_signal_7290) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_3543), .Q (new_AGEMA_signal_7294) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (Midori_rounds_n11), .Q (new_AGEMA_signal_7298) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_3780), .Q (new_AGEMA_signal_7302) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_3781), .Q (new_AGEMA_signal_7306) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (Midori_rounds_SelectedKey_46_), .Q (new_AGEMA_signal_7310) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_7314) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_2637), .Q (new_AGEMA_signal_7318) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (Midori_rounds_n10), .Q (new_AGEMA_signal_7322) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_7326) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_3465), .Q (new_AGEMA_signal_7330) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (Midori_rounds_SelectedKey_42_), .Q (new_AGEMA_signal_7334) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_2628), .Q (new_AGEMA_signal_7338) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_2629), .Q (new_AGEMA_signal_7342) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (Midori_rounds_n9), .Q (new_AGEMA_signal_7346) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_7350) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_7354) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (Midori_rounds_SelectedKey_38_), .Q (new_AGEMA_signal_7358) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_2620), .Q (new_AGEMA_signal_7362) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_7366) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (Midori_rounds_n8), .Q (new_AGEMA_signal_7370) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_7374) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_7378) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (Midori_rounds_SelectedKey_34_), .Q (new_AGEMA_signal_7382) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_7386) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_2613), .Q (new_AGEMA_signal_7390) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (Midori_rounds_n7), .Q (new_AGEMA_signal_7394) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_3546), .Q (new_AGEMA_signal_7398) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_3547), .Q (new_AGEMA_signal_7402) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (Midori_rounds_SelectedKey_30_), .Q (new_AGEMA_signal_7406) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_7410) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_2605), .Q (new_AGEMA_signal_7414) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (Midori_rounds_SelectedKey_2_), .Q (new_AGEMA_signal_7418) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_7422) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_1845), .Q (new_AGEMA_signal_7426) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (Midori_rounds_n6), .Q (new_AGEMA_signal_7430) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_7434) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_7438) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (Midori_rounds_SelectedKey_26_), .Q (new_AGEMA_signal_7442) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_1864), .Q (new_AGEMA_signal_7446) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_1865), .Q (new_AGEMA_signal_7450) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (Midori_rounds_n5), .Q (new_AGEMA_signal_7454) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_7458) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_3549), .Q (new_AGEMA_signal_7462) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (Midori_rounds_SelectedKey_22_), .Q (new_AGEMA_signal_7466) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_2590), .Q (new_AGEMA_signal_7470) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_7474) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (Midori_rounds_n4), .Q (new_AGEMA_signal_7478) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_7482) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_7486) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (Midori_rounds_SelectedKey_18_), .Q (new_AGEMA_signal_7490) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_7494) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_2583), .Q (new_AGEMA_signal_7498) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (Midori_rounds_n3), .Q (new_AGEMA_signal_7502) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_3550), .Q (new_AGEMA_signal_7506) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_3551), .Q (new_AGEMA_signal_7510) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (Midori_rounds_SelectedKey_14_), .Q (new_AGEMA_signal_7514) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (new_AGEMA_signal_1860), .Q (new_AGEMA_signal_7518) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_1861), .Q (new_AGEMA_signal_7522) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (Midori_rounds_n2), .Q (new_AGEMA_signal_7526) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_7530) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_7534) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (Midori_rounds_SelectedKey_10_), .Q (new_AGEMA_signal_7538) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_7542) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_1855), .Q (new_AGEMA_signal_7546) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (Midori_rounds_n1), .Q (new_AGEMA_signal_7550) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (new_AGEMA_signal_3554), .Q (new_AGEMA_signal_7554) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_3555), .Q (new_AGEMA_signal_7558) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (Midori_add_Result_Start[0]), .Q (new_AGEMA_signal_7563) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_2376), .Q (new_AGEMA_signal_7567) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_2377), .Q (new_AGEMA_signal_7571) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (Midori_add_Result_Start[2]), .Q (new_AGEMA_signal_7575) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_2288), .Q (new_AGEMA_signal_7579) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_2289), .Q (new_AGEMA_signal_7583) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (Midori_add_Result_Start[4]), .Q (new_AGEMA_signal_7587) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_2200), .Q (new_AGEMA_signal_7591) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_2201), .Q (new_AGEMA_signal_7595) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (Midori_add_Result_Start[6]), .Q (new_AGEMA_signal_7599) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_2136), .Q (new_AGEMA_signal_7603) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_2137), .Q (new_AGEMA_signal_7607) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (Midori_add_Result_Start[8]), .Q (new_AGEMA_signal_7611) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_2128), .Q (new_AGEMA_signal_7615) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_2129), .Q (new_AGEMA_signal_7619) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (Midori_add_Result_Start[10]), .Q (new_AGEMA_signal_7623) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_2372), .Q (new_AGEMA_signal_7627) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_2373), .Q (new_AGEMA_signal_7631) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (Midori_add_Result_Start[12]), .Q (new_AGEMA_signal_7635) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_2364), .Q (new_AGEMA_signal_7639) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_2365), .Q (new_AGEMA_signal_7643) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (Midori_add_Result_Start[14]), .Q (new_AGEMA_signal_7647) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_2356), .Q (new_AGEMA_signal_7651) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_2357), .Q (new_AGEMA_signal_7655) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (Midori_add_Result_Start[16]), .Q (new_AGEMA_signal_7659) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_2348), .Q (new_AGEMA_signal_7663) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_2349), .Q (new_AGEMA_signal_7667) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (Midori_add_Result_Start[18]), .Q (new_AGEMA_signal_7671) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_2340), .Q (new_AGEMA_signal_7675) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_2341), .Q (new_AGEMA_signal_7679) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (Midori_add_Result_Start[20]), .Q (new_AGEMA_signal_7683) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_2328), .Q (new_AGEMA_signal_7687) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_2329), .Q (new_AGEMA_signal_7691) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (Midori_add_Result_Start[22]), .Q (new_AGEMA_signal_7695) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_2320), .Q (new_AGEMA_signal_7699) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_2321), .Q (new_AGEMA_signal_7703) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (clk), .D (Midori_add_Result_Start[24]), .Q (new_AGEMA_signal_7707) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_2312), .Q (new_AGEMA_signal_7711) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_2313), .Q (new_AGEMA_signal_7715) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (clk), .D (Midori_add_Result_Start[26]), .Q (new_AGEMA_signal_7719) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_2304), .Q (new_AGEMA_signal_7723) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_2305), .Q (new_AGEMA_signal_7727) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (clk), .D (Midori_add_Result_Start[28]), .Q (new_AGEMA_signal_7731) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_2296), .Q (new_AGEMA_signal_7735) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_2297), .Q (new_AGEMA_signal_7739) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (clk), .D (Midori_add_Result_Start[30]), .Q (new_AGEMA_signal_7743) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_2284), .Q (new_AGEMA_signal_7747) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_2285), .Q (new_AGEMA_signal_7751) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (clk), .D (Midori_add_Result_Start[32]), .Q (new_AGEMA_signal_7755) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_2276), .Q (new_AGEMA_signal_7759) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_2277), .Q (new_AGEMA_signal_7763) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (clk), .D (Midori_add_Result_Start[34]), .Q (new_AGEMA_signal_7767) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_2268), .Q (new_AGEMA_signal_7771) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_2269), .Q (new_AGEMA_signal_7775) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (clk), .D (Midori_add_Result_Start[36]), .Q (new_AGEMA_signal_7779) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_2260), .Q (new_AGEMA_signal_7783) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_2261), .Q (new_AGEMA_signal_7787) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (clk), .D (Midori_add_Result_Start[38]), .Q (new_AGEMA_signal_7791) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_2252), .Q (new_AGEMA_signal_7795) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_2253), .Q (new_AGEMA_signal_7799) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (clk), .D (Midori_add_Result_Start[40]), .Q (new_AGEMA_signal_7803) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_2240), .Q (new_AGEMA_signal_7807) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_2241), .Q (new_AGEMA_signal_7811) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (clk), .D (Midori_add_Result_Start[42]), .Q (new_AGEMA_signal_7815) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_2232), .Q (new_AGEMA_signal_7819) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_2233), .Q (new_AGEMA_signal_7823) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (clk), .D (Midori_add_Result_Start[44]), .Q (new_AGEMA_signal_7827) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_2224), .Q (new_AGEMA_signal_7831) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_2225), .Q (new_AGEMA_signal_7835) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (clk), .D (Midori_add_Result_Start[46]), .Q (new_AGEMA_signal_7839) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_2216), .Q (new_AGEMA_signal_7843) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_2217), .Q (new_AGEMA_signal_7847) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (clk), .D (Midori_add_Result_Start[48]), .Q (new_AGEMA_signal_7851) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_2208), .Q (new_AGEMA_signal_7855) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_2209), .Q (new_AGEMA_signal_7859) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (clk), .D (Midori_add_Result_Start[50]), .Q (new_AGEMA_signal_7863) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_2196), .Q (new_AGEMA_signal_7867) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_2197), .Q (new_AGEMA_signal_7871) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (Midori_add_Result_Start[52]), .Q (new_AGEMA_signal_7875) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_2188), .Q (new_AGEMA_signal_7879) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_2189), .Q (new_AGEMA_signal_7883) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (clk), .D (Midori_add_Result_Start[54]), .Q (new_AGEMA_signal_7887) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_2180), .Q (new_AGEMA_signal_7891) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_2181), .Q (new_AGEMA_signal_7895) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (Midori_add_Result_Start[56]), .Q (new_AGEMA_signal_7899) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_2172), .Q (new_AGEMA_signal_7903) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_2173), .Q (new_AGEMA_signal_7907) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (clk), .D (Midori_add_Result_Start[58]), .Q (new_AGEMA_signal_7911) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_2164), .Q (new_AGEMA_signal_7915) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_2165), .Q (new_AGEMA_signal_7919) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (clk), .D (Midori_add_Result_Start[60]), .Q (new_AGEMA_signal_7923) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_2152), .Q (new_AGEMA_signal_7927) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_2153), .Q (new_AGEMA_signal_7931) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (clk), .D (Midori_add_Result_Start[62]), .Q (new_AGEMA_signal_7935) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_2144), .Q (new_AGEMA_signal_7939) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_2145), .Q (new_AGEMA_signal_7943) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C (clk), .D (controller_roundCounter_N7), .Q (new_AGEMA_signal_8092) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C (clk), .D (controller_roundCounter_N8), .Q (new_AGEMA_signal_8096) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C (clk), .D (controller_roundCounter_n2), .Q (new_AGEMA_signal_8100) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C (clk), .D (controller_roundCounter_N10), .Q (new_AGEMA_signal_8104) ) ;

    /* cells in depth 2 */
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .a ({new_AGEMA_signal_2389, new_AGEMA_signal_2388, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_5590, new_AGEMA_signal_5589, new_AGEMA_signal_5588}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_rounds_sub_sBox_PRINCE_0_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .a ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, Midori_rounds_sub_sBox_PRINCE_0_n10}), .b ({new_AGEMA_signal_5593, new_AGEMA_signal_5592, new_AGEMA_signal_5591}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, Midori_rounds_sub_sBox_PRINCE_0_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .a ({new_AGEMA_signal_5596, new_AGEMA_signal_5595, new_AGEMA_signal_5594}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, Midori_rounds_sub_sBox_PRINCE_0_n4}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, Midori_rounds_sub_sBox_PRINCE_0_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .a ({new_AGEMA_signal_5599, new_AGEMA_signal_5598, new_AGEMA_signal_5597}), .b ({new_AGEMA_signal_1875, new_AGEMA_signal_1874, Midori_rounds_sub_sBox_PRINCE_0_n1}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_sub_sBox_PRINCE_0_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .a ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_5602, new_AGEMA_signal_5601, new_AGEMA_signal_5600}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, Midori_rounds_sub_sBox_PRINCE_1_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .a ({new_AGEMA_signal_1887, new_AGEMA_signal_1886, Midori_rounds_sub_sBox_PRINCE_1_n10}), .b ({new_AGEMA_signal_5605, new_AGEMA_signal_5604, new_AGEMA_signal_5603}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, Midori_rounds_sub_sBox_PRINCE_1_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .a ({new_AGEMA_signal_5608, new_AGEMA_signal_5607, new_AGEMA_signal_5606}), .b ({new_AGEMA_signal_2395, new_AGEMA_signal_2394, Midori_rounds_sub_sBox_PRINCE_1_n4}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, Midori_rounds_sub_sBox_PRINCE_1_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .a ({new_AGEMA_signal_5611, new_AGEMA_signal_5610, new_AGEMA_signal_5609}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, Midori_rounds_sub_sBox_PRINCE_1_n1}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_1_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .a ({new_AGEMA_signal_2413, new_AGEMA_signal_2412, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_5614, new_AGEMA_signal_5613, new_AGEMA_signal_5612}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, Midori_rounds_sub_sBox_PRINCE_2_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .a ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, Midori_rounds_sub_sBox_PRINCE_2_n10}), .b ({new_AGEMA_signal_5617, new_AGEMA_signal_5616, new_AGEMA_signal_5615}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, Midori_rounds_sub_sBox_PRINCE_2_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .a ({new_AGEMA_signal_5620, new_AGEMA_signal_5619, new_AGEMA_signal_5618}), .b ({new_AGEMA_signal_2407, new_AGEMA_signal_2406, Midori_rounds_sub_sBox_PRINCE_2_n4}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_rounds_sub_sBox_PRINCE_2_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .a ({new_AGEMA_signal_5623, new_AGEMA_signal_5622, new_AGEMA_signal_5621}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, Midori_rounds_sub_sBox_PRINCE_2_n1}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_sub_sBox_PRINCE_2_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .a ({new_AGEMA_signal_2425, new_AGEMA_signal_2424, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_5626, new_AGEMA_signal_5625, new_AGEMA_signal_5624}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_rounds_sub_sBox_PRINCE_3_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .a ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_3_n10}), .b ({new_AGEMA_signal_5629, new_AGEMA_signal_5628, new_AGEMA_signal_5627}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, Midori_rounds_sub_sBox_PRINCE_3_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .a ({new_AGEMA_signal_5632, new_AGEMA_signal_5631, new_AGEMA_signal_5630}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, Midori_rounds_sub_sBox_PRINCE_3_n4}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, Midori_rounds_sub_sBox_PRINCE_3_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .a ({new_AGEMA_signal_5635, new_AGEMA_signal_5634, new_AGEMA_signal_5633}), .b ({new_AGEMA_signal_1923, new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_3_n1}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_3_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .a ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_5638, new_AGEMA_signal_5637, new_AGEMA_signal_5636}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, Midori_rounds_sub_sBox_PRINCE_4_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .a ({new_AGEMA_signal_1935, new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_4_n10}), .b ({new_AGEMA_signal_5641, new_AGEMA_signal_5640, new_AGEMA_signal_5639}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, Midori_rounds_sub_sBox_PRINCE_4_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .a ({new_AGEMA_signal_5644, new_AGEMA_signal_5643, new_AGEMA_signal_5642}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, Midori_rounds_sub_sBox_PRINCE_4_n4}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, Midori_rounds_sub_sBox_PRINCE_4_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .a ({new_AGEMA_signal_5647, new_AGEMA_signal_5646, new_AGEMA_signal_5645}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_4_n1}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_sub_sBox_PRINCE_4_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .a ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_5650, new_AGEMA_signal_5649, new_AGEMA_signal_5648}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, Midori_rounds_sub_sBox_PRINCE_5_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .a ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n10}), .b ({new_AGEMA_signal_5653, new_AGEMA_signal_5652, new_AGEMA_signal_5651}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, Midori_rounds_sub_sBox_PRINCE_5_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .a ({new_AGEMA_signal_5656, new_AGEMA_signal_5655, new_AGEMA_signal_5654}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, Midori_rounds_sub_sBox_PRINCE_5_n4}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_rounds_sub_sBox_PRINCE_5_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .a ({new_AGEMA_signal_5659, new_AGEMA_signal_5658, new_AGEMA_signal_5657}), .b ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_5_n1}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_5_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .a ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_5662, new_AGEMA_signal_5661, new_AGEMA_signal_5660}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_rounds_sub_sBox_PRINCE_6_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .a ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_6_n10}), .b ({new_AGEMA_signal_5665, new_AGEMA_signal_5664, new_AGEMA_signal_5663}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, Midori_rounds_sub_sBox_PRINCE_6_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .a ({new_AGEMA_signal_5668, new_AGEMA_signal_5667, new_AGEMA_signal_5666}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, Midori_rounds_sub_sBox_PRINCE_6_n4}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, Midori_rounds_sub_sBox_PRINCE_6_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .a ({new_AGEMA_signal_5671, new_AGEMA_signal_5670, new_AGEMA_signal_5669}), .b ({new_AGEMA_signal_1971, new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_6_n1}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_rounds_sub_sBox_PRINCE_6_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .a ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_5674, new_AGEMA_signal_5673, new_AGEMA_signal_5672}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, Midori_rounds_sub_sBox_PRINCE_7_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .a ({new_AGEMA_signal_1983, new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_7_n10}), .b ({new_AGEMA_signal_5677, new_AGEMA_signal_5676, new_AGEMA_signal_5675}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, Midori_rounds_sub_sBox_PRINCE_7_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .a ({new_AGEMA_signal_5680, new_AGEMA_signal_5679, new_AGEMA_signal_5678}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, Midori_rounds_sub_sBox_PRINCE_7_n4}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, Midori_rounds_sub_sBox_PRINCE_7_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .a ({new_AGEMA_signal_5683, new_AGEMA_signal_5682, new_AGEMA_signal_5681}), .b ({new_AGEMA_signal_1987, new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_7_n1}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_rounds_sub_sBox_PRINCE_7_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .a ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_5686, new_AGEMA_signal_5685, new_AGEMA_signal_5684}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, Midori_rounds_sub_sBox_PRINCE_8_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .a ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_8_n10}), .b ({new_AGEMA_signal_5689, new_AGEMA_signal_5688, new_AGEMA_signal_5687}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, Midori_rounds_sub_sBox_PRINCE_8_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .a ({new_AGEMA_signal_5692, new_AGEMA_signal_5691, new_AGEMA_signal_5690}), .b ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, Midori_rounds_sub_sBox_PRINCE_8_n4}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_rounds_sub_sBox_PRINCE_8_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .a ({new_AGEMA_signal_5695, new_AGEMA_signal_5694, new_AGEMA_signal_5693}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_8_n1}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_rounds_sub_sBox_PRINCE_8_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .a ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_5698, new_AGEMA_signal_5697, new_AGEMA_signal_5696}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_rounds_sub_sBox_PRINCE_9_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, Midori_rounds_sub_sBox_PRINCE_9_n10}), .b ({new_AGEMA_signal_5701, new_AGEMA_signal_5700, new_AGEMA_signal_5699}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, Midori_rounds_sub_sBox_PRINCE_9_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .a ({new_AGEMA_signal_5704, new_AGEMA_signal_5703, new_AGEMA_signal_5702}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, Midori_rounds_sub_sBox_PRINCE_9_n4}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, Midori_rounds_sub_sBox_PRINCE_9_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .a ({new_AGEMA_signal_5707, new_AGEMA_signal_5706, new_AGEMA_signal_5705}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, Midori_rounds_sub_sBox_PRINCE_9_n1}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_rounds_sub_sBox_PRINCE_9_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .a ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_5710, new_AGEMA_signal_5709, new_AGEMA_signal_5708}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, Midori_rounds_sub_sBox_PRINCE_10_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, Midori_rounds_sub_sBox_PRINCE_10_n10}), .b ({new_AGEMA_signal_5713, new_AGEMA_signal_5712, new_AGEMA_signal_5711}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, Midori_rounds_sub_sBox_PRINCE_10_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .a ({new_AGEMA_signal_5716, new_AGEMA_signal_5715, new_AGEMA_signal_5714}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, Midori_rounds_sub_sBox_PRINCE_10_n4}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, Midori_rounds_sub_sBox_PRINCE_10_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .a ({new_AGEMA_signal_5719, new_AGEMA_signal_5718, new_AGEMA_signal_5717}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, Midori_rounds_sub_sBox_PRINCE_10_n1}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_rounds_sub_sBox_PRINCE_10_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .a ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_5722, new_AGEMA_signal_5721, new_AGEMA_signal_5720}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, Midori_rounds_sub_sBox_PRINCE_11_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, Midori_rounds_sub_sBox_PRINCE_11_n10}), .b ({new_AGEMA_signal_5725, new_AGEMA_signal_5724, new_AGEMA_signal_5723}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, Midori_rounds_sub_sBox_PRINCE_11_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .a ({new_AGEMA_signal_5728, new_AGEMA_signal_5727, new_AGEMA_signal_5726}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, Midori_rounds_sub_sBox_PRINCE_11_n4}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_rounds_sub_sBox_PRINCE_11_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .a ({new_AGEMA_signal_5731, new_AGEMA_signal_5730, new_AGEMA_signal_5729}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, Midori_rounds_sub_sBox_PRINCE_11_n1}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_rounds_sub_sBox_PRINCE_11_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .a ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_5734, new_AGEMA_signal_5733, new_AGEMA_signal_5732}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_rounds_sub_sBox_PRINCE_12_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, Midori_rounds_sub_sBox_PRINCE_12_n10}), .b ({new_AGEMA_signal_5737, new_AGEMA_signal_5736, new_AGEMA_signal_5735}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, Midori_rounds_sub_sBox_PRINCE_12_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .a ({new_AGEMA_signal_5740, new_AGEMA_signal_5739, new_AGEMA_signal_5738}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, Midori_rounds_sub_sBox_PRINCE_12_n4}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, Midori_rounds_sub_sBox_PRINCE_12_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .a ({new_AGEMA_signal_5743, new_AGEMA_signal_5742, new_AGEMA_signal_5741}), .b ({new_AGEMA_signal_2067, new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_12_n1}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_rounds_sub_sBox_PRINCE_12_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_5746, new_AGEMA_signal_5745, new_AGEMA_signal_5744}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, Midori_rounds_sub_sBox_PRINCE_13_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .a ({new_AGEMA_signal_2079, new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_13_n10}), .b ({new_AGEMA_signal_5749, new_AGEMA_signal_5748, new_AGEMA_signal_5747}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, Midori_rounds_sub_sBox_PRINCE_13_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .a ({new_AGEMA_signal_5752, new_AGEMA_signal_5751, new_AGEMA_signal_5750}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, Midori_rounds_sub_sBox_PRINCE_13_n4}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, Midori_rounds_sub_sBox_PRINCE_13_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .a ({new_AGEMA_signal_5755, new_AGEMA_signal_5754, new_AGEMA_signal_5753}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_13_n1}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_rounds_sub_sBox_PRINCE_13_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .a ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_5758, new_AGEMA_signal_5757, new_AGEMA_signal_5756}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, Midori_rounds_sub_sBox_PRINCE_14_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .a ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, Midori_rounds_sub_sBox_PRINCE_14_n10}), .b ({new_AGEMA_signal_5761, new_AGEMA_signal_5760, new_AGEMA_signal_5759}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, Midori_rounds_sub_sBox_PRINCE_14_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .a ({new_AGEMA_signal_5764, new_AGEMA_signal_5763, new_AGEMA_signal_5762}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, Midori_rounds_sub_sBox_PRINCE_14_n4}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_rounds_sub_sBox_PRINCE_14_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .a ({new_AGEMA_signal_5767, new_AGEMA_signal_5766, new_AGEMA_signal_5765}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_14_n1}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_rounds_sub_sBox_PRINCE_14_n2}) ) ;
    or_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .a ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_5770, new_AGEMA_signal_5769, new_AGEMA_signal_5768}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_rounds_sub_sBox_PRINCE_15_n14}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .a ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_15_n10}), .b ({new_AGEMA_signal_5773, new_AGEMA_signal_5772, new_AGEMA_signal_5771}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, Midori_rounds_sub_sBox_PRINCE_15_n11}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .a ({new_AGEMA_signal_5776, new_AGEMA_signal_5775, new_AGEMA_signal_5774}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, Midori_rounds_sub_sBox_PRINCE_15_n4}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, Midori_rounds_sub_sBox_PRINCE_15_n5}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .a ({new_AGEMA_signal_5779, new_AGEMA_signal_5778, new_AGEMA_signal_5777}), .b ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, Midori_rounds_sub_sBox_PRINCE_15_n1}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_rounds_sub_sBox_PRINCE_15_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (new_AGEMA_signal_5789), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (new_AGEMA_signal_5801), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (new_AGEMA_signal_5813), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (new_AGEMA_signal_5825), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (new_AGEMA_signal_5837), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (new_AGEMA_signal_5849), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (new_AGEMA_signal_5861), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (new_AGEMA_signal_5873), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (new_AGEMA_signal_5885), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (new_AGEMA_signal_5897), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (new_AGEMA_signal_5909), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (new_AGEMA_signal_5933), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_5957), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_5969), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (new_AGEMA_signal_5981), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_5993), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_6005), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (new_AGEMA_signal_6017), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_6029), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_6041), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_6053), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_6065), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_6077), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (new_AGEMA_signal_6089), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_6101), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_6113), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (new_AGEMA_signal_6125), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_6137), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_6149), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (new_AGEMA_signal_6161), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_6173), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_6185), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (new_AGEMA_signal_6197), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_6209), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_6221), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (new_AGEMA_signal_6233), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (new_AGEMA_signal_6239), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_6245), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_6257), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_6266), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (new_AGEMA_signal_6269), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_6281), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (new_AGEMA_signal_6287), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_6290), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_6293), .Q (new_AGEMA_signal_6294) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (new_AGEMA_signal_6299), .Q (new_AGEMA_signal_6300) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_6303) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (new_AGEMA_signal_6305), .Q (new_AGEMA_signal_6306) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_6312) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_6314), .Q (new_AGEMA_signal_6315) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_6317), .Q (new_AGEMA_signal_6318) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_6321) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_6324) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_6327) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_6329), .Q (new_AGEMA_signal_6330) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_6333) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_6336) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_6338), .Q (new_AGEMA_signal_6339) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_6341), .Q (new_AGEMA_signal_6342) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_6345) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (new_AGEMA_signal_6347), .Q (new_AGEMA_signal_6348) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_6351) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_6353), .Q (new_AGEMA_signal_6354) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_6360) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_6363) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_6365), .Q (new_AGEMA_signal_6366) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_6369) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (new_AGEMA_signal_6371), .Q (new_AGEMA_signal_6372) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_6375) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_6377), .Q (new_AGEMA_signal_6378) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_6381) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_6384) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_6387) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_6389), .Q (new_AGEMA_signal_6390) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_6393) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_6396) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_6399) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_6401), .Q (new_AGEMA_signal_6402) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_6408) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_6411) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_6413), .Q (new_AGEMA_signal_6414) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_6417) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_6419), .Q (new_AGEMA_signal_6420) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_6423) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_6425), .Q (new_AGEMA_signal_6426) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_6429) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_6432) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_6435) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_6437), .Q (new_AGEMA_signal_6438) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_6441) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_6443), .Q (new_AGEMA_signal_6444) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_6447) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (new_AGEMA_signal_6449), .Q (new_AGEMA_signal_6450) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_6455), .Q (new_AGEMA_signal_6456) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_6459) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_6462) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_6465) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_6467), .Q (new_AGEMA_signal_6468) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_6471) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_6473), .Q (new_AGEMA_signal_6474) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_6477) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_6479), .Q (new_AGEMA_signal_6480) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_6483) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (new_AGEMA_signal_6485), .Q (new_AGEMA_signal_6486) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_6489) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_6491), .Q (new_AGEMA_signal_6492) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_6495) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_6497), .Q (new_AGEMA_signal_6498) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_6503), .Q (new_AGEMA_signal_6504) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_6507) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_6509), .Q (new_AGEMA_signal_6510) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_6513) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_6515), .Q (new_AGEMA_signal_6516) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_6519) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (new_AGEMA_signal_6521), .Q (new_AGEMA_signal_6522) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_6525) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_6527), .Q (new_AGEMA_signal_6528) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_6530), .Q (new_AGEMA_signal_6531) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_6533), .Q (new_AGEMA_signal_6534) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_6537) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_6539), .Q (new_AGEMA_signal_6540) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_6543) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_6545), .Q (new_AGEMA_signal_6546) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_6551), .Q (new_AGEMA_signal_6552) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_6554), .Q (new_AGEMA_signal_6555) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (new_AGEMA_signal_6557), .Q (new_AGEMA_signal_6558) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_6561) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_6563), .Q (new_AGEMA_signal_6564) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_6566), .Q (new_AGEMA_signal_6567) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_6569), .Q (new_AGEMA_signal_6570) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_6572), .Q (new_AGEMA_signal_6573) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_6575), .Q (new_AGEMA_signal_6576) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_6578), .Q (new_AGEMA_signal_6579) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_6581), .Q (new_AGEMA_signal_6582) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_6584), .Q (new_AGEMA_signal_6585) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_6587), .Q (new_AGEMA_signal_6588) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_6590), .Q (new_AGEMA_signal_6591) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (new_AGEMA_signal_6593), .Q (new_AGEMA_signal_6594) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_6597) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_6599), .Q (new_AGEMA_signal_6600) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_6602), .Q (new_AGEMA_signal_6603) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_6605), .Q (new_AGEMA_signal_6606) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_6608), .Q (new_AGEMA_signal_6609) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_6611), .Q (new_AGEMA_signal_6612) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_6614), .Q (new_AGEMA_signal_6615) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_6617), .Q (new_AGEMA_signal_6618) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_6620), .Q (new_AGEMA_signal_6621) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_6623), .Q (new_AGEMA_signal_6624) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_6626), .Q (new_AGEMA_signal_6627) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (new_AGEMA_signal_6629), .Q (new_AGEMA_signal_6630) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_6633) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_6635), .Q (new_AGEMA_signal_6636) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_6638), .Q (new_AGEMA_signal_6639) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_6641), .Q (new_AGEMA_signal_6642) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_6644), .Q (new_AGEMA_signal_6645) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n15), .Q (new_AGEMA_signal_6647) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_2380), .Q (new_AGEMA_signal_6648) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_2381), .Q (new_AGEMA_signal_6649) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_6650) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_6651) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_6652) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n6), .Q (new_AGEMA_signal_6653) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_2384), .Q (new_AGEMA_signal_6654) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_2385), .Q (new_AGEMA_signal_6655) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n15), .Q (new_AGEMA_signal_6656) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_2392), .Q (new_AGEMA_signal_6657) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_2393), .Q (new_AGEMA_signal_6658) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_6659) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_6660) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_6661) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n6), .Q (new_AGEMA_signal_6662) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_2396), .Q (new_AGEMA_signal_6663) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_2397), .Q (new_AGEMA_signal_6664) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n15), .Q (new_AGEMA_signal_6665) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (new_AGEMA_signal_2404), .Q (new_AGEMA_signal_6666) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_6667) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_6668) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_5613), .Q (new_AGEMA_signal_6669) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_6670) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n6), .Q (new_AGEMA_signal_6671) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_2408), .Q (new_AGEMA_signal_6672) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_2409), .Q (new_AGEMA_signal_6673) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n15), .Q (new_AGEMA_signal_6674) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_2416), .Q (new_AGEMA_signal_6675) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_2417), .Q (new_AGEMA_signal_6676) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_6677) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_6678) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_6679) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n6), .Q (new_AGEMA_signal_6680) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_2420), .Q (new_AGEMA_signal_6681) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_2421), .Q (new_AGEMA_signal_6682) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n15), .Q (new_AGEMA_signal_6683) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_2428), .Q (new_AGEMA_signal_6684) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_2429), .Q (new_AGEMA_signal_6685) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_6686) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_6687) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_6688) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n6), .Q (new_AGEMA_signal_6689) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_2432), .Q (new_AGEMA_signal_6690) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_2433), .Q (new_AGEMA_signal_6691) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n15), .Q (new_AGEMA_signal_6692) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_2440), .Q (new_AGEMA_signal_6693) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_6694) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_6695) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_5649), .Q (new_AGEMA_signal_6696) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_6697) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n6), .Q (new_AGEMA_signal_6698) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_2444), .Q (new_AGEMA_signal_6699) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_2445), .Q (new_AGEMA_signal_6700) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n15), .Q (new_AGEMA_signal_6701) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (new_AGEMA_signal_2452), .Q (new_AGEMA_signal_6702) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_2453), .Q (new_AGEMA_signal_6703) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_6704) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_6705) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_6706) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n6), .Q (new_AGEMA_signal_6707) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_6708) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_2457), .Q (new_AGEMA_signal_6709) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n15), .Q (new_AGEMA_signal_6710) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_2464), .Q (new_AGEMA_signal_6711) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_2465), .Q (new_AGEMA_signal_6712) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_6713) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (new_AGEMA_signal_5673), .Q (new_AGEMA_signal_6714) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_5674), .Q (new_AGEMA_signal_6715) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n6), .Q (new_AGEMA_signal_6716) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_6717) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_2469), .Q (new_AGEMA_signal_6718) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n15), .Q (new_AGEMA_signal_6719) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_2476), .Q (new_AGEMA_signal_6720) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_2477), .Q (new_AGEMA_signal_6721) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_6722) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_5685), .Q (new_AGEMA_signal_6723) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_6724) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n6), .Q (new_AGEMA_signal_6725) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_2480), .Q (new_AGEMA_signal_6726) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_2481), .Q (new_AGEMA_signal_6727) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n15), .Q (new_AGEMA_signal_6728) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_2488), .Q (new_AGEMA_signal_6729) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_2489), .Q (new_AGEMA_signal_6730) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_6731) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_6732) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_6733) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n6), .Q (new_AGEMA_signal_6734) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_2492), .Q (new_AGEMA_signal_6735) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_2493), .Q (new_AGEMA_signal_6736) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n15), .Q (new_AGEMA_signal_6737) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (new_AGEMA_signal_2500), .Q (new_AGEMA_signal_6738) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_2501), .Q (new_AGEMA_signal_6739) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_6740) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_6741) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_6742) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n6), .Q (new_AGEMA_signal_6743) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_2504), .Q (new_AGEMA_signal_6744) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_2505), .Q (new_AGEMA_signal_6745) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n15), .Q (new_AGEMA_signal_6746) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_2512), .Q (new_AGEMA_signal_6747) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_2513), .Q (new_AGEMA_signal_6748) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_6749) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_6750) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_6751) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n6), .Q (new_AGEMA_signal_6752) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_2516), .Q (new_AGEMA_signal_6753) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_2517), .Q (new_AGEMA_signal_6754) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n15), .Q (new_AGEMA_signal_6755) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_2524), .Q (new_AGEMA_signal_6756) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_2525), .Q (new_AGEMA_signal_6757) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_6758) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_5733), .Q (new_AGEMA_signal_6759) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_6760) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n6), .Q (new_AGEMA_signal_6761) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_2528), .Q (new_AGEMA_signal_6762) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_2529), .Q (new_AGEMA_signal_6763) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n15), .Q (new_AGEMA_signal_6764) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_2536), .Q (new_AGEMA_signal_6765) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_2537), .Q (new_AGEMA_signal_6766) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_6767) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_5745), .Q (new_AGEMA_signal_6768) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_6769) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n6), .Q (new_AGEMA_signal_6770) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_2540), .Q (new_AGEMA_signal_6771) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_2541), .Q (new_AGEMA_signal_6772) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n15), .Q (new_AGEMA_signal_6773) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (new_AGEMA_signal_2548), .Q (new_AGEMA_signal_6774) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_2549), .Q (new_AGEMA_signal_6775) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_6776) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_5757), .Q (new_AGEMA_signal_6777) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_6778) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n6), .Q (new_AGEMA_signal_6779) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_2552), .Q (new_AGEMA_signal_6780) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_2553), .Q (new_AGEMA_signal_6781) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n15), .Q (new_AGEMA_signal_6782) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_2560), .Q (new_AGEMA_signal_6783) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_2561), .Q (new_AGEMA_signal_6784) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_6785) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_6786) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_6787) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n6), .Q (new_AGEMA_signal_6788) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_2564), .Q (new_AGEMA_signal_6789) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_2565), .Q (new_AGEMA_signal_6790) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_6791), .Q (new_AGEMA_signal_6792) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_6794), .Q (new_AGEMA_signal_6795) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_6798), .Q (new_AGEMA_signal_6799) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_6802), .Q (new_AGEMA_signal_6803) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_6806), .Q (new_AGEMA_signal_6807) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_6810), .Q (new_AGEMA_signal_6811) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_6814), .Q (new_AGEMA_signal_6815) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_6818), .Q (new_AGEMA_signal_6819) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_6822), .Q (new_AGEMA_signal_6823) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_6826), .Q (new_AGEMA_signal_6827) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_6830), .Q (new_AGEMA_signal_6831) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_6834), .Q (new_AGEMA_signal_6835) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_6838), .Q (new_AGEMA_signal_6839) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_6842), .Q (new_AGEMA_signal_6843) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_6846), .Q (new_AGEMA_signal_6847) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_6850), .Q (new_AGEMA_signal_6851) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_6854), .Q (new_AGEMA_signal_6855) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_6858), .Q (new_AGEMA_signal_6859) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_6862), .Q (new_AGEMA_signal_6863) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_6866), .Q (new_AGEMA_signal_6867) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_6870), .Q (new_AGEMA_signal_6871) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_6874), .Q (new_AGEMA_signal_6875) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_6878), .Q (new_AGEMA_signal_6879) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_6882), .Q (new_AGEMA_signal_6883) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_6886), .Q (new_AGEMA_signal_6887) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_6890), .Q (new_AGEMA_signal_6891) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_6894), .Q (new_AGEMA_signal_6895) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_6898), .Q (new_AGEMA_signal_6899) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_6902), .Q (new_AGEMA_signal_6903) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_6906), .Q (new_AGEMA_signal_6907) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_6910), .Q (new_AGEMA_signal_6911) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_6914), .Q (new_AGEMA_signal_6915) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_6918), .Q (new_AGEMA_signal_6919) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_6922), .Q (new_AGEMA_signal_6923) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_6926), .Q (new_AGEMA_signal_6927) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_6930), .Q (new_AGEMA_signal_6931) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_6934), .Q (new_AGEMA_signal_6935) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_6938), .Q (new_AGEMA_signal_6939) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_6942), .Q (new_AGEMA_signal_6943) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_6946), .Q (new_AGEMA_signal_6947) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_6950), .Q (new_AGEMA_signal_6951) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_6954), .Q (new_AGEMA_signal_6955) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_6958), .Q (new_AGEMA_signal_6959) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_6962), .Q (new_AGEMA_signal_6963) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_6966), .Q (new_AGEMA_signal_6967) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_6970), .Q (new_AGEMA_signal_6971) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_6974), .Q (new_AGEMA_signal_6975) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_6978), .Q (new_AGEMA_signal_6979) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_6982), .Q (new_AGEMA_signal_6983) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_6986), .Q (new_AGEMA_signal_6987) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_6990), .Q (new_AGEMA_signal_6991) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_6994), .Q (new_AGEMA_signal_6995) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_6998), .Q (new_AGEMA_signal_6999) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_7002), .Q (new_AGEMA_signal_7003) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_7006), .Q (new_AGEMA_signal_7007) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_7010), .Q (new_AGEMA_signal_7011) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_7014), .Q (new_AGEMA_signal_7015) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_7018), .Q (new_AGEMA_signal_7019) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_7022), .Q (new_AGEMA_signal_7023) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_7026), .Q (new_AGEMA_signal_7027) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_7030), .Q (new_AGEMA_signal_7031) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_7034), .Q (new_AGEMA_signal_7035) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_7038), .Q (new_AGEMA_signal_7039) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_7042), .Q (new_AGEMA_signal_7043) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_7046), .Q (new_AGEMA_signal_7047) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_7050), .Q (new_AGEMA_signal_7051) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_7054), .Q (new_AGEMA_signal_7055) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_7058), .Q (new_AGEMA_signal_7059) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_7062), .Q (new_AGEMA_signal_7063) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_7066), .Q (new_AGEMA_signal_7067) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_7070), .Q (new_AGEMA_signal_7071) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_7074), .Q (new_AGEMA_signal_7075) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_7078), .Q (new_AGEMA_signal_7079) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_7082), .Q (new_AGEMA_signal_7083) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_7086), .Q (new_AGEMA_signal_7087) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_7090), .Q (new_AGEMA_signal_7091) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_7094), .Q (new_AGEMA_signal_7095) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_7098), .Q (new_AGEMA_signal_7099) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_7102), .Q (new_AGEMA_signal_7103) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_7106), .Q (new_AGEMA_signal_7107) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_7110), .Q (new_AGEMA_signal_7111) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_7114), .Q (new_AGEMA_signal_7115) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_7118), .Q (new_AGEMA_signal_7119) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_7122), .Q (new_AGEMA_signal_7123) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_7126), .Q (new_AGEMA_signal_7127) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_7130), .Q (new_AGEMA_signal_7131) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_7134), .Q (new_AGEMA_signal_7135) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_7138), .Q (new_AGEMA_signal_7139) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_7142), .Q (new_AGEMA_signal_7143) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_7146), .Q (new_AGEMA_signal_7147) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_7150), .Q (new_AGEMA_signal_7151) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_7154), .Q (new_AGEMA_signal_7155) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_7158), .Q (new_AGEMA_signal_7159) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_7162), .Q (new_AGEMA_signal_7163) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_7166), .Q (new_AGEMA_signal_7167) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_7170), .Q (new_AGEMA_signal_7171) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_7174), .Q (new_AGEMA_signal_7175) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_7178), .Q (new_AGEMA_signal_7179) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_7182), .Q (new_AGEMA_signal_7183) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_7187) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_7190), .Q (new_AGEMA_signal_7191) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_7194), .Q (new_AGEMA_signal_7195) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_7198), .Q (new_AGEMA_signal_7199) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_7202), .Q (new_AGEMA_signal_7203) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_7206), .Q (new_AGEMA_signal_7207) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_7210), .Q (new_AGEMA_signal_7211) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_7214), .Q (new_AGEMA_signal_7215) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_7218), .Q (new_AGEMA_signal_7219) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_7222), .Q (new_AGEMA_signal_7223) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_7226), .Q (new_AGEMA_signal_7227) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_7230), .Q (new_AGEMA_signal_7231) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_7234), .Q (new_AGEMA_signal_7235) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_7238), .Q (new_AGEMA_signal_7239) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_7242), .Q (new_AGEMA_signal_7243) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_7246), .Q (new_AGEMA_signal_7247) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_7250), .Q (new_AGEMA_signal_7251) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_7254), .Q (new_AGEMA_signal_7255) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_7258), .Q (new_AGEMA_signal_7259) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_7262), .Q (new_AGEMA_signal_7263) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_7266), .Q (new_AGEMA_signal_7267) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_7270), .Q (new_AGEMA_signal_7271) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_7274), .Q (new_AGEMA_signal_7275) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_7278), .Q (new_AGEMA_signal_7279) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_7282), .Q (new_AGEMA_signal_7283) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_7286), .Q (new_AGEMA_signal_7287) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_7290), .Q (new_AGEMA_signal_7291) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_7294), .Q (new_AGEMA_signal_7295) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_7298), .Q (new_AGEMA_signal_7299) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_7302), .Q (new_AGEMA_signal_7303) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_7306), .Q (new_AGEMA_signal_7307) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_7310), .Q (new_AGEMA_signal_7311) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_7314), .Q (new_AGEMA_signal_7315) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_7318), .Q (new_AGEMA_signal_7319) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_7322), .Q (new_AGEMA_signal_7323) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_7326), .Q (new_AGEMA_signal_7327) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_7330), .Q (new_AGEMA_signal_7331) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_7334), .Q (new_AGEMA_signal_7335) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_7338), .Q (new_AGEMA_signal_7339) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_7342), .Q (new_AGEMA_signal_7343) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_7346), .Q (new_AGEMA_signal_7347) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_7350), .Q (new_AGEMA_signal_7351) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_7354), .Q (new_AGEMA_signal_7355) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_7358), .Q (new_AGEMA_signal_7359) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_7362), .Q (new_AGEMA_signal_7363) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_7366), .Q (new_AGEMA_signal_7367) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_7370), .Q (new_AGEMA_signal_7371) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_7374), .Q (new_AGEMA_signal_7375) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_7378), .Q (new_AGEMA_signal_7379) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_7382), .Q (new_AGEMA_signal_7383) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_7386), .Q (new_AGEMA_signal_7387) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_7390), .Q (new_AGEMA_signal_7391) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_7394), .Q (new_AGEMA_signal_7395) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_7398), .Q (new_AGEMA_signal_7399) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_7402), .Q (new_AGEMA_signal_7403) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_7406), .Q (new_AGEMA_signal_7407) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_7410), .Q (new_AGEMA_signal_7411) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_7414), .Q (new_AGEMA_signal_7415) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_7418), .Q (new_AGEMA_signal_7419) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_7422), .Q (new_AGEMA_signal_7423) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_7426), .Q (new_AGEMA_signal_7427) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_7430), .Q (new_AGEMA_signal_7431) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_7434), .Q (new_AGEMA_signal_7435) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_7438), .Q (new_AGEMA_signal_7439) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_7442), .Q (new_AGEMA_signal_7443) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_7447) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_7450), .Q (new_AGEMA_signal_7451) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_7454), .Q (new_AGEMA_signal_7455) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_7458), .Q (new_AGEMA_signal_7459) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_7462), .Q (new_AGEMA_signal_7463) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_7466), .Q (new_AGEMA_signal_7467) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_7470), .Q (new_AGEMA_signal_7471) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_7474), .Q (new_AGEMA_signal_7475) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_7478), .Q (new_AGEMA_signal_7479) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_7482), .Q (new_AGEMA_signal_7483) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_7487) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_7490), .Q (new_AGEMA_signal_7491) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_7494), .Q (new_AGEMA_signal_7495) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_7498), .Q (new_AGEMA_signal_7499) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_7502), .Q (new_AGEMA_signal_7503) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_7506), .Q (new_AGEMA_signal_7507) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_7510), .Q (new_AGEMA_signal_7511) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_7514), .Q (new_AGEMA_signal_7515) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_7518), .Q (new_AGEMA_signal_7519) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_7522), .Q (new_AGEMA_signal_7523) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_7526), .Q (new_AGEMA_signal_7527) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_7530), .Q (new_AGEMA_signal_7531) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_7534), .Q (new_AGEMA_signal_7535) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_7538), .Q (new_AGEMA_signal_7539) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_7542), .Q (new_AGEMA_signal_7543) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_7546), .Q (new_AGEMA_signal_7547) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_7550), .Q (new_AGEMA_signal_7551) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_7554), .Q (new_AGEMA_signal_7555) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_7558), .Q (new_AGEMA_signal_7559) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_7563), .Q (new_AGEMA_signal_7564) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_7567), .Q (new_AGEMA_signal_7568) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (new_AGEMA_signal_7571), .Q (new_AGEMA_signal_7572) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_7575), .Q (new_AGEMA_signal_7576) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_7579), .Q (new_AGEMA_signal_7580) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_7583), .Q (new_AGEMA_signal_7584) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_7587), .Q (new_AGEMA_signal_7588) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_7591), .Q (new_AGEMA_signal_7592) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_7595), .Q (new_AGEMA_signal_7596) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_7599), .Q (new_AGEMA_signal_7600) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_7603), .Q (new_AGEMA_signal_7604) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_7607), .Q (new_AGEMA_signal_7608) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_7611), .Q (new_AGEMA_signal_7612) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_7616) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_7619), .Q (new_AGEMA_signal_7620) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_7623), .Q (new_AGEMA_signal_7624) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_7627), .Q (new_AGEMA_signal_7628) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_7631), .Q (new_AGEMA_signal_7632) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_7635), .Q (new_AGEMA_signal_7636) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_7639), .Q (new_AGEMA_signal_7640) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_7643), .Q (new_AGEMA_signal_7644) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_7647), .Q (new_AGEMA_signal_7648) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_7651), .Q (new_AGEMA_signal_7652) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_7655), .Q (new_AGEMA_signal_7656) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_7659), .Q (new_AGEMA_signal_7660) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_7663), .Q (new_AGEMA_signal_7664) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_7667), .Q (new_AGEMA_signal_7668) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_7671), .Q (new_AGEMA_signal_7672) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_7675), .Q (new_AGEMA_signal_7676) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_7679), .Q (new_AGEMA_signal_7680) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_7683), .Q (new_AGEMA_signal_7684) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_7687), .Q (new_AGEMA_signal_7688) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_7691), .Q (new_AGEMA_signal_7692) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_7695), .Q (new_AGEMA_signal_7696) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_7699), .Q (new_AGEMA_signal_7700) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_7703), .Q (new_AGEMA_signal_7704) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_7707), .Q (new_AGEMA_signal_7708) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_7711), .Q (new_AGEMA_signal_7712) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_7715), .Q (new_AGEMA_signal_7716) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_7719), .Q (new_AGEMA_signal_7720) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_7723), .Q (new_AGEMA_signal_7724) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_7727), .Q (new_AGEMA_signal_7728) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_7731), .Q (new_AGEMA_signal_7732) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_7735), .Q (new_AGEMA_signal_7736) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_7739), .Q (new_AGEMA_signal_7740) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_7743), .Q (new_AGEMA_signal_7744) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_7747), .Q (new_AGEMA_signal_7748) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_7751), .Q (new_AGEMA_signal_7752) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_7755), .Q (new_AGEMA_signal_7756) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_7759), .Q (new_AGEMA_signal_7760) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_7763), .Q (new_AGEMA_signal_7764) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_7767), .Q (new_AGEMA_signal_7768) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_7771), .Q (new_AGEMA_signal_7772) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_7775), .Q (new_AGEMA_signal_7776) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_7779), .Q (new_AGEMA_signal_7780) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_7783), .Q (new_AGEMA_signal_7784) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_7787), .Q (new_AGEMA_signal_7788) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_7791), .Q (new_AGEMA_signal_7792) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_7795), .Q (new_AGEMA_signal_7796) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_7799), .Q (new_AGEMA_signal_7800) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_7803), .Q (new_AGEMA_signal_7804) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_7807), .Q (new_AGEMA_signal_7808) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_7811), .Q (new_AGEMA_signal_7812) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_7815), .Q (new_AGEMA_signal_7816) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_7819), .Q (new_AGEMA_signal_7820) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_7823), .Q (new_AGEMA_signal_7824) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_7827), .Q (new_AGEMA_signal_7828) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_7831), .Q (new_AGEMA_signal_7832) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_7835), .Q (new_AGEMA_signal_7836) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_7839), .Q (new_AGEMA_signal_7840) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_7843), .Q (new_AGEMA_signal_7844) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_7847), .Q (new_AGEMA_signal_7848) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_7851), .Q (new_AGEMA_signal_7852) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_7855), .Q (new_AGEMA_signal_7856) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_7859), .Q (new_AGEMA_signal_7860) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_7863), .Q (new_AGEMA_signal_7864) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_7867), .Q (new_AGEMA_signal_7868) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_7871), .Q (new_AGEMA_signal_7872) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_7875), .Q (new_AGEMA_signal_7876) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_7879), .Q (new_AGEMA_signal_7880) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_7883), .Q (new_AGEMA_signal_7884) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_7887), .Q (new_AGEMA_signal_7888) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_7891), .Q (new_AGEMA_signal_7892) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_7895), .Q (new_AGEMA_signal_7896) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_7899), .Q (new_AGEMA_signal_7900) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_7903), .Q (new_AGEMA_signal_7904) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_7907), .Q (new_AGEMA_signal_7908) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_7911), .Q (new_AGEMA_signal_7912) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_7915), .Q (new_AGEMA_signal_7916) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_7919), .Q (new_AGEMA_signal_7920) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_7923), .Q (new_AGEMA_signal_7924) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_7927), .Q (new_AGEMA_signal_7928) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_7931), .Q (new_AGEMA_signal_7932) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_7935), .Q (new_AGEMA_signal_7936) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_7939), .Q (new_AGEMA_signal_7940) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_7943), .Q (new_AGEMA_signal_7944) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n13), .Q (new_AGEMA_signal_7950) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_7952) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_2389), .Q (new_AGEMA_signal_7954) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n13), .Q (new_AGEMA_signal_7959) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_7961) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_2401), .Q (new_AGEMA_signal_7963) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n13), .Q (new_AGEMA_signal_7968) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_2412), .Q (new_AGEMA_signal_7970) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_2413), .Q (new_AGEMA_signal_7972) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n13), .Q (new_AGEMA_signal_7977) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_2424), .Q (new_AGEMA_signal_7979) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_2425), .Q (new_AGEMA_signal_7981) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n13), .Q (new_AGEMA_signal_7986) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_2436), .Q (new_AGEMA_signal_7988) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_2437), .Q (new_AGEMA_signal_7990) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n13), .Q (new_AGEMA_signal_7995) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_2448), .Q (new_AGEMA_signal_7997) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_2449), .Q (new_AGEMA_signal_7999) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n13), .Q (new_AGEMA_signal_8004) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_8006) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_2461), .Q (new_AGEMA_signal_8008) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n13), .Q (new_AGEMA_signal_8013) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_2472), .Q (new_AGEMA_signal_8015) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_2473), .Q (new_AGEMA_signal_8017) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n13), .Q (new_AGEMA_signal_8022) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_8024) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_2485), .Q (new_AGEMA_signal_8026) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n13), .Q (new_AGEMA_signal_8031) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_8033) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_8035) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n13), .Q (new_AGEMA_signal_8040) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_8042) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_2509), .Q (new_AGEMA_signal_8044) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n13), .Q (new_AGEMA_signal_8049) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_2520), .Q (new_AGEMA_signal_8051) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_2521), .Q (new_AGEMA_signal_8053) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n13), .Q (new_AGEMA_signal_8058) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_2532), .Q (new_AGEMA_signal_8060) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_2533), .Q (new_AGEMA_signal_8062) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n13), .Q (new_AGEMA_signal_8067) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_2544), .Q (new_AGEMA_signal_8069) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_2545), .Q (new_AGEMA_signal_8071) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n13), .Q (new_AGEMA_signal_8076) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_2556), .Q (new_AGEMA_signal_8078) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_2557), .Q (new_AGEMA_signal_8080) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n13), .Q (new_AGEMA_signal_8085) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_2568), .Q (new_AGEMA_signal_8087) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_2569), .Q (new_AGEMA_signal_8089) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_8092), .Q (new_AGEMA_signal_8093) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_8096), .Q (new_AGEMA_signal_8097) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_8100), .Q (new_AGEMA_signal_8101) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_8104), .Q (new_AGEMA_signal_8105) ) ;

    /* cells in depth 3 */
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U128 ( .a ({new_AGEMA_signal_5788, new_AGEMA_signal_5785, new_AGEMA_signal_5782}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_5525, new_AGEMA_signal_5524, new_AGEMA_signal_5515}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U126 ( .a ({new_AGEMA_signal_5797, new_AGEMA_signal_5794, new_AGEMA_signal_5791}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_5527, new_AGEMA_signal_5526, new_AGEMA_signal_5516}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U124 ( .a ({new_AGEMA_signal_5806, new_AGEMA_signal_5803, new_AGEMA_signal_5800}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_5529, new_AGEMA_signal_5528, new_AGEMA_signal_5488}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U122 ( .a ({new_AGEMA_signal_5815, new_AGEMA_signal_5812, new_AGEMA_signal_5809}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_5531, new_AGEMA_signal_5530, new_AGEMA_signal_5489}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U120 ( .a ({new_AGEMA_signal_5824, new_AGEMA_signal_5821, new_AGEMA_signal_5818}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_5533, new_AGEMA_signal_5532, new_AGEMA_signal_5517}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U119 ( .a ({new_AGEMA_signal_5833, new_AGEMA_signal_5830, new_AGEMA_signal_5827}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5490}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U117 ( .a ({new_AGEMA_signal_5842, new_AGEMA_signal_5839, new_AGEMA_signal_5836}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_5537, new_AGEMA_signal_5536, new_AGEMA_signal_5491}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U115 ( .a ({new_AGEMA_signal_5851, new_AGEMA_signal_5848, new_AGEMA_signal_5845}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_5539, new_AGEMA_signal_5538, new_AGEMA_signal_5492}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U113 ( .a ({new_AGEMA_signal_5860, new_AGEMA_signal_5857, new_AGEMA_signal_5854}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5493}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U111 ( .a ({new_AGEMA_signal_5869, new_AGEMA_signal_5866, new_AGEMA_signal_5863}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_5543, new_AGEMA_signal_5542, new_AGEMA_signal_5494}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U108 ( .a ({new_AGEMA_signal_5878, new_AGEMA_signal_5875, new_AGEMA_signal_5872}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_5545, new_AGEMA_signal_5544, new_AGEMA_signal_5495}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U106 ( .a ({new_AGEMA_signal_5887, new_AGEMA_signal_5884, new_AGEMA_signal_5881}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_5547, new_AGEMA_signal_5546, new_AGEMA_signal_5496}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U104 ( .a ({new_AGEMA_signal_5896, new_AGEMA_signal_5893, new_AGEMA_signal_5890}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_5549, new_AGEMA_signal_5548, new_AGEMA_signal_5497}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U102 ( .a ({new_AGEMA_signal_5905, new_AGEMA_signal_5902, new_AGEMA_signal_5899}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_5551, new_AGEMA_signal_5550, new_AGEMA_signal_5498}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U100 ( .a ({new_AGEMA_signal_5914, new_AGEMA_signal_5911, new_AGEMA_signal_5908}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5499}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U98 ( .a ({new_AGEMA_signal_5923, new_AGEMA_signal_5920, new_AGEMA_signal_5917}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_5555, new_AGEMA_signal_5554, new_AGEMA_signal_5518}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U97 ( .a ({new_AGEMA_signal_5932, new_AGEMA_signal_5929, new_AGEMA_signal_5926}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_5557, new_AGEMA_signal_5556, new_AGEMA_signal_5500}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U95 ( .a ({new_AGEMA_signal_5941, new_AGEMA_signal_5938, new_AGEMA_signal_5935}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5501}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U93 ( .a ({new_AGEMA_signal_5950, new_AGEMA_signal_5947, new_AGEMA_signal_5944}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_5561, new_AGEMA_signal_5560, new_AGEMA_signal_5502}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U91 ( .a ({new_AGEMA_signal_5959, new_AGEMA_signal_5956, new_AGEMA_signal_5953}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_5563, new_AGEMA_signal_5562, new_AGEMA_signal_5503}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U89 ( .a ({new_AGEMA_signal_5968, new_AGEMA_signal_5965, new_AGEMA_signal_5962}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_5565, new_AGEMA_signal_5564, new_AGEMA_signal_5504}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U86 ( .a ({new_AGEMA_signal_5977, new_AGEMA_signal_5974, new_AGEMA_signal_5971}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_5567, new_AGEMA_signal_5566, new_AGEMA_signal_5505}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U84 ( .a ({new_AGEMA_signal_5986, new_AGEMA_signal_5983, new_AGEMA_signal_5980}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_5569, new_AGEMA_signal_5568, new_AGEMA_signal_5506}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U82 ( .a ({new_AGEMA_signal_5995, new_AGEMA_signal_5992, new_AGEMA_signal_5989}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5507}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U80 ( .a ({new_AGEMA_signal_6004, new_AGEMA_signal_6001, new_AGEMA_signal_5998}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_5573, new_AGEMA_signal_5572, new_AGEMA_signal_5508}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U78 ( .a ({new_AGEMA_signal_6013, new_AGEMA_signal_6010, new_AGEMA_signal_6007}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_5575, new_AGEMA_signal_5574, new_AGEMA_signal_5509}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U76 ( .a ({new_AGEMA_signal_6022, new_AGEMA_signal_6019, new_AGEMA_signal_6016}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5519}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U75 ( .a ({new_AGEMA_signal_6031, new_AGEMA_signal_6028, new_AGEMA_signal_6025}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_5579, new_AGEMA_signal_5578, new_AGEMA_signal_5510}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U73 ( .a ({new_AGEMA_signal_6040, new_AGEMA_signal_6037, new_AGEMA_signal_6034}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_5581, new_AGEMA_signal_5580, new_AGEMA_signal_5511}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U71 ( .a ({new_AGEMA_signal_6049, new_AGEMA_signal_6046, new_AGEMA_signal_6043}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_5583, new_AGEMA_signal_5582, new_AGEMA_signal_5512}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U69 ( .a ({new_AGEMA_signal_6058, new_AGEMA_signal_6055, new_AGEMA_signal_6052}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_5585, new_AGEMA_signal_5584, new_AGEMA_signal_5513}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U67 ( .a ({new_AGEMA_signal_6067, new_AGEMA_signal_6064, new_AGEMA_signal_6061}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_5587, new_AGEMA_signal_5586, new_AGEMA_signal_5514}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U144 ( .a ({new_AGEMA_signal_6076, new_AGEMA_signal_6073, new_AGEMA_signal_6070}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_ResultXORkey[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U142 ( .a ({new_AGEMA_signal_6085, new_AGEMA_signal_6082, new_AGEMA_signal_6079}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, Midori_rounds_sub_ResultXORkey[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U140 ( .a ({new_AGEMA_signal_6094, new_AGEMA_signal_6091, new_AGEMA_signal_6088}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_ResultXORkey[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U138 ( .a ({new_AGEMA_signal_6103, new_AGEMA_signal_6100, new_AGEMA_signal_6097}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, Midori_rounds_sub_ResultXORkey[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U136 ( .a ({new_AGEMA_signal_6112, new_AGEMA_signal_6109, new_AGEMA_signal_6106}), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_ResultXORkey[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U135 ( .a ({new_AGEMA_signal_6121, new_AGEMA_signal_6118, new_AGEMA_signal_6115}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, Midori_rounds_sub_ResultXORkey[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U133 ( .a ({new_AGEMA_signal_6130, new_AGEMA_signal_6127, new_AGEMA_signal_6124}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_ResultXORkey[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U131 ( .a ({new_AGEMA_signal_6139, new_AGEMA_signal_6136, new_AGEMA_signal_6133}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, Midori_rounds_sub_ResultXORkey[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U129 ( .a ({new_AGEMA_signal_6148, new_AGEMA_signal_6145, new_AGEMA_signal_6142}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_ResultXORkey[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U127 ( .a ({new_AGEMA_signal_6157, new_AGEMA_signal_6154, new_AGEMA_signal_6151}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, Midori_rounds_sub_ResultXORkey[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U124 ( .a ({new_AGEMA_signal_6166, new_AGEMA_signal_6163, new_AGEMA_signal_6160}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_ResultXORkey[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U122 ( .a ({new_AGEMA_signal_6175, new_AGEMA_signal_6172, new_AGEMA_signal_6169}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, Midori_rounds_sub_ResultXORkey[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U120 ( .a ({new_AGEMA_signal_6184, new_AGEMA_signal_6181, new_AGEMA_signal_6178}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_ResultXORkey[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U118 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6190, new_AGEMA_signal_6187}), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, Midori_rounds_sub_ResultXORkey[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U116 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6199, new_AGEMA_signal_6196}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_sub_ResultXORkey[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U114 ( .a ({new_AGEMA_signal_6211, new_AGEMA_signal_6208, new_AGEMA_signal_6205}), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, Midori_rounds_sub_ResultXORkey[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U113 ( .a ({new_AGEMA_signal_6220, new_AGEMA_signal_6217, new_AGEMA_signal_6214}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, Midori_rounds_sub_ResultXORkey[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U111 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6226, new_AGEMA_signal_6223}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, Midori_rounds_sub_ResultXORkey[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U109 ( .a ({new_AGEMA_signal_6238, new_AGEMA_signal_6235, new_AGEMA_signal_6232}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, Midori_rounds_sub_ResultXORkey[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U107 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6244, new_AGEMA_signal_6241}), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, Midori_rounds_sub_ResultXORkey[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U105 ( .a ({new_AGEMA_signal_6256, new_AGEMA_signal_6253, new_AGEMA_signal_6250}), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, Midori_rounds_sub_ResultXORkey[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U102 ( .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6262, new_AGEMA_signal_6259}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, Midori_rounds_sub_ResultXORkey[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U100 ( .a ({new_AGEMA_signal_6274, new_AGEMA_signal_6271, new_AGEMA_signal_6268}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_sub_ResultXORkey[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U98 ( .a ({new_AGEMA_signal_6283, new_AGEMA_signal_6280, new_AGEMA_signal_6277}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, Midori_rounds_sub_ResultXORkey[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U96 ( .a ({new_AGEMA_signal_6292, new_AGEMA_signal_6289, new_AGEMA_signal_6286}), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_sub_ResultXORkey[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U94 ( .a ({new_AGEMA_signal_6301, new_AGEMA_signal_6298, new_AGEMA_signal_6295}), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, Midori_rounds_sub_ResultXORkey[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U92 ( .a ({new_AGEMA_signal_6310, new_AGEMA_signal_6307, new_AGEMA_signal_6304}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_sub_ResultXORkey[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U91 ( .a ({new_AGEMA_signal_6319, new_AGEMA_signal_6316, new_AGEMA_signal_6313}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, Midori_rounds_sub_ResultXORkey[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U89 ( .a ({new_AGEMA_signal_6328, new_AGEMA_signal_6325, new_AGEMA_signal_6322}), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_sub_ResultXORkey[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U87 ( .a ({new_AGEMA_signal_6337, new_AGEMA_signal_6334, new_AGEMA_signal_6331}), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, Midori_rounds_sub_ResultXORkey[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U85 ( .a ({new_AGEMA_signal_6346, new_AGEMA_signal_6343, new_AGEMA_signal_6340}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_sub_ResultXORkey[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U83 ( .a ({new_AGEMA_signal_6355, new_AGEMA_signal_6352, new_AGEMA_signal_6349}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, Midori_rounds_sub_ResultXORkey[11]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U80 ( .a ({new_AGEMA_signal_6076, new_AGEMA_signal_6073, new_AGEMA_signal_6070}), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_mul_ResultXORkey[9]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U77 ( .a ({new_AGEMA_signal_6085, new_AGEMA_signal_6082, new_AGEMA_signal_6079}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, Midori_rounds_mul_ResultXORkey[7]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U75 ( .a ({new_AGEMA_signal_6094, new_AGEMA_signal_6091, new_AGEMA_signal_6088}), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, Midori_rounds_mul_ResultXORkey[63]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U73 ( .a ({new_AGEMA_signal_6103, new_AGEMA_signal_6100, new_AGEMA_signal_6097}), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_mul_ResultXORkey[61]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U70 ( .a ({new_AGEMA_signal_6112, new_AGEMA_signal_6109, new_AGEMA_signal_6106}), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, Midori_rounds_mul_ResultXORkey[5]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U69 ( .a ({new_AGEMA_signal_6121, new_AGEMA_signal_6118, new_AGEMA_signal_6115}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, Midori_rounds_mul_ResultXORkey[59]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U67 ( .a ({new_AGEMA_signal_6130, new_AGEMA_signal_6127, new_AGEMA_signal_6124}), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, Midori_rounds_mul_ResultXORkey[57]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U64 ( .a ({new_AGEMA_signal_6139, new_AGEMA_signal_6136, new_AGEMA_signal_6133}), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, Midori_rounds_mul_ResultXORkey[55]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U62 ( .a ({new_AGEMA_signal_6148, new_AGEMA_signal_6145, new_AGEMA_signal_6142}), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, Midori_rounds_mul_ResultXORkey[53]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U59 ( .a ({new_AGEMA_signal_6157, new_AGEMA_signal_6154, new_AGEMA_signal_6151}), .b ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, Midori_rounds_mul_ResultXORkey[51]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U55 ( .a ({new_AGEMA_signal_6166, new_AGEMA_signal_6163, new_AGEMA_signal_6160}), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, Midori_rounds_mul_ResultXORkey[49]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U52 ( .a ({new_AGEMA_signal_6175, new_AGEMA_signal_6172, new_AGEMA_signal_6169}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, Midori_rounds_mul_ResultXORkey[47]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U50 ( .a ({new_AGEMA_signal_6184, new_AGEMA_signal_6181, new_AGEMA_signal_6178}), .b ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, Midori_rounds_mul_ResultXORkey[45]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U47 ( .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6190, new_AGEMA_signal_6187}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_mul_ResultXORkey[43]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U45 ( .a ({new_AGEMA_signal_6202, new_AGEMA_signal_6199, new_AGEMA_signal_6196}), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, Midori_rounds_mul_ResultXORkey[41]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U42 ( .a ({new_AGEMA_signal_6211, new_AGEMA_signal_6208, new_AGEMA_signal_6205}), .b ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_mul_ResultXORkey[3]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U41 ( .a ({new_AGEMA_signal_6220, new_AGEMA_signal_6217, new_AGEMA_signal_6214}), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, Midori_rounds_mul_ResultXORkey[39]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U39 ( .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6226, new_AGEMA_signal_6223}), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_mul_ResultXORkey[37]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U36 ( .a ({new_AGEMA_signal_6238, new_AGEMA_signal_6235, new_AGEMA_signal_6232}), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, Midori_rounds_mul_ResultXORkey[35]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U34 ( .a ({new_AGEMA_signal_6247, new_AGEMA_signal_6244, new_AGEMA_signal_6241}), .b ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, Midori_rounds_mul_ResultXORkey[33]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U31 ( .a ({new_AGEMA_signal_6256, new_AGEMA_signal_6253, new_AGEMA_signal_6250}), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, Midori_rounds_mul_ResultXORkey[31]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U28 ( .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6262, new_AGEMA_signal_6259}), .b ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, Midori_rounds_mul_ResultXORkey[29]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U25 ( .a ({new_AGEMA_signal_6274, new_AGEMA_signal_6271, new_AGEMA_signal_6268}), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_mul_ResultXORkey[27]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U23 ( .a ({new_AGEMA_signal_6283, new_AGEMA_signal_6280, new_AGEMA_signal_6277}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, Midori_rounds_mul_ResultXORkey[25]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U20 ( .a ({new_AGEMA_signal_6292, new_AGEMA_signal_6289, new_AGEMA_signal_6286}), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_mul_ResultXORkey[23]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U18 ( .a ({new_AGEMA_signal_6301, new_AGEMA_signal_6298, new_AGEMA_signal_6295}), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, Midori_rounds_mul_ResultXORkey[21]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U15 ( .a ({new_AGEMA_signal_6310, new_AGEMA_signal_6307, new_AGEMA_signal_6304}), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, Midori_rounds_mul_ResultXORkey[1]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U14 ( .a ({new_AGEMA_signal_6319, new_AGEMA_signal_6316, new_AGEMA_signal_6313}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, Midori_rounds_mul_ResultXORkey[19]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U12 ( .a ({new_AGEMA_signal_6328, new_AGEMA_signal_6325, new_AGEMA_signal_6322}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, Midori_rounds_mul_ResultXORkey[17]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U9 ( .a ({new_AGEMA_signal_6337, new_AGEMA_signal_6334, new_AGEMA_signal_6331}), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, Midori_rounds_mul_ResultXORkey[15]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U7 ( .a ({new_AGEMA_signal_6346, new_AGEMA_signal_6343, new_AGEMA_signal_6340}), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, Midori_rounds_mul_ResultXORkey[13]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U4 ( .a ({new_AGEMA_signal_6355, new_AGEMA_signal_6352, new_AGEMA_signal_6349}), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, Midori_rounds_mul_ResultXORkey[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_round_Result[1]}), .a ({new_AGEMA_signal_6367, new_AGEMA_signal_6364, new_AGEMA_signal_6361}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, Midori_rounds_roundResult_Reg_SFF_1_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, Midori_rounds_round_Result[3]}), .a ({new_AGEMA_signal_6376, new_AGEMA_signal_6373, new_AGEMA_signal_6370}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, Midori_rounds_roundResult_Reg_SFF_3_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_round_Result[5]}), .a ({new_AGEMA_signal_6385, new_AGEMA_signal_6382, new_AGEMA_signal_6379}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, Midori_rounds_roundResult_Reg_SFF_5_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, Midori_rounds_round_Result[7]}), .a ({new_AGEMA_signal_6394, new_AGEMA_signal_6391, new_AGEMA_signal_6388}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, Midori_rounds_roundResult_Reg_SFF_7_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_round_Result[9]}), .a ({new_AGEMA_signal_6403, new_AGEMA_signal_6400, new_AGEMA_signal_6397}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, Midori_rounds_roundResult_Reg_SFF_9_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, Midori_rounds_round_Result[11]}), .a ({new_AGEMA_signal_6412, new_AGEMA_signal_6409, new_AGEMA_signal_6406}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, Midori_rounds_roundResult_Reg_SFF_11_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_round_Result[13]}), .a ({new_AGEMA_signal_6421, new_AGEMA_signal_6418, new_AGEMA_signal_6415}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, Midori_rounds_roundResult_Reg_SFF_13_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, Midori_rounds_round_Result[15]}), .a ({new_AGEMA_signal_6430, new_AGEMA_signal_6427, new_AGEMA_signal_6424}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, Midori_rounds_roundResult_Reg_SFF_15_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_round_Result[17]}), .a ({new_AGEMA_signal_6439, new_AGEMA_signal_6436, new_AGEMA_signal_6433}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, Midori_rounds_roundResult_Reg_SFF_17_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, Midori_rounds_round_Result[19]}), .a ({new_AGEMA_signal_6448, new_AGEMA_signal_6445, new_AGEMA_signal_6442}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, Midori_rounds_roundResult_Reg_SFF_19_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_round_Result[21]}), .a ({new_AGEMA_signal_6457, new_AGEMA_signal_6454, new_AGEMA_signal_6451}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, Midori_rounds_roundResult_Reg_SFF_21_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, Midori_rounds_round_Result[23]}), .a ({new_AGEMA_signal_6466, new_AGEMA_signal_6463, new_AGEMA_signal_6460}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, Midori_rounds_roundResult_Reg_SFF_23_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_round_Result[25]}), .a ({new_AGEMA_signal_6475, new_AGEMA_signal_6472, new_AGEMA_signal_6469}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, Midori_rounds_roundResult_Reg_SFF_25_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, Midori_rounds_round_Result[27]}), .a ({new_AGEMA_signal_6484, new_AGEMA_signal_6481, new_AGEMA_signal_6478}), .c ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, Midori_rounds_roundResult_Reg_SFF_27_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_round_Result[29]}), .a ({new_AGEMA_signal_6493, new_AGEMA_signal_6490, new_AGEMA_signal_6487}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, Midori_rounds_roundResult_Reg_SFF_29_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, Midori_rounds_round_Result[31]}), .a ({new_AGEMA_signal_6502, new_AGEMA_signal_6499, new_AGEMA_signal_6496}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, Midori_rounds_roundResult_Reg_SFF_31_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_round_Result[33]}), .a ({new_AGEMA_signal_6511, new_AGEMA_signal_6508, new_AGEMA_signal_6505}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, Midori_rounds_roundResult_Reg_SFF_33_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, Midori_rounds_round_Result[35]}), .a ({new_AGEMA_signal_6520, new_AGEMA_signal_6517, new_AGEMA_signal_6514}), .c ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, Midori_rounds_roundResult_Reg_SFF_35_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_round_Result[37]}), .a ({new_AGEMA_signal_6529, new_AGEMA_signal_6526, new_AGEMA_signal_6523}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, Midori_rounds_roundResult_Reg_SFF_37_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, Midori_rounds_round_Result[39]}), .a ({new_AGEMA_signal_6538, new_AGEMA_signal_6535, new_AGEMA_signal_6532}), .c ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, Midori_rounds_roundResult_Reg_SFF_39_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_round_Result[41]}), .a ({new_AGEMA_signal_6547, new_AGEMA_signal_6544, new_AGEMA_signal_6541}), .c ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, Midori_rounds_roundResult_Reg_SFF_41_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, Midori_rounds_round_Result[43]}), .a ({new_AGEMA_signal_6556, new_AGEMA_signal_6553, new_AGEMA_signal_6550}), .c ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, Midori_rounds_roundResult_Reg_SFF_43_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_round_Result[45]}), .a ({new_AGEMA_signal_6565, new_AGEMA_signal_6562, new_AGEMA_signal_6559}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, Midori_rounds_roundResult_Reg_SFF_45_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, Midori_rounds_round_Result[47]}), .a ({new_AGEMA_signal_6574, new_AGEMA_signal_6571, new_AGEMA_signal_6568}), .c ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, Midori_rounds_roundResult_Reg_SFF_47_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_round_Result[49]}), .a ({new_AGEMA_signal_6583, new_AGEMA_signal_6580, new_AGEMA_signal_6577}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, Midori_rounds_roundResult_Reg_SFF_49_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, Midori_rounds_round_Result[51]}), .a ({new_AGEMA_signal_6592, new_AGEMA_signal_6589, new_AGEMA_signal_6586}), .c ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, Midori_rounds_roundResult_Reg_SFF_51_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_round_Result[53]}), .a ({new_AGEMA_signal_6601, new_AGEMA_signal_6598, new_AGEMA_signal_6595}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, Midori_rounds_roundResult_Reg_SFF_53_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, Midori_rounds_round_Result[55]}), .a ({new_AGEMA_signal_6610, new_AGEMA_signal_6607, new_AGEMA_signal_6604}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, Midori_rounds_roundResult_Reg_SFF_55_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_round_Result[57]}), .a ({new_AGEMA_signal_6619, new_AGEMA_signal_6616, new_AGEMA_signal_6613}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Midori_rounds_roundResult_Reg_SFF_57_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, Midori_rounds_round_Result[59]}), .a ({new_AGEMA_signal_6628, new_AGEMA_signal_6625, new_AGEMA_signal_6622}), .c ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Midori_rounds_roundResult_Reg_SFF_59_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_round_Result[61]}), .a ({new_AGEMA_signal_6637, new_AGEMA_signal_6634, new_AGEMA_signal_6631}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Midori_rounds_roundResult_Reg_SFF_61_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1 ( .s (new_AGEMA_signal_6358), .b ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, Midori_rounds_round_Result[63]}), .a ({new_AGEMA_signal_6646, new_AGEMA_signal_6643, new_AGEMA_signal_6640}), .c ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Midori_rounds_roundResult_Reg_SFF_63_DQ}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .a ({new_AGEMA_signal_6649, new_AGEMA_signal_6648, new_AGEMA_signal_6647}), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, Midori_rounds_sub_sBox_PRINCE_0_n14}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .a ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, Midori_rounds_sub_sBox_PRINCE_0_n11}), .b ({new_AGEMA_signal_6652, new_AGEMA_signal_6651, new_AGEMA_signal_6650}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, Midori_rounds_sub_sBox_PRINCE_0_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .a ({new_AGEMA_signal_6655, new_AGEMA_signal_6654, new_AGEMA_signal_6653}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2678, Midori_rounds_sub_sBox_PRINCE_0_n5}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .a ({new_AGEMA_signal_6652, new_AGEMA_signal_6651, new_AGEMA_signal_6650}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, Midori_rounds_sub_sBox_PRINCE_0_n2}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_rounds_sub_sBox_PRINCE_0_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .a ({new_AGEMA_signal_6658, new_AGEMA_signal_6657, new_AGEMA_signal_6656}), .b ({new_AGEMA_signal_2685, new_AGEMA_signal_2684, Midori_rounds_sub_sBox_PRINCE_1_n14}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .a ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, Midori_rounds_sub_sBox_PRINCE_1_n11}), .b ({new_AGEMA_signal_6661, new_AGEMA_signal_6660, new_AGEMA_signal_6659}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_rounds_sub_sBox_PRINCE_1_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .a ({new_AGEMA_signal_6664, new_AGEMA_signal_6663, new_AGEMA_signal_6662}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, Midori_rounds_sub_sBox_PRINCE_1_n5}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .a ({new_AGEMA_signal_6661, new_AGEMA_signal_6660, new_AGEMA_signal_6659}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, Midori_rounds_sub_sBox_PRINCE_1_n2}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, Midori_rounds_sub_sBox_PRINCE_1_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .a ({new_AGEMA_signal_6667, new_AGEMA_signal_6666, new_AGEMA_signal_6665}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, Midori_rounds_sub_sBox_PRINCE_2_n14}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .a ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, Midori_rounds_sub_sBox_PRINCE_2_n11}), .b ({new_AGEMA_signal_6670, new_AGEMA_signal_6669, new_AGEMA_signal_6668}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, Midori_rounds_sub_sBox_PRINCE_2_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .a ({new_AGEMA_signal_6673, new_AGEMA_signal_6672, new_AGEMA_signal_6671}), .b ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, Midori_rounds_sub_sBox_PRINCE_2_n5}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .a ({new_AGEMA_signal_6670, new_AGEMA_signal_6669, new_AGEMA_signal_6668}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, Midori_rounds_sub_sBox_PRINCE_2_n2}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, Midori_rounds_sub_sBox_PRINCE_2_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .a ({new_AGEMA_signal_6676, new_AGEMA_signal_6675, new_AGEMA_signal_6674}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, Midori_rounds_sub_sBox_PRINCE_3_n14}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .a ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, Midori_rounds_sub_sBox_PRINCE_3_n11}), .b ({new_AGEMA_signal_6679, new_AGEMA_signal_6678, new_AGEMA_signal_6677}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, Midori_rounds_sub_sBox_PRINCE_3_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .a ({new_AGEMA_signal_6682, new_AGEMA_signal_6681, new_AGEMA_signal_6680}), .b ({new_AGEMA_signal_2709, new_AGEMA_signal_2708, Midori_rounds_sub_sBox_PRINCE_3_n5}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .a ({new_AGEMA_signal_6679, new_AGEMA_signal_6678, new_AGEMA_signal_6677}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, Midori_rounds_sub_sBox_PRINCE_3_n2}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_rounds_sub_sBox_PRINCE_3_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .a ({new_AGEMA_signal_6685, new_AGEMA_signal_6684, new_AGEMA_signal_6683}), .b ({new_AGEMA_signal_2715, new_AGEMA_signal_2714, Midori_rounds_sub_sBox_PRINCE_4_n14}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .a ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, Midori_rounds_sub_sBox_PRINCE_4_n11}), .b ({new_AGEMA_signal_6688, new_AGEMA_signal_6687, new_AGEMA_signal_6686}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_rounds_sub_sBox_PRINCE_4_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .a ({new_AGEMA_signal_6691, new_AGEMA_signal_6690, new_AGEMA_signal_6689}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, Midori_rounds_sub_sBox_PRINCE_4_n5}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .a ({new_AGEMA_signal_6688, new_AGEMA_signal_6687, new_AGEMA_signal_6686}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, Midori_rounds_sub_sBox_PRINCE_4_n2}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, Midori_rounds_sub_sBox_PRINCE_4_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .a ({new_AGEMA_signal_6694, new_AGEMA_signal_6693, new_AGEMA_signal_6692}), .b ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, Midori_rounds_sub_sBox_PRINCE_5_n14}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .a ({new_AGEMA_signal_2439, new_AGEMA_signal_2438, Midori_rounds_sub_sBox_PRINCE_5_n11}), .b ({new_AGEMA_signal_6697, new_AGEMA_signal_6696, new_AGEMA_signal_6695}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, Midori_rounds_sub_sBox_PRINCE_5_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .a ({new_AGEMA_signal_6700, new_AGEMA_signal_6699, new_AGEMA_signal_6698}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, Midori_rounds_sub_sBox_PRINCE_5_n5}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .a ({new_AGEMA_signal_6697, new_AGEMA_signal_6696, new_AGEMA_signal_6695}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, Midori_rounds_sub_sBox_PRINCE_5_n2}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, Midori_rounds_sub_sBox_PRINCE_5_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .a ({new_AGEMA_signal_6703, new_AGEMA_signal_6702, new_AGEMA_signal_6701}), .b ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, Midori_rounds_sub_sBox_PRINCE_6_n14}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .a ({new_AGEMA_signal_2451, new_AGEMA_signal_2450, Midori_rounds_sub_sBox_PRINCE_6_n11}), .b ({new_AGEMA_signal_6706, new_AGEMA_signal_6705, new_AGEMA_signal_6704}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, Midori_rounds_sub_sBox_PRINCE_6_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .a ({new_AGEMA_signal_6709, new_AGEMA_signal_6708, new_AGEMA_signal_6707}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, Midori_rounds_sub_sBox_PRINCE_6_n5}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .a ({new_AGEMA_signal_6706, new_AGEMA_signal_6705, new_AGEMA_signal_6704}), .b ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, Midori_rounds_sub_sBox_PRINCE_6_n2}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_rounds_sub_sBox_PRINCE_6_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .a ({new_AGEMA_signal_6712, new_AGEMA_signal_6711, new_AGEMA_signal_6710}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, Midori_rounds_sub_sBox_PRINCE_7_n14}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .a ({new_AGEMA_signal_2463, new_AGEMA_signal_2462, Midori_rounds_sub_sBox_PRINCE_7_n11}), .b ({new_AGEMA_signal_6715, new_AGEMA_signal_6714, new_AGEMA_signal_6713}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_rounds_sub_sBox_PRINCE_7_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .a ({new_AGEMA_signal_6718, new_AGEMA_signal_6717, new_AGEMA_signal_6716}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, Midori_rounds_sub_sBox_PRINCE_7_n5}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .a ({new_AGEMA_signal_6715, new_AGEMA_signal_6714, new_AGEMA_signal_6713}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, Midori_rounds_sub_sBox_PRINCE_7_n2}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, Midori_rounds_sub_sBox_PRINCE_7_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .a ({new_AGEMA_signal_6721, new_AGEMA_signal_6720, new_AGEMA_signal_6719}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, Midori_rounds_sub_sBox_PRINCE_8_n14}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .a ({new_AGEMA_signal_2475, new_AGEMA_signal_2474, Midori_rounds_sub_sBox_PRINCE_8_n11}), .b ({new_AGEMA_signal_6724, new_AGEMA_signal_6723, new_AGEMA_signal_6722}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, Midori_rounds_sub_sBox_PRINCE_8_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .a ({new_AGEMA_signal_6727, new_AGEMA_signal_6726, new_AGEMA_signal_6725}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, Midori_rounds_sub_sBox_PRINCE_8_n5}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .a ({new_AGEMA_signal_6724, new_AGEMA_signal_6723, new_AGEMA_signal_6722}), .b ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, Midori_rounds_sub_sBox_PRINCE_8_n2}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, Midori_rounds_sub_sBox_PRINCE_8_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .a ({new_AGEMA_signal_6730, new_AGEMA_signal_6729, new_AGEMA_signal_6728}), .b ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, Midori_rounds_sub_sBox_PRINCE_9_n14}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .a ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, Midori_rounds_sub_sBox_PRINCE_9_n11}), .b ({new_AGEMA_signal_6733, new_AGEMA_signal_6732, new_AGEMA_signal_6731}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, Midori_rounds_sub_sBox_PRINCE_9_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .a ({new_AGEMA_signal_6736, new_AGEMA_signal_6735, new_AGEMA_signal_6734}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, Midori_rounds_sub_sBox_PRINCE_9_n5}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .a ({new_AGEMA_signal_6733, new_AGEMA_signal_6732, new_AGEMA_signal_6731}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, Midori_rounds_sub_sBox_PRINCE_9_n2}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_rounds_sub_sBox_PRINCE_9_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .a ({new_AGEMA_signal_6739, new_AGEMA_signal_6738, new_AGEMA_signal_6737}), .b ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, Midori_rounds_sub_sBox_PRINCE_10_n14}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .a ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, Midori_rounds_sub_sBox_PRINCE_10_n11}), .b ({new_AGEMA_signal_6742, new_AGEMA_signal_6741, new_AGEMA_signal_6740}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_rounds_sub_sBox_PRINCE_10_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .a ({new_AGEMA_signal_6745, new_AGEMA_signal_6744, new_AGEMA_signal_6743}), .b ({new_AGEMA_signal_2779, new_AGEMA_signal_2778, Midori_rounds_sub_sBox_PRINCE_10_n5}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .a ({new_AGEMA_signal_6742, new_AGEMA_signal_6741, new_AGEMA_signal_6740}), .b ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, Midori_rounds_sub_sBox_PRINCE_10_n2}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, Midori_rounds_sub_sBox_PRINCE_10_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .a ({new_AGEMA_signal_6748, new_AGEMA_signal_6747, new_AGEMA_signal_6746}), .b ({new_AGEMA_signal_2785, new_AGEMA_signal_2784, Midori_rounds_sub_sBox_PRINCE_11_n14}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .a ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, Midori_rounds_sub_sBox_PRINCE_11_n11}), .b ({new_AGEMA_signal_6751, new_AGEMA_signal_6750, new_AGEMA_signal_6749}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, Midori_rounds_sub_sBox_PRINCE_11_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .a ({new_AGEMA_signal_6754, new_AGEMA_signal_6753, new_AGEMA_signal_6752}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, Midori_rounds_sub_sBox_PRINCE_11_n5}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .a ({new_AGEMA_signal_6751, new_AGEMA_signal_6750, new_AGEMA_signal_6749}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, Midori_rounds_sub_sBox_PRINCE_11_n2}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, Midori_rounds_sub_sBox_PRINCE_11_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .a ({new_AGEMA_signal_6757, new_AGEMA_signal_6756, new_AGEMA_signal_6755}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, Midori_rounds_sub_sBox_PRINCE_12_n14}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .a ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, Midori_rounds_sub_sBox_PRINCE_12_n11}), .b ({new_AGEMA_signal_6760, new_AGEMA_signal_6759, new_AGEMA_signal_6758}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, Midori_rounds_sub_sBox_PRINCE_12_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .a ({new_AGEMA_signal_6763, new_AGEMA_signal_6762, new_AGEMA_signal_6761}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, Midori_rounds_sub_sBox_PRINCE_12_n5}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .a ({new_AGEMA_signal_6760, new_AGEMA_signal_6759, new_AGEMA_signal_6758}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, Midori_rounds_sub_sBox_PRINCE_12_n2}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_rounds_sub_sBox_PRINCE_12_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .a ({new_AGEMA_signal_6766, new_AGEMA_signal_6765, new_AGEMA_signal_6764}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, Midori_rounds_sub_sBox_PRINCE_13_n14}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .a ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, Midori_rounds_sub_sBox_PRINCE_13_n11}), .b ({new_AGEMA_signal_6769, new_AGEMA_signal_6768, new_AGEMA_signal_6767}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_rounds_sub_sBox_PRINCE_13_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .a ({new_AGEMA_signal_6772, new_AGEMA_signal_6771, new_AGEMA_signal_6770}), .b ({new_AGEMA_signal_2809, new_AGEMA_signal_2808, Midori_rounds_sub_sBox_PRINCE_13_n5}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .a ({new_AGEMA_signal_6769, new_AGEMA_signal_6768, new_AGEMA_signal_6767}), .b ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, Midori_rounds_sub_sBox_PRINCE_13_n2}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, Midori_rounds_sub_sBox_PRINCE_13_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .a ({new_AGEMA_signal_6775, new_AGEMA_signal_6774, new_AGEMA_signal_6773}), .b ({new_AGEMA_signal_2815, new_AGEMA_signal_2814, Midori_rounds_sub_sBox_PRINCE_14_n14}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .a ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, Midori_rounds_sub_sBox_PRINCE_14_n11}), .b ({new_AGEMA_signal_6778, new_AGEMA_signal_6777, new_AGEMA_signal_6776}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, Midori_rounds_sub_sBox_PRINCE_14_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .a ({new_AGEMA_signal_6781, new_AGEMA_signal_6780, new_AGEMA_signal_6779}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, Midori_rounds_sub_sBox_PRINCE_14_n5}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .a ({new_AGEMA_signal_6778, new_AGEMA_signal_6777, new_AGEMA_signal_6776}), .b ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, Midori_rounds_sub_sBox_PRINCE_14_n2}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, Midori_rounds_sub_sBox_PRINCE_14_n3}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .a ({new_AGEMA_signal_6784, new_AGEMA_signal_6783, new_AGEMA_signal_6782}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, Midori_rounds_sub_sBox_PRINCE_15_n14}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .a ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, Midori_rounds_sub_sBox_PRINCE_15_n11}), .b ({new_AGEMA_signal_6787, new_AGEMA_signal_6786, new_AGEMA_signal_6785}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, Midori_rounds_sub_sBox_PRINCE_15_n12}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .a ({new_AGEMA_signal_6790, new_AGEMA_signal_6789, new_AGEMA_signal_6788}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, Midori_rounds_sub_sBox_PRINCE_15_n5}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .a ({new_AGEMA_signal_6787, new_AGEMA_signal_6786, new_AGEMA_signal_6785}), .b ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, Midori_rounds_sub_sBox_PRINCE_15_n2}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_rounds_sub_sBox_PRINCE_15_n3}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_1_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, Midori_rounds_SR_Result[1]}), .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, Midori_rounds_sub_ResultXORkey[1]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_3_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2889, new_AGEMA_signal_2888, Midori_rounds_SR_Result[3]}), .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, Midori_rounds_sub_ResultXORkey[3]}), .c ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_5_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, Midori_rounds_SR_Result[5]}), .a ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, Midori_rounds_sub_ResultXORkey[5]}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_7_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, Midori_rounds_SR_Result[7]}), .a ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, Midori_rounds_sub_ResultXORkey[7]}), .c ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_9_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, Midori_rounds_SR_Result[9]}), .a ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, Midori_rounds_sub_ResultXORkey[9]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_11_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, Midori_rounds_SR_Result[11]}), .a ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, Midori_rounds_sub_ResultXORkey[11]}), .c ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_13_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2901, new_AGEMA_signal_2900, Midori_rounds_SR_Result[13]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, Midori_rounds_sub_ResultXORkey[13]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_15_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, Midori_rounds_SR_Result[15]}), .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, Midori_rounds_sub_ResultXORkey[15]}), .c ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_17_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, Midori_rounds_SR_Result[17]}), .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, Midori_rounds_sub_ResultXORkey[17]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_19_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, Midori_rounds_SR_Result[19]}), .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, Midori_rounds_sub_ResultXORkey[19]}), .c ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_21_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, Midori_rounds_SR_Result[21]}), .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, Midori_rounds_sub_ResultXORkey[21]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_23_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2857, new_AGEMA_signal_2856, Midori_rounds_SR_Result[23]}), .a ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, Midori_rounds_sub_ResultXORkey[23]}), .c ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_25_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, Midori_rounds_SR_Result[25]}), .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, Midori_rounds_sub_ResultXORkey[25]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_27_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, Midori_rounds_SR_Result[27]}), .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, Midori_rounds_sub_ResultXORkey[27]}), .c ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_29_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, Midori_rounds_SR_Result[29]}), .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, Midori_rounds_sub_ResultXORkey[29]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_31_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, Midori_rounds_SR_Result[31]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, Midori_rounds_sub_ResultXORkey[31]}), .c ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_33_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, Midori_rounds_SR_Result[33]}), .a ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, Midori_rounds_sub_ResultXORkey[33]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_35_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, Midori_rounds_SR_Result[35]}), .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, Midori_rounds_sub_ResultXORkey[35]}), .c ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_37_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2869, new_AGEMA_signal_2868, Midori_rounds_SR_Result[37]}), .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, Midori_rounds_sub_ResultXORkey[37]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_39_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, Midori_rounds_SR_Result[39]}), .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, Midori_rounds_sub_ResultXORkey[39]}), .c ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_41_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, Midori_rounds_SR_Result[41]}), .a ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, Midori_rounds_sub_ResultXORkey[41]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_43_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, Midori_rounds_SR_Result[43]}), .a ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, Midori_rounds_sub_ResultXORkey[43]}), .c ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_45_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2845, new_AGEMA_signal_2844, Midori_rounds_SR_Result[45]}), .a ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, Midori_rounds_sub_ResultXORkey[45]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_47_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, Midori_rounds_SR_Result[47]}), .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, Midori_rounds_sub_ResultXORkey[47]}), .c ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_49_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, Midori_rounds_SR_Result[49]}), .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, Midori_rounds_sub_ResultXORkey[49]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_51_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2833, new_AGEMA_signal_2832, Midori_rounds_SR_Result[51]}), .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, Midori_rounds_sub_ResultXORkey[51]}), .c ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_53_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, Midori_rounds_SR_Result[53]}), .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, Midori_rounds_sub_ResultXORkey[53]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_55_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2913, new_AGEMA_signal_2912, Midori_rounds_SR_Result[55]}), .a ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, Midori_rounds_sub_ResultXORkey[55]}), .c ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_57_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2877, new_AGEMA_signal_2876, Midori_rounds_SR_Result[57]}), .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, Midori_rounds_sub_ResultXORkey[57]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_59_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, Midori_rounds_SR_Result[59]}), .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, Midori_rounds_sub_ResultXORkey[59]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_61_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, Midori_rounds_SR_Result[61]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, Midori_rounds_sub_ResultXORkey[61]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_63_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, Midori_rounds_SR_Result[63]}), .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, Midori_rounds_sub_ResultXORkey[63]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U24 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U22 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U20 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U18 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U17 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, Midori_rounds_mul_MC1_n6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U14 ( .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U13 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, Midori_rounds_mul_input[61]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, Midori_rounds_mul_MC1_n4}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U12 ( .a ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, Midori_rounds_mul_input[59]}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U10 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U9 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, Midori_rounds_mul_input[53]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, Midori_rounds_mul_MC1_n8}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U6 ( .a ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U5 ( .a ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, Midori_rounds_mul_input[55]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, Midori_rounds_mul_MC1_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U24 ( .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U22 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U20 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U18 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U17 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, Midori_rounds_mul_MC2_n6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U14 ( .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U13 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, Midori_rounds_mul_input[45]}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, Midori_rounds_mul_MC2_n4}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U12 ( .a ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, Midori_rounds_mul_input[43]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U10 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U9 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, Midori_rounds_mul_input[37]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, Midori_rounds_mul_MC2_n8}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U6 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U5 ( .a ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, Midori_rounds_mul_input[39]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, Midori_rounds_mul_MC2_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U24 ( .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U22 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U20 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U18 ( .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U17 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, Midori_rounds_mul_MC3_n6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U14 ( .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U13 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, Midori_rounds_mul_input[29]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, Midori_rounds_mul_MC3_n4}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U12 ( .a ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, Midori_rounds_mul_input[27]}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U10 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U9 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, Midori_rounds_mul_input[21]}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, Midori_rounds_mul_MC3_n8}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U6 ( .a ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U5 ( .a ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, Midori_rounds_mul_input[23]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, Midori_rounds_mul_MC3_n2}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U24 ( .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U22 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U20 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U18 ( .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U17 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, Midori_rounds_mul_MC4_n6}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U14 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U13 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, Midori_rounds_mul_input[13]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, Midori_rounds_mul_MC4_n4}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U12 ( .a ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, Midori_rounds_mul_input[11]}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U10 ( .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U9 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, Midori_rounds_mul_input[5]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, Midori_rounds_mul_MC4_n8}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U6 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U5 ( .a ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, Midori_rounds_mul_input[7]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, Midori_rounds_mul_MC4_n2}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_1_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, Midori_rounds_mul_ResultXORkey[1]}), .a ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, Midori_rounds_round_Result[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_3_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, Midori_rounds_mul_ResultXORkey[3]}), .a ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, Midori_rounds_round_Result[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_5_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, Midori_rounds_mul_ResultXORkey[5]}), .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, Midori_rounds_round_Result[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_7_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, Midori_rounds_mul_ResultXORkey[7]}), .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, Midori_rounds_round_Result[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_9_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, Midori_rounds_mul_ResultXORkey[9]}), .a ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, Midori_rounds_round_Result[9]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_11_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, Midori_rounds_mul_ResultXORkey[11]}), .a ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, Midori_rounds_round_Result[11]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_13_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, Midori_rounds_mul_ResultXORkey[13]}), .a ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, Midori_rounds_round_Result[13]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_15_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, Midori_rounds_mul_ResultXORkey[15]}), .a ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, Midori_rounds_round_Result[15]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_17_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, Midori_rounds_mul_ResultXORkey[17]}), .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, Midori_rounds_round_Result[17]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_19_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, Midori_rounds_mul_ResultXORkey[19]}), .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, Midori_rounds_round_Result[19]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_21_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, Midori_rounds_mul_ResultXORkey[21]}), .a ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, Midori_rounds_round_Result[21]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_23_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, Midori_rounds_mul_ResultXORkey[23]}), .a ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, Midori_rounds_round_Result[23]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_25_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, Midori_rounds_mul_ResultXORkey[25]}), .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, Midori_rounds_round_Result[25]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_27_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, Midori_rounds_mul_ResultXORkey[27]}), .a ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, Midori_rounds_round_Result[27]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_29_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, Midori_rounds_mul_ResultXORkey[29]}), .a ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, Midori_rounds_round_Result[29]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_31_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, Midori_rounds_mul_ResultXORkey[31]}), .a ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, Midori_rounds_round_Result[31]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_33_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, Midori_rounds_mul_ResultXORkey[33]}), .a ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, Midori_rounds_round_Result[33]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_35_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, Midori_rounds_mul_ResultXORkey[35]}), .a ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, Midori_rounds_round_Result[35]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_37_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, Midori_rounds_mul_ResultXORkey[37]}), .a ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, Midori_rounds_round_Result[37]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_39_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, Midori_rounds_mul_ResultXORkey[39]}), .a ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, Midori_rounds_round_Result[39]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_41_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, Midori_rounds_mul_ResultXORkey[41]}), .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, Midori_rounds_round_Result[41]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_43_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, Midori_rounds_mul_ResultXORkey[43]}), .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, Midori_rounds_round_Result[43]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_45_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, Midori_rounds_mul_ResultXORkey[45]}), .a ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, Midori_rounds_round_Result[45]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_47_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, Midori_rounds_mul_ResultXORkey[47]}), .a ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, Midori_rounds_round_Result[47]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_49_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, Midori_rounds_mul_ResultXORkey[49]}), .a ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, Midori_rounds_round_Result[49]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_51_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, Midori_rounds_mul_ResultXORkey[51]}), .a ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, Midori_rounds_round_Result[51]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_53_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, Midori_rounds_mul_ResultXORkey[53]}), .a ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, Midori_rounds_round_Result[53]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_55_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, Midori_rounds_mul_ResultXORkey[55]}), .a ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, Midori_rounds_round_Result[55]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_57_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, Midori_rounds_mul_ResultXORkey[57]}), .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, Midori_rounds_round_Result[57]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_59_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, Midori_rounds_mul_ResultXORkey[59]}), .a ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, Midori_rounds_round_Result[59]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_61_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, Midori_rounds_mul_ResultXORkey[61]}), .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, Midori_rounds_round_Result[61]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_63_U1 ( .s (new_AGEMA_signal_6793), .b ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, Midori_rounds_mul_ResultXORkey[63]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, Midori_rounds_round_Result[63]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_5781), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_5805), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_5817), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_5829), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_5841), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_5853), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_5865), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_5877), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_5901), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_5925), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_5949), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_5973), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_5997), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_6021), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_6045), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_6057), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_6069), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_6081), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_6093), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_6105), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_6114), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_6117), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_6129), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_6138), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_6141), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_6165), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (new_AGEMA_signal_6189), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (new_AGEMA_signal_6201), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_6210), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (new_AGEMA_signal_6213), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (new_AGEMA_signal_6225), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_6234), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (new_AGEMA_signal_6237), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (new_AGEMA_signal_6249), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_6261), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_6273), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_6285), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_6297), .Q (new_AGEMA_signal_6298) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_6301) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_6304) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_6307) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_6309), .Q (new_AGEMA_signal_6310) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_6319) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_6321), .Q (new_AGEMA_signal_6322) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_6325) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_6331) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_6333), .Q (new_AGEMA_signal_6334) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_6337) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_6340) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_6343) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_6345), .Q (new_AGEMA_signal_6346) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_6349) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_6352) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_6355) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_6357), .Q (new_AGEMA_signal_6358) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_6367) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_6369), .Q (new_AGEMA_signal_6370) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_6373) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_6376) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_6379) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_6381), .Q (new_AGEMA_signal_6382) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_6385) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_6388) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_6391) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_6393), .Q (new_AGEMA_signal_6394) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_6397) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_6403) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_6405), .Q (new_AGEMA_signal_6406) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_6412) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_6415) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_6417), .Q (new_AGEMA_signal_6418) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_6421) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_6424) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_6426), .Q (new_AGEMA_signal_6427) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_6429), .Q (new_AGEMA_signal_6430) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_6433) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_6436) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_6439) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_6441), .Q (new_AGEMA_signal_6442) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_6445) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_6447), .Q (new_AGEMA_signal_6448) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_6450), .Q (new_AGEMA_signal_6451) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_6454) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_6460) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_6463) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_6466) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_6469) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_6471), .Q (new_AGEMA_signal_6472) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_6474), .Q (new_AGEMA_signal_6475) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_6477), .Q (new_AGEMA_signal_6478) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_6481) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_6484) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_6487) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_6489), .Q (new_AGEMA_signal_6490) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_6493) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_6495), .Q (new_AGEMA_signal_6496) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_6498), .Q (new_AGEMA_signal_6499) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_6501), .Q (new_AGEMA_signal_6502) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_6508) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_6511) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_6513), .Q (new_AGEMA_signal_6514) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_6517) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_6519), .Q (new_AGEMA_signal_6520) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_6522), .Q (new_AGEMA_signal_6523) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_6525), .Q (new_AGEMA_signal_6526) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_6529) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_6532) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_6535) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_6537), .Q (new_AGEMA_signal_6538) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_6541) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_6544) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_6546), .Q (new_AGEMA_signal_6547) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_6549), .Q (new_AGEMA_signal_6550) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_6553) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_6555), .Q (new_AGEMA_signal_6556) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_6559) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_6561), .Q (new_AGEMA_signal_6562) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_6564), .Q (new_AGEMA_signal_6565) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_6567), .Q (new_AGEMA_signal_6568) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_6570), .Q (new_AGEMA_signal_6571) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_6573), .Q (new_AGEMA_signal_6574) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_6577) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_6579), .Q (new_AGEMA_signal_6580) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_6582), .Q (new_AGEMA_signal_6583) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_6585), .Q (new_AGEMA_signal_6586) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_6588), .Q (new_AGEMA_signal_6589) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_6591), .Q (new_AGEMA_signal_6592) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_6594), .Q (new_AGEMA_signal_6595) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_6597), .Q (new_AGEMA_signal_6598) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_6600), .Q (new_AGEMA_signal_6601) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_6603), .Q (new_AGEMA_signal_6604) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_6606), .Q (new_AGEMA_signal_6607) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_6609), .Q (new_AGEMA_signal_6610) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_6612), .Q (new_AGEMA_signal_6613) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_6615), .Q (new_AGEMA_signal_6616) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_6618), .Q (new_AGEMA_signal_6619) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_6621), .Q (new_AGEMA_signal_6622) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_6624), .Q (new_AGEMA_signal_6625) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_6627), .Q (new_AGEMA_signal_6628) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_6630), .Q (new_AGEMA_signal_6631) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_6633), .Q (new_AGEMA_signal_6634) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_6636), .Q (new_AGEMA_signal_6637) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_6639), .Q (new_AGEMA_signal_6640) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_6642), .Q (new_AGEMA_signal_6643) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_6645), .Q (new_AGEMA_signal_6646) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_6793) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_6795), .Q (new_AGEMA_signal_6796) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_6799), .Q (new_AGEMA_signal_6800) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_6803), .Q (new_AGEMA_signal_6804) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_6807), .Q (new_AGEMA_signal_6808) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_6811), .Q (new_AGEMA_signal_6812) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_6815), .Q (new_AGEMA_signal_6816) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_6819), .Q (new_AGEMA_signal_6820) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_6823), .Q (new_AGEMA_signal_6824) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_6827), .Q (new_AGEMA_signal_6828) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_6831), .Q (new_AGEMA_signal_6832) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_6835), .Q (new_AGEMA_signal_6836) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_6839), .Q (new_AGEMA_signal_6840) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_6843), .Q (new_AGEMA_signal_6844) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_6847), .Q (new_AGEMA_signal_6848) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_6851), .Q (new_AGEMA_signal_6852) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_6855), .Q (new_AGEMA_signal_6856) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_6859), .Q (new_AGEMA_signal_6860) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_6863), .Q (new_AGEMA_signal_6864) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_6867), .Q (new_AGEMA_signal_6868) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_6871), .Q (new_AGEMA_signal_6872) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_6875), .Q (new_AGEMA_signal_6876) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_6879), .Q (new_AGEMA_signal_6880) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_6883), .Q (new_AGEMA_signal_6884) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_6887), .Q (new_AGEMA_signal_6888) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_6891), .Q (new_AGEMA_signal_6892) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_6895), .Q (new_AGEMA_signal_6896) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_6899), .Q (new_AGEMA_signal_6900) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_6903), .Q (new_AGEMA_signal_6904) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_6907), .Q (new_AGEMA_signal_6908) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_6911), .Q (new_AGEMA_signal_6912) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_6915), .Q (new_AGEMA_signal_6916) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_6919), .Q (new_AGEMA_signal_6920) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_6923), .Q (new_AGEMA_signal_6924) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_6927), .Q (new_AGEMA_signal_6928) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_6931), .Q (new_AGEMA_signal_6932) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_6935), .Q (new_AGEMA_signal_6936) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_6939), .Q (new_AGEMA_signal_6940) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_6943), .Q (new_AGEMA_signal_6944) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_6947), .Q (new_AGEMA_signal_6948) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_6951), .Q (new_AGEMA_signal_6952) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_6955), .Q (new_AGEMA_signal_6956) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_6959), .Q (new_AGEMA_signal_6960) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_6963), .Q (new_AGEMA_signal_6964) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_6967), .Q (new_AGEMA_signal_6968) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_6971), .Q (new_AGEMA_signal_6972) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_6975), .Q (new_AGEMA_signal_6976) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_6979), .Q (new_AGEMA_signal_6980) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_6983), .Q (new_AGEMA_signal_6984) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_6987), .Q (new_AGEMA_signal_6988) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_6991), .Q (new_AGEMA_signal_6992) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_6995), .Q (new_AGEMA_signal_6996) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_6999), .Q (new_AGEMA_signal_7000) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_7003), .Q (new_AGEMA_signal_7004) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_7007), .Q (new_AGEMA_signal_7008) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_7011), .Q (new_AGEMA_signal_7012) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_7015), .Q (new_AGEMA_signal_7016) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_7019), .Q (new_AGEMA_signal_7020) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_7023), .Q (new_AGEMA_signal_7024) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_7027), .Q (new_AGEMA_signal_7028) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_7031), .Q (new_AGEMA_signal_7032) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_7035), .Q (new_AGEMA_signal_7036) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_7039), .Q (new_AGEMA_signal_7040) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_7043), .Q (new_AGEMA_signal_7044) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_7047), .Q (new_AGEMA_signal_7048) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_7051), .Q (new_AGEMA_signal_7052) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_7055), .Q (new_AGEMA_signal_7056) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_7059), .Q (new_AGEMA_signal_7060) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_7063), .Q (new_AGEMA_signal_7064) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_7067), .Q (new_AGEMA_signal_7068) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_7071), .Q (new_AGEMA_signal_7072) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_7075), .Q (new_AGEMA_signal_7076) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_7079), .Q (new_AGEMA_signal_7080) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_7083), .Q (new_AGEMA_signal_7084) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_7087), .Q (new_AGEMA_signal_7088) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_7091), .Q (new_AGEMA_signal_7092) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_7095), .Q (new_AGEMA_signal_7096) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_7099), .Q (new_AGEMA_signal_7100) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_7103), .Q (new_AGEMA_signal_7104) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_7107), .Q (new_AGEMA_signal_7108) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_7111), .Q (new_AGEMA_signal_7112) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_7115), .Q (new_AGEMA_signal_7116) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_7119), .Q (new_AGEMA_signal_7120) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_7123), .Q (new_AGEMA_signal_7124) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_7127), .Q (new_AGEMA_signal_7128) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_7131), .Q (new_AGEMA_signal_7132) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_7135), .Q (new_AGEMA_signal_7136) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_7139), .Q (new_AGEMA_signal_7140) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_7143), .Q (new_AGEMA_signal_7144) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_7148) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_7152) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_7155), .Q (new_AGEMA_signal_7156) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_7159), .Q (new_AGEMA_signal_7160) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_7163), .Q (new_AGEMA_signal_7164) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_7167), .Q (new_AGEMA_signal_7168) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_7171), .Q (new_AGEMA_signal_7172) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_7175), .Q (new_AGEMA_signal_7176) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_7179), .Q (new_AGEMA_signal_7180) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_7184) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_7188) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_7191), .Q (new_AGEMA_signal_7192) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_7195), .Q (new_AGEMA_signal_7196) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_7199), .Q (new_AGEMA_signal_7200) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_7203), .Q (new_AGEMA_signal_7204) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_7207), .Q (new_AGEMA_signal_7208) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_7211), .Q (new_AGEMA_signal_7212) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_7215), .Q (new_AGEMA_signal_7216) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_7219), .Q (new_AGEMA_signal_7220) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_7223), .Q (new_AGEMA_signal_7224) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_7227), .Q (new_AGEMA_signal_7228) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_7231), .Q (new_AGEMA_signal_7232) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_7235), .Q (new_AGEMA_signal_7236) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_7239), .Q (new_AGEMA_signal_7240) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_7243), .Q (new_AGEMA_signal_7244) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_7247), .Q (new_AGEMA_signal_7248) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_7251), .Q (new_AGEMA_signal_7252) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_7256) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_7260) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_7263), .Q (new_AGEMA_signal_7264) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_7267), .Q (new_AGEMA_signal_7268) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_7271), .Q (new_AGEMA_signal_7272) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_7275), .Q (new_AGEMA_signal_7276) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_7279), .Q (new_AGEMA_signal_7280) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (new_AGEMA_signal_7283), .Q (new_AGEMA_signal_7284) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_7287), .Q (new_AGEMA_signal_7288) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_7292) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_7296) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_7299), .Q (new_AGEMA_signal_7300) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_7303), .Q (new_AGEMA_signal_7304) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_7307), .Q (new_AGEMA_signal_7308) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_7311), .Q (new_AGEMA_signal_7312) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_7315), .Q (new_AGEMA_signal_7316) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_7319), .Q (new_AGEMA_signal_7320) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_7323), .Q (new_AGEMA_signal_7324) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_7328) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_7332) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_7336) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_7339), .Q (new_AGEMA_signal_7340) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_7344) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_7347), .Q (new_AGEMA_signal_7348) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_7351), .Q (new_AGEMA_signal_7352) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_7355), .Q (new_AGEMA_signal_7356) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_7359), .Q (new_AGEMA_signal_7360) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_7363), .Q (new_AGEMA_signal_7364) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_7368) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_7371), .Q (new_AGEMA_signal_7372) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_7376) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_7379), .Q (new_AGEMA_signal_7380) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_7384) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_7387), .Q (new_AGEMA_signal_7388) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_7391), .Q (new_AGEMA_signal_7392) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_7395), .Q (new_AGEMA_signal_7396) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_7399), .Q (new_AGEMA_signal_7400) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_7403), .Q (new_AGEMA_signal_7404) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_7408) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_7411), .Q (new_AGEMA_signal_7412) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_7416) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_7419), .Q (new_AGEMA_signal_7420) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_7424) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_7427), .Q (new_AGEMA_signal_7428) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_7431), .Q (new_AGEMA_signal_7432) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_7435), .Q (new_AGEMA_signal_7436) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_7439), .Q (new_AGEMA_signal_7440) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_7443), .Q (new_AGEMA_signal_7444) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_7448) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_7451), .Q (new_AGEMA_signal_7452) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_7456) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_7459), .Q (new_AGEMA_signal_7460) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_7464) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_7467), .Q (new_AGEMA_signal_7468) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_7471), .Q (new_AGEMA_signal_7472) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_7475), .Q (new_AGEMA_signal_7476) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_7479), .Q (new_AGEMA_signal_7480) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_7483), .Q (new_AGEMA_signal_7484) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_7488) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_7491), .Q (new_AGEMA_signal_7492) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_7496) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_7499), .Q (new_AGEMA_signal_7500) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_7504) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_7507), .Q (new_AGEMA_signal_7508) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_7511), .Q (new_AGEMA_signal_7512) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_7515), .Q (new_AGEMA_signal_7516) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_7519), .Q (new_AGEMA_signal_7520) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_7523), .Q (new_AGEMA_signal_7524) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_7528) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_7531), .Q (new_AGEMA_signal_7532) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_7536) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_7539), .Q (new_AGEMA_signal_7540) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_7543), .Q (new_AGEMA_signal_7544) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_7547), .Q (new_AGEMA_signal_7548) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_7551), .Q (new_AGEMA_signal_7552) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_7555), .Q (new_AGEMA_signal_7556) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_7559), .Q (new_AGEMA_signal_7560) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_7564), .Q (new_AGEMA_signal_7565) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_7568), .Q (new_AGEMA_signal_7569) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_7572), .Q (new_AGEMA_signal_7573) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_7576), .Q (new_AGEMA_signal_7577) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_7580), .Q (new_AGEMA_signal_7581) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_7584), .Q (new_AGEMA_signal_7585) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_7589) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_7592), .Q (new_AGEMA_signal_7593) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_7596), .Q (new_AGEMA_signal_7597) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_7600), .Q (new_AGEMA_signal_7601) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_7604), .Q (new_AGEMA_signal_7605) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_7608), .Q (new_AGEMA_signal_7609) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_7612), .Q (new_AGEMA_signal_7613) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_7617) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_7620), .Q (new_AGEMA_signal_7621) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_7624), .Q (new_AGEMA_signal_7625) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_7628), .Q (new_AGEMA_signal_7629) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_7632), .Q (new_AGEMA_signal_7633) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_7636), .Q (new_AGEMA_signal_7637) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_7640), .Q (new_AGEMA_signal_7641) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_7644), .Q (new_AGEMA_signal_7645) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_7648), .Q (new_AGEMA_signal_7649) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_7652), .Q (new_AGEMA_signal_7653) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_7656), .Q (new_AGEMA_signal_7657) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_7660), .Q (new_AGEMA_signal_7661) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_7664), .Q (new_AGEMA_signal_7665) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_7668), .Q (new_AGEMA_signal_7669) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_7672), .Q (new_AGEMA_signal_7673) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_7676), .Q (new_AGEMA_signal_7677) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_7680), .Q (new_AGEMA_signal_7681) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_7684), .Q (new_AGEMA_signal_7685) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_7688), .Q (new_AGEMA_signal_7689) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_7692), .Q (new_AGEMA_signal_7693) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_7697) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_7700), .Q (new_AGEMA_signal_7701) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_7704), .Q (new_AGEMA_signal_7705) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_7708), .Q (new_AGEMA_signal_7709) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_7712), .Q (new_AGEMA_signal_7713) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_7716), .Q (new_AGEMA_signal_7717) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_7720), .Q (new_AGEMA_signal_7721) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_7724), .Q (new_AGEMA_signal_7725) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_7728), .Q (new_AGEMA_signal_7729) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_7732), .Q (new_AGEMA_signal_7733) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_7736), .Q (new_AGEMA_signal_7737) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_7740), .Q (new_AGEMA_signal_7741) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_7744), .Q (new_AGEMA_signal_7745) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_7748), .Q (new_AGEMA_signal_7749) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_7752), .Q (new_AGEMA_signal_7753) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_7756), .Q (new_AGEMA_signal_7757) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_7760), .Q (new_AGEMA_signal_7761) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_7764), .Q (new_AGEMA_signal_7765) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_7768), .Q (new_AGEMA_signal_7769) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_7772), .Q (new_AGEMA_signal_7773) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_7776), .Q (new_AGEMA_signal_7777) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_7780), .Q (new_AGEMA_signal_7781) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_7784), .Q (new_AGEMA_signal_7785) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_7788), .Q (new_AGEMA_signal_7789) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_7792), .Q (new_AGEMA_signal_7793) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_7796), .Q (new_AGEMA_signal_7797) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_7800), .Q (new_AGEMA_signal_7801) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_7804), .Q (new_AGEMA_signal_7805) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_7808), .Q (new_AGEMA_signal_7809) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_7812), .Q (new_AGEMA_signal_7813) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_7816), .Q (new_AGEMA_signal_7817) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_7820), .Q (new_AGEMA_signal_7821) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_7824), .Q (new_AGEMA_signal_7825) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_7828), .Q (new_AGEMA_signal_7829) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_7832), .Q (new_AGEMA_signal_7833) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_7836), .Q (new_AGEMA_signal_7837) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_7840), .Q (new_AGEMA_signal_7841) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_7844), .Q (new_AGEMA_signal_7845) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_7848), .Q (new_AGEMA_signal_7849) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_7852), .Q (new_AGEMA_signal_7853) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_7856), .Q (new_AGEMA_signal_7857) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_7860), .Q (new_AGEMA_signal_7861) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_7864), .Q (new_AGEMA_signal_7865) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_7868), .Q (new_AGEMA_signal_7869) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_7872), .Q (new_AGEMA_signal_7873) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_7876), .Q (new_AGEMA_signal_7877) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_7880), .Q (new_AGEMA_signal_7881) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_7884), .Q (new_AGEMA_signal_7885) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_7888), .Q (new_AGEMA_signal_7889) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_7892), .Q (new_AGEMA_signal_7893) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_7896), .Q (new_AGEMA_signal_7897) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_7900), .Q (new_AGEMA_signal_7901) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_7904), .Q (new_AGEMA_signal_7905) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_7908), .Q (new_AGEMA_signal_7909) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_7912), .Q (new_AGEMA_signal_7913) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_7916), .Q (new_AGEMA_signal_7917) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_7920), .Q (new_AGEMA_signal_7921) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_7924), .Q (new_AGEMA_signal_7925) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_7928), .Q (new_AGEMA_signal_7929) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_7932), .Q (new_AGEMA_signal_7933) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_7936), .Q (new_AGEMA_signal_7937) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_7940), .Q (new_AGEMA_signal_7941) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_7944), .Q (new_AGEMA_signal_7945) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_6647), .Q (new_AGEMA_signal_7947) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_7948) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_6649), .Q (new_AGEMA_signal_7949) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_7950), .Q (new_AGEMA_signal_7951) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_7952), .Q (new_AGEMA_signal_7953) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_7954), .Q (new_AGEMA_signal_7955) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_6656), .Q (new_AGEMA_signal_7956) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_6657), .Q (new_AGEMA_signal_7957) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (new_AGEMA_signal_6658), .Q (new_AGEMA_signal_7958) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_7959), .Q (new_AGEMA_signal_7960) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (clk), .D (new_AGEMA_signal_7961), .Q (new_AGEMA_signal_7962) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_7963), .Q (new_AGEMA_signal_7964) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_6665), .Q (new_AGEMA_signal_7965) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_6666), .Q (new_AGEMA_signal_7966) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_7967) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_7968), .Q (new_AGEMA_signal_7969) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_7970), .Q (new_AGEMA_signal_7971) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_7972), .Q (new_AGEMA_signal_7973) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_6674), .Q (new_AGEMA_signal_7974) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_6675), .Q (new_AGEMA_signal_7975) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_6676), .Q (new_AGEMA_signal_7976) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (new_AGEMA_signal_7977), .Q (new_AGEMA_signal_7978) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_7979), .Q (new_AGEMA_signal_7980) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (clk), .D (new_AGEMA_signal_7981), .Q (new_AGEMA_signal_7982) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_6683), .Q (new_AGEMA_signal_7983) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_7984) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_6685), .Q (new_AGEMA_signal_7985) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_7986), .Q (new_AGEMA_signal_7987) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_7988), .Q (new_AGEMA_signal_7989) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_7990), .Q (new_AGEMA_signal_7991) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_6692), .Q (new_AGEMA_signal_7992) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_6693), .Q (new_AGEMA_signal_7993) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_6694), .Q (new_AGEMA_signal_7994) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_7995), .Q (new_AGEMA_signal_7996) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (new_AGEMA_signal_7997), .Q (new_AGEMA_signal_7998) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_7999), .Q (new_AGEMA_signal_8000) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_6701), .Q (new_AGEMA_signal_8001) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (clk), .D (new_AGEMA_signal_6702), .Q (new_AGEMA_signal_8002) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_8003) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_8004), .Q (new_AGEMA_signal_8005) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_8006), .Q (new_AGEMA_signal_8007) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_8008), .Q (new_AGEMA_signal_8009) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_6710), .Q (new_AGEMA_signal_8010) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_6711), .Q (new_AGEMA_signal_8011) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_6712), .Q (new_AGEMA_signal_8012) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_8013), .Q (new_AGEMA_signal_8014) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_8015), .Q (new_AGEMA_signal_8016) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C (clk), .D (new_AGEMA_signal_8017), .Q (new_AGEMA_signal_8018) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_6719), .Q (new_AGEMA_signal_8019) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_8020) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_6721), .Q (new_AGEMA_signal_8021) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_8022), .Q (new_AGEMA_signal_8023) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_8024), .Q (new_AGEMA_signal_8025) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_8026), .Q (new_AGEMA_signal_8027) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_6728), .Q (new_AGEMA_signal_8028) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_6729), .Q (new_AGEMA_signal_8029) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_6730), .Q (new_AGEMA_signal_8030) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_8031), .Q (new_AGEMA_signal_8032) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C (clk), .D (new_AGEMA_signal_8033), .Q (new_AGEMA_signal_8034) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_8035), .Q (new_AGEMA_signal_8036) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_6737), .Q (new_AGEMA_signal_8037) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_6738), .Q (new_AGEMA_signal_8038) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_8039) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_8040), .Q (new_AGEMA_signal_8041) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_8042), .Q (new_AGEMA_signal_8043) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_8044), .Q (new_AGEMA_signal_8045) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_6746), .Q (new_AGEMA_signal_8046) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_6747), .Q (new_AGEMA_signal_8047) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_6748), .Q (new_AGEMA_signal_8048) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C (clk), .D (new_AGEMA_signal_8049), .Q (new_AGEMA_signal_8050) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_8051), .Q (new_AGEMA_signal_8052) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_8053), .Q (new_AGEMA_signal_8054) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_6755), .Q (new_AGEMA_signal_8055) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_8056) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_6757), .Q (new_AGEMA_signal_8057) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_8058), .Q (new_AGEMA_signal_8059) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_8060), .Q (new_AGEMA_signal_8061) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_8062), .Q (new_AGEMA_signal_8063) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_6764), .Q (new_AGEMA_signal_8064) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_6765), .Q (new_AGEMA_signal_8065) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C (clk), .D (new_AGEMA_signal_6766), .Q (new_AGEMA_signal_8066) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_8067), .Q (new_AGEMA_signal_8068) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C (clk), .D (new_AGEMA_signal_8069), .Q (new_AGEMA_signal_8070) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_8071), .Q (new_AGEMA_signal_8072) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_6773), .Q (new_AGEMA_signal_8073) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_6774), .Q (new_AGEMA_signal_8074) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_8075) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_8076), .Q (new_AGEMA_signal_8077) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_8078), .Q (new_AGEMA_signal_8079) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_8080), .Q (new_AGEMA_signal_8081) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C (clk), .D (new_AGEMA_signal_6782), .Q (new_AGEMA_signal_8082) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_6783), .Q (new_AGEMA_signal_8083) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_6784), .Q (new_AGEMA_signal_8084) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_8085), .Q (new_AGEMA_signal_8086) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_8087), .Q (new_AGEMA_signal_8088) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_8089), .Q (new_AGEMA_signal_8090) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C (clk), .D (new_AGEMA_signal_8093), .Q (new_AGEMA_signal_8094) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C (clk), .D (new_AGEMA_signal_8097), .Q (new_AGEMA_signal_8098) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_8101), .Q (new_AGEMA_signal_8102) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_8105), .Q (new_AGEMA_signal_8106) ) ;

    /* cells in depth 4 */
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U127 ( .a ({new_AGEMA_signal_6805, new_AGEMA_signal_6801, new_AGEMA_signal_6797}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .c ({DataOut_s2[8], DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U125 ( .a ({new_AGEMA_signal_6817, new_AGEMA_signal_6813, new_AGEMA_signal_6809}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .c ({DataOut_s2[6], DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U123 ( .a ({new_AGEMA_signal_6829, new_AGEMA_signal_6825, new_AGEMA_signal_6821}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .c ({DataOut_s2[62], DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U121 ( .a ({new_AGEMA_signal_6841, new_AGEMA_signal_6837, new_AGEMA_signal_6833}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .c ({DataOut_s2[60], DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U118 ( .a ({new_AGEMA_signal_6853, new_AGEMA_signal_6849, new_AGEMA_signal_6845}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .c ({DataOut_s2[58], DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U116 ( .a ({new_AGEMA_signal_6865, new_AGEMA_signal_6861, new_AGEMA_signal_6857}), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .c ({DataOut_s2[56], DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U114 ( .a ({new_AGEMA_signal_6877, new_AGEMA_signal_6873, new_AGEMA_signal_6869}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .c ({DataOut_s2[54], DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U112 ( .a ({new_AGEMA_signal_6889, new_AGEMA_signal_6885, new_AGEMA_signal_6881}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .c ({DataOut_s2[52], DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U110 ( .a ({new_AGEMA_signal_6901, new_AGEMA_signal_6897, new_AGEMA_signal_6893}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .c ({DataOut_s2[50], DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U109 ( .a ({new_AGEMA_signal_6913, new_AGEMA_signal_6909, new_AGEMA_signal_6905}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .c ({DataOut_s2[4], DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U107 ( .a ({new_AGEMA_signal_6925, new_AGEMA_signal_6921, new_AGEMA_signal_6917}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .c ({DataOut_s2[48], DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U105 ( .a ({new_AGEMA_signal_6937, new_AGEMA_signal_6933, new_AGEMA_signal_6929}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .c ({DataOut_s2[46], DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U103 ( .a ({new_AGEMA_signal_6949, new_AGEMA_signal_6945, new_AGEMA_signal_6941}), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .c ({DataOut_s2[44], DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U101 ( .a ({new_AGEMA_signal_6961, new_AGEMA_signal_6957, new_AGEMA_signal_6953}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .c ({DataOut_s2[42], DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U99 ( .a ({new_AGEMA_signal_6973, new_AGEMA_signal_6969, new_AGEMA_signal_6965}), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .c ({DataOut_s2[40], DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U96 ( .a ({new_AGEMA_signal_6985, new_AGEMA_signal_6981, new_AGEMA_signal_6977}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .c ({DataOut_s2[38], DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U94 ( .a ({new_AGEMA_signal_6997, new_AGEMA_signal_6993, new_AGEMA_signal_6989}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .c ({DataOut_s2[36], DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U92 ( .a ({new_AGEMA_signal_7009, new_AGEMA_signal_7005, new_AGEMA_signal_7001}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .c ({DataOut_s2[34], DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U90 ( .a ({new_AGEMA_signal_7021, new_AGEMA_signal_7017, new_AGEMA_signal_7013}), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .c ({DataOut_s2[32], DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U88 ( .a ({new_AGEMA_signal_7033, new_AGEMA_signal_7029, new_AGEMA_signal_7025}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .c ({DataOut_s2[30], DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U87 ( .a ({new_AGEMA_signal_7045, new_AGEMA_signal_7041, new_AGEMA_signal_7037}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .c ({DataOut_s2[2], DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U85 ( .a ({new_AGEMA_signal_7057, new_AGEMA_signal_7053, new_AGEMA_signal_7049}), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .c ({DataOut_s2[28], DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U83 ( .a ({new_AGEMA_signal_7069, new_AGEMA_signal_7065, new_AGEMA_signal_7061}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .c ({DataOut_s2[26], DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U81 ( .a ({new_AGEMA_signal_7081, new_AGEMA_signal_7077, new_AGEMA_signal_7073}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .c ({DataOut_s2[24], DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U79 ( .a ({new_AGEMA_signal_7093, new_AGEMA_signal_7089, new_AGEMA_signal_7085}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .c ({DataOut_s2[22], DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U77 ( .a ({new_AGEMA_signal_7105, new_AGEMA_signal_7101, new_AGEMA_signal_7097}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .c ({DataOut_s2[20], DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U74 ( .a ({new_AGEMA_signal_7117, new_AGEMA_signal_7113, new_AGEMA_signal_7109}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .c ({DataOut_s2[18], DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U72 ( .a ({new_AGEMA_signal_7129, new_AGEMA_signal_7125, new_AGEMA_signal_7121}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .c ({DataOut_s2[16], DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U70 ( .a ({new_AGEMA_signal_7141, new_AGEMA_signal_7137, new_AGEMA_signal_7133}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .c ({DataOut_s2[14], DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U68 ( .a ({new_AGEMA_signal_7153, new_AGEMA_signal_7149, new_AGEMA_signal_7145}), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .c ({DataOut_s2[12], DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U66 ( .a ({new_AGEMA_signal_7165, new_AGEMA_signal_7161, new_AGEMA_signal_7157}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .c ({DataOut_s2[10], DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_U65 ( .a ({new_AGEMA_signal_7177, new_AGEMA_signal_7173, new_AGEMA_signal_7169}), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .c ({DataOut_s2[0], DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U143 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .b ({new_AGEMA_signal_7189, new_AGEMA_signal_7185, new_AGEMA_signal_7181}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, Midori_rounds_sub_ResultXORkey[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U141 ( .a ({new_AGEMA_signal_7201, new_AGEMA_signal_7197, new_AGEMA_signal_7193}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .c ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, Midori_rounds_sub_ResultXORkey[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U139 ( .a ({new_AGEMA_signal_7213, new_AGEMA_signal_7209, new_AGEMA_signal_7205}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .c ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, Midori_rounds_sub_ResultXORkey[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U137 ( .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .b ({new_AGEMA_signal_7225, new_AGEMA_signal_7221, new_AGEMA_signal_7217}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_sub_ResultXORkey[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U134 ( .a ({new_AGEMA_signal_7237, new_AGEMA_signal_7233, new_AGEMA_signal_7229}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .c ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, Midori_rounds_sub_ResultXORkey[58]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U132 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .b ({new_AGEMA_signal_7249, new_AGEMA_signal_7245, new_AGEMA_signal_7241}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, Midori_rounds_sub_ResultXORkey[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U130 ( .a ({new_AGEMA_signal_7261, new_AGEMA_signal_7257, new_AGEMA_signal_7253}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .c ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, Midori_rounds_sub_ResultXORkey[54]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U128 ( .a ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .b ({new_AGEMA_signal_7273, new_AGEMA_signal_7269, new_AGEMA_signal_7265}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, Midori_rounds_sub_ResultXORkey[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U126 ( .a ({new_AGEMA_signal_7285, new_AGEMA_signal_7281, new_AGEMA_signal_7277}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .c ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, Midori_rounds_sub_ResultXORkey[50]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U125 ( .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .b ({new_AGEMA_signal_7297, new_AGEMA_signal_7293, new_AGEMA_signal_7289}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_sub_ResultXORkey[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U123 ( .a ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .b ({new_AGEMA_signal_7309, new_AGEMA_signal_7305, new_AGEMA_signal_7301}), .c ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, Midori_rounds_sub_ResultXORkey[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U121 ( .a ({new_AGEMA_signal_7321, new_AGEMA_signal_7317, new_AGEMA_signal_7313}), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .c ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, Midori_rounds_sub_ResultXORkey[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U119 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .b ({new_AGEMA_signal_7333, new_AGEMA_signal_7329, new_AGEMA_signal_7325}), .c ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, Midori_rounds_sub_ResultXORkey[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U117 ( .a ({new_AGEMA_signal_7345, new_AGEMA_signal_7341, new_AGEMA_signal_7337}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .c ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, Midori_rounds_sub_ResultXORkey[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U115 ( .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .b ({new_AGEMA_signal_7357, new_AGEMA_signal_7353, new_AGEMA_signal_7349}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, Midori_rounds_sub_ResultXORkey[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U112 ( .a ({new_AGEMA_signal_7369, new_AGEMA_signal_7365, new_AGEMA_signal_7361}), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_sub_ResultXORkey[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U110 ( .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .b ({new_AGEMA_signal_7381, new_AGEMA_signal_7377, new_AGEMA_signal_7373}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_sub_ResultXORkey[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U108 ( .a ({new_AGEMA_signal_7393, new_AGEMA_signal_7389, new_AGEMA_signal_7385}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_sub_ResultXORkey[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U106 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .b ({new_AGEMA_signal_7405, new_AGEMA_signal_7401, new_AGEMA_signal_7397}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, Midori_rounds_sub_ResultXORkey[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U104 ( .a ({new_AGEMA_signal_7417, new_AGEMA_signal_7413, new_AGEMA_signal_7409}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_sub_ResultXORkey[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U103 ( .a ({new_AGEMA_signal_7429, new_AGEMA_signal_7425, new_AGEMA_signal_7421}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, Midori_rounds_sub_ResultXORkey[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U101 ( .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .b ({new_AGEMA_signal_7441, new_AGEMA_signal_7437, new_AGEMA_signal_7433}), .c ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, Midori_rounds_sub_ResultXORkey[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U99 ( .a ({new_AGEMA_signal_7453, new_AGEMA_signal_7449, new_AGEMA_signal_7445}), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, Midori_rounds_sub_ResultXORkey[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U97 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .b ({new_AGEMA_signal_7465, new_AGEMA_signal_7461, new_AGEMA_signal_7457}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_sub_ResultXORkey[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U95 ( .a ({new_AGEMA_signal_7477, new_AGEMA_signal_7473, new_AGEMA_signal_7469}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, Midori_rounds_sub_ResultXORkey[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U93 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7485, new_AGEMA_signal_7481}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, Midori_rounds_sub_ResultXORkey[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U90 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7497, new_AGEMA_signal_7493}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .c ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, Midori_rounds_sub_ResultXORkey[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U88 ( .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7509, new_AGEMA_signal_7505}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, Midori_rounds_sub_ResultXORkey[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U86 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7521, new_AGEMA_signal_7517}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .c ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, Midori_rounds_sub_ResultXORkey[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U84 ( .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7533, new_AGEMA_signal_7529}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, Midori_rounds_sub_ResultXORkey[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U82 ( .a ({new_AGEMA_signal_7549, new_AGEMA_signal_7545, new_AGEMA_signal_7541}), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .c ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, Midori_rounds_sub_ResultXORkey[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U81 ( .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .b ({new_AGEMA_signal_7561, new_AGEMA_signal_7557, new_AGEMA_signal_7553}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_sub_ResultXORkey[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U79 ( .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}), .b ({new_AGEMA_signal_7189, new_AGEMA_signal_7185, new_AGEMA_signal_7181}), .c ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, Midori_rounds_mul_ResultXORkey[8]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U76 ( .a ({new_AGEMA_signal_7201, new_AGEMA_signal_7197, new_AGEMA_signal_7193}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_mul_ResultXORkey[6]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U74 ( .a ({new_AGEMA_signal_7213, new_AGEMA_signal_7209, new_AGEMA_signal_7205}), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, Midori_rounds_mul_ResultXORkey[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U72 ( .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}), .b ({new_AGEMA_signal_7225, new_AGEMA_signal_7221, new_AGEMA_signal_7217}), .c ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, Midori_rounds_mul_ResultXORkey[60]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U68 ( .a ({new_AGEMA_signal_7237, new_AGEMA_signal_7233, new_AGEMA_signal_7229}), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_mul_ResultXORkey[58]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U66 ( .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}), .b ({new_AGEMA_signal_7249, new_AGEMA_signal_7245, new_AGEMA_signal_7241}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, Midori_rounds_mul_ResultXORkey[56]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U63 ( .a ({new_AGEMA_signal_7261, new_AGEMA_signal_7257, new_AGEMA_signal_7253}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_mul_ResultXORkey[54]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U61 ( .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}), .b ({new_AGEMA_signal_7273, new_AGEMA_signal_7269, new_AGEMA_signal_7265}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, Midori_rounds_mul_ResultXORkey[52]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U58 ( .a ({new_AGEMA_signal_7285, new_AGEMA_signal_7281, new_AGEMA_signal_7277}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_mul_ResultXORkey[50]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U57 ( .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}), .b ({new_AGEMA_signal_7297, new_AGEMA_signal_7293, new_AGEMA_signal_7289}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, Midori_rounds_mul_ResultXORkey[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U54 ( .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}), .b ({new_AGEMA_signal_7309, new_AGEMA_signal_7305, new_AGEMA_signal_7301}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, Midori_rounds_mul_ResultXORkey[48]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U51 ( .a ({new_AGEMA_signal_7321, new_AGEMA_signal_7317, new_AGEMA_signal_7313}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_mul_ResultXORkey[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U49 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}), .b ({new_AGEMA_signal_7333, new_AGEMA_signal_7329, new_AGEMA_signal_7325}), .c ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, Midori_rounds_mul_ResultXORkey[44]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U46 ( .a ({new_AGEMA_signal_7345, new_AGEMA_signal_7341, new_AGEMA_signal_7337}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, Midori_rounds_mul_ResultXORkey[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U44 ( .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}), .b ({new_AGEMA_signal_7357, new_AGEMA_signal_7353, new_AGEMA_signal_7349}), .c ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, Midori_rounds_mul_ResultXORkey[40]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U40 ( .a ({new_AGEMA_signal_7369, new_AGEMA_signal_7365, new_AGEMA_signal_7361}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, Midori_rounds_mul_ResultXORkey[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U38 ( .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}), .b ({new_AGEMA_signal_7381, new_AGEMA_signal_7377, new_AGEMA_signal_7373}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, Midori_rounds_mul_ResultXORkey[36]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U35 ( .a ({new_AGEMA_signal_7393, new_AGEMA_signal_7389, new_AGEMA_signal_7385}), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_mul_ResultXORkey[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U33 ( .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}), .b ({new_AGEMA_signal_7405, new_AGEMA_signal_7401, new_AGEMA_signal_7397}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, Midori_rounds_mul_ResultXORkey[32]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U30 ( .a ({new_AGEMA_signal_7417, new_AGEMA_signal_7413, new_AGEMA_signal_7409}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_mul_ResultXORkey[30]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U29 ( .a ({new_AGEMA_signal_7429, new_AGEMA_signal_7425, new_AGEMA_signal_7421}), .b ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, Midori_rounds_mul_ResultXORkey[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U27 ( .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}), .b ({new_AGEMA_signal_7441, new_AGEMA_signal_7437, new_AGEMA_signal_7433}), .c ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, Midori_rounds_mul_ResultXORkey[28]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U24 ( .a ({new_AGEMA_signal_7453, new_AGEMA_signal_7449, new_AGEMA_signal_7445}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, Midori_rounds_mul_ResultXORkey[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U22 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}), .b ({new_AGEMA_signal_7465, new_AGEMA_signal_7461, new_AGEMA_signal_7457}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, Midori_rounds_mul_ResultXORkey[24]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U19 ( .a ({new_AGEMA_signal_7477, new_AGEMA_signal_7473, new_AGEMA_signal_7469}), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, Midori_rounds_mul_ResultXORkey[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U17 ( .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7485, new_AGEMA_signal_7481}), .c ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, Midori_rounds_mul_ResultXORkey[20]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U13 ( .a ({new_AGEMA_signal_7501, new_AGEMA_signal_7497, new_AGEMA_signal_7493}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_mul_ResultXORkey[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U11 ( .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7509, new_AGEMA_signal_7505}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, Midori_rounds_mul_ResultXORkey[16]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U8 ( .a ({new_AGEMA_signal_7525, new_AGEMA_signal_7521, new_AGEMA_signal_7517}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_mul_ResultXORkey[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U6 ( .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7533, new_AGEMA_signal_7529}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, Midori_rounds_mul_ResultXORkey[12]}) ) ;
    xor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U3 ( .a ({new_AGEMA_signal_7549, new_AGEMA_signal_7545, new_AGEMA_signal_7541}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_mul_ResultXORkey[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_U2 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}), .b ({new_AGEMA_signal_7561, new_AGEMA_signal_7557, new_AGEMA_signal_7553}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, Midori_rounds_mul_ResultXORkey[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, Midori_rounds_round_Result[0]}), .a ({new_AGEMA_signal_7574, new_AGEMA_signal_7570, new_AGEMA_signal_7566}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_roundResult_Reg_SFF_0_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, Midori_rounds_round_Result[2]}), .a ({new_AGEMA_signal_7586, new_AGEMA_signal_7582, new_AGEMA_signal_7578}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_roundResult_Reg_SFF_2_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, Midori_rounds_round_Result[4]}), .a ({new_AGEMA_signal_7598, new_AGEMA_signal_7594, new_AGEMA_signal_7590}), .c ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, Midori_rounds_roundResult_Reg_SFF_4_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, Midori_rounds_round_Result[6]}), .a ({new_AGEMA_signal_7610, new_AGEMA_signal_7606, new_AGEMA_signal_7602}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_roundResult_Reg_SFF_6_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, Midori_rounds_round_Result[8]}), .a ({new_AGEMA_signal_7622, new_AGEMA_signal_7618, new_AGEMA_signal_7614}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, Midori_rounds_roundResult_Reg_SFF_8_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, Midori_rounds_round_Result[10]}), .a ({new_AGEMA_signal_7634, new_AGEMA_signal_7630, new_AGEMA_signal_7626}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_roundResult_Reg_SFF_10_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, Midori_rounds_round_Result[12]}), .a ({new_AGEMA_signal_7646, new_AGEMA_signal_7642, new_AGEMA_signal_7638}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_roundResult_Reg_SFF_12_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, Midori_rounds_round_Result[14]}), .a ({new_AGEMA_signal_7658, new_AGEMA_signal_7654, new_AGEMA_signal_7650}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_roundResult_Reg_SFF_14_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, Midori_rounds_round_Result[16]}), .a ({new_AGEMA_signal_7670, new_AGEMA_signal_7666, new_AGEMA_signal_7662}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, Midori_rounds_roundResult_Reg_SFF_16_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, Midori_rounds_round_Result[18]}), .a ({new_AGEMA_signal_7682, new_AGEMA_signal_7678, new_AGEMA_signal_7674}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_roundResult_Reg_SFF_18_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_round_Result[20]}), .a ({new_AGEMA_signal_7694, new_AGEMA_signal_7690, new_AGEMA_signal_7686}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_roundResult_Reg_SFF_20_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, Midori_rounds_round_Result[22]}), .a ({new_AGEMA_signal_7706, new_AGEMA_signal_7702, new_AGEMA_signal_7698}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_roundResult_Reg_SFF_22_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, Midori_rounds_round_Result[24]}), .a ({new_AGEMA_signal_7718, new_AGEMA_signal_7714, new_AGEMA_signal_7710}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, Midori_rounds_roundResult_Reg_SFF_24_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, Midori_rounds_round_Result[26]}), .a ({new_AGEMA_signal_7730, new_AGEMA_signal_7726, new_AGEMA_signal_7722}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, Midori_rounds_roundResult_Reg_SFF_26_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, Midori_rounds_round_Result[28]}), .a ({new_AGEMA_signal_7742, new_AGEMA_signal_7738, new_AGEMA_signal_7734}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, Midori_rounds_roundResult_Reg_SFF_28_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, Midori_rounds_round_Result[30]}), .a ({new_AGEMA_signal_7754, new_AGEMA_signal_7750, new_AGEMA_signal_7746}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, Midori_rounds_roundResult_Reg_SFF_30_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, Midori_rounds_round_Result[32]}), .a ({new_AGEMA_signal_7766, new_AGEMA_signal_7762, new_AGEMA_signal_7758}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_roundResult_Reg_SFF_32_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, Midori_rounds_round_Result[34]}), .a ({new_AGEMA_signal_7778, new_AGEMA_signal_7774, new_AGEMA_signal_7770}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, Midori_rounds_roundResult_Reg_SFF_34_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, Midori_rounds_round_Result[36]}), .a ({new_AGEMA_signal_7790, new_AGEMA_signal_7786, new_AGEMA_signal_7782}), .c ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, Midori_rounds_roundResult_Reg_SFF_36_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, Midori_rounds_round_Result[38]}), .a ({new_AGEMA_signal_7802, new_AGEMA_signal_7798, new_AGEMA_signal_7794}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, Midori_rounds_roundResult_Reg_SFF_38_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, Midori_rounds_round_Result[40]}), .a ({new_AGEMA_signal_7814, new_AGEMA_signal_7810, new_AGEMA_signal_7806}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, Midori_rounds_roundResult_Reg_SFF_40_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, Midori_rounds_round_Result[42]}), .a ({new_AGEMA_signal_7826, new_AGEMA_signal_7822, new_AGEMA_signal_7818}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, Midori_rounds_roundResult_Reg_SFF_42_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, Midori_rounds_round_Result[44]}), .a ({new_AGEMA_signal_7838, new_AGEMA_signal_7834, new_AGEMA_signal_7830}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_roundResult_Reg_SFF_44_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, Midori_rounds_round_Result[46]}), .a ({new_AGEMA_signal_7850, new_AGEMA_signal_7846, new_AGEMA_signal_7842}), .c ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, Midori_rounds_roundResult_Reg_SFF_46_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_round_Result[48]}), .a ({new_AGEMA_signal_7862, new_AGEMA_signal_7858, new_AGEMA_signal_7854}), .c ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, Midori_rounds_roundResult_Reg_SFF_48_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, Midori_rounds_round_Result[50]}), .a ({new_AGEMA_signal_7874, new_AGEMA_signal_7870, new_AGEMA_signal_7866}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, Midori_rounds_roundResult_Reg_SFF_50_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, Midori_rounds_round_Result[52]}), .a ({new_AGEMA_signal_7886, new_AGEMA_signal_7882, new_AGEMA_signal_7878}), .c ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, Midori_rounds_roundResult_Reg_SFF_52_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, Midori_rounds_round_Result[54]}), .a ({new_AGEMA_signal_7898, new_AGEMA_signal_7894, new_AGEMA_signal_7890}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, Midori_rounds_roundResult_Reg_SFF_54_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, Midori_rounds_round_Result[56]}), .a ({new_AGEMA_signal_7910, new_AGEMA_signal_7906, new_AGEMA_signal_7902}), .c ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, Midori_rounds_roundResult_Reg_SFF_56_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, Midori_rounds_round_Result[58]}), .a ({new_AGEMA_signal_7922, new_AGEMA_signal_7918, new_AGEMA_signal_7914}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Midori_rounds_roundResult_Reg_SFF_58_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_round_Result[60]}), .a ({new_AGEMA_signal_7934, new_AGEMA_signal_7930, new_AGEMA_signal_7926}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, Midori_rounds_roundResult_Reg_SFF_60_DQ}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1 ( .s (new_AGEMA_signal_7562), .b ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, Midori_rounds_round_Result[62]}), .a ({new_AGEMA_signal_7946, new_AGEMA_signal_7942, new_AGEMA_signal_7938}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Midori_rounds_roundResult_Reg_SFF_62_DQ}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .a ({new_AGEMA_signal_7949, new_AGEMA_signal_7948, new_AGEMA_signal_7947}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, Midori_rounds_sub_sBox_PRINCE_0_n12}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .a ({new_AGEMA_signal_7955, new_AGEMA_signal_7953, new_AGEMA_signal_7951}), .b ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, Midori_rounds_sub_sBox_PRINCE_0_n3}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .a ({new_AGEMA_signal_7958, new_AGEMA_signal_7957, new_AGEMA_signal_7956}), .b ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, Midori_rounds_sub_sBox_PRINCE_1_n12}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .a ({new_AGEMA_signal_7964, new_AGEMA_signal_7962, new_AGEMA_signal_7960}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2690, Midori_rounds_sub_sBox_PRINCE_1_n3}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .a ({new_AGEMA_signal_7967, new_AGEMA_signal_7966, new_AGEMA_signal_7965}), .b ({new_AGEMA_signal_2697, new_AGEMA_signal_2696, Midori_rounds_sub_sBox_PRINCE_2_n12}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .a ({new_AGEMA_signal_7973, new_AGEMA_signal_7971, new_AGEMA_signal_7969}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, Midori_rounds_sub_sBox_PRINCE_2_n3}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .a ({new_AGEMA_signal_7976, new_AGEMA_signal_7975, new_AGEMA_signal_7974}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, Midori_rounds_sub_sBox_PRINCE_3_n12}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .a ({new_AGEMA_signal_7982, new_AGEMA_signal_7980, new_AGEMA_signal_7978}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, Midori_rounds_sub_sBox_PRINCE_3_n3}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .a ({new_AGEMA_signal_7985, new_AGEMA_signal_7984, new_AGEMA_signal_7983}), .b ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, Midori_rounds_sub_sBox_PRINCE_4_n12}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .a ({new_AGEMA_signal_7991, new_AGEMA_signal_7989, new_AGEMA_signal_7987}), .b ({new_AGEMA_signal_2721, new_AGEMA_signal_2720, Midori_rounds_sub_sBox_PRINCE_4_n3}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .a ({new_AGEMA_signal_7994, new_AGEMA_signal_7993, new_AGEMA_signal_7992}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, Midori_rounds_sub_sBox_PRINCE_5_n12}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .a ({new_AGEMA_signal_8000, new_AGEMA_signal_7998, new_AGEMA_signal_7996}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, Midori_rounds_sub_sBox_PRINCE_5_n3}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .a ({new_AGEMA_signal_8003, new_AGEMA_signal_8002, new_AGEMA_signal_8001}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, Midori_rounds_sub_sBox_PRINCE_6_n12}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .a ({new_AGEMA_signal_8009, new_AGEMA_signal_8007, new_AGEMA_signal_8005}), .b ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, Midori_rounds_sub_sBox_PRINCE_6_n3}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .a ({new_AGEMA_signal_8012, new_AGEMA_signal_8011, new_AGEMA_signal_8010}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, Midori_rounds_sub_sBox_PRINCE_7_n12}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .a ({new_AGEMA_signal_8018, new_AGEMA_signal_8016, new_AGEMA_signal_8014}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, Midori_rounds_sub_sBox_PRINCE_7_n3}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .a ({new_AGEMA_signal_8021, new_AGEMA_signal_8020, new_AGEMA_signal_8019}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, Midori_rounds_sub_sBox_PRINCE_8_n12}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .a ({new_AGEMA_signal_8027, new_AGEMA_signal_8025, new_AGEMA_signal_8023}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, Midori_rounds_sub_sBox_PRINCE_8_n3}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .a ({new_AGEMA_signal_8030, new_AGEMA_signal_8029, new_AGEMA_signal_8028}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, Midori_rounds_sub_sBox_PRINCE_9_n12}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .a ({new_AGEMA_signal_8036, new_AGEMA_signal_8034, new_AGEMA_signal_8032}), .b ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, Midori_rounds_sub_sBox_PRINCE_9_n3}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .a ({new_AGEMA_signal_8039, new_AGEMA_signal_8038, new_AGEMA_signal_8037}), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, Midori_rounds_sub_sBox_PRINCE_10_n12}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .a ({new_AGEMA_signal_8045, new_AGEMA_signal_8043, new_AGEMA_signal_8041}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, Midori_rounds_sub_sBox_PRINCE_10_n3}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .a ({new_AGEMA_signal_8048, new_AGEMA_signal_8047, new_AGEMA_signal_8046}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, Midori_rounds_sub_sBox_PRINCE_11_n12}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .a ({new_AGEMA_signal_8054, new_AGEMA_signal_8052, new_AGEMA_signal_8050}), .b ({new_AGEMA_signal_2791, new_AGEMA_signal_2790, Midori_rounds_sub_sBox_PRINCE_11_n3}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .a ({new_AGEMA_signal_8057, new_AGEMA_signal_8056, new_AGEMA_signal_8055}), .b ({new_AGEMA_signal_2797, new_AGEMA_signal_2796, Midori_rounds_sub_sBox_PRINCE_12_n12}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .a ({new_AGEMA_signal_8063, new_AGEMA_signal_8061, new_AGEMA_signal_8059}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, Midori_rounds_sub_sBox_PRINCE_12_n3}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .a ({new_AGEMA_signal_8066, new_AGEMA_signal_8065, new_AGEMA_signal_8064}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, Midori_rounds_sub_sBox_PRINCE_13_n12}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .a ({new_AGEMA_signal_8072, new_AGEMA_signal_8070, new_AGEMA_signal_8068}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, Midori_rounds_sub_sBox_PRINCE_13_n3}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .a ({new_AGEMA_signal_8075, new_AGEMA_signal_8074, new_AGEMA_signal_8073}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, Midori_rounds_sub_sBox_PRINCE_14_n12}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .a ({new_AGEMA_signal_8081, new_AGEMA_signal_8079, new_AGEMA_signal_8077}), .b ({new_AGEMA_signal_2821, new_AGEMA_signal_2820, Midori_rounds_sub_sBox_PRINCE_14_n3}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}) ) ;
    nand_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .a ({new_AGEMA_signal_8084, new_AGEMA_signal_8083, new_AGEMA_signal_8082}), .b ({new_AGEMA_signal_2827, new_AGEMA_signal_2826, Midori_rounds_sub_sBox_PRINCE_15_n12}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}) ) ;
    nor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .a ({new_AGEMA_signal_8090, new_AGEMA_signal_8088, new_AGEMA_signal_8086}), .b ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, Midori_rounds_sub_sBox_PRINCE_15_n3}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_0_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2895, new_AGEMA_signal_2894, Midori_rounds_SR_Result[0]}), .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, Midori_rounds_sub_ResultXORkey[0]}), .c ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_2_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, Midori_rounds_SR_Result[2]}), .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, Midori_rounds_sub_ResultXORkey[2]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_4_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, Midori_rounds_SR_Result[4]}), .a ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, Midori_rounds_sub_ResultXORkey[4]}), .c ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_6_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, Midori_rounds_SR_Result[6]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, Midori_rounds_sub_ResultXORkey[6]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_8_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, Midori_rounds_SR_Result[8]}), .a ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, Midori_rounds_sub_ResultXORkey[8]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_10_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2851, new_AGEMA_signal_2850, Midori_rounds_SR_Result[10]}), .a ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, Midori_rounds_sub_ResultXORkey[10]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_12_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, Midori_rounds_SR_Result[12]}), .a ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, Midori_rounds_sub_ResultXORkey[12]}), .c ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_14_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, Midori_rounds_SR_Result[14]}), .a ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, Midori_rounds_sub_ResultXORkey[14]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_16_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, Midori_rounds_SR_Result[16]}), .a ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, Midori_rounds_sub_ResultXORkey[16]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_18_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2907, new_AGEMA_signal_2906, Midori_rounds_SR_Result[18]}), .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, Midori_rounds_sub_ResultXORkey[18]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_20_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2863, new_AGEMA_signal_2862, Midori_rounds_SR_Result[20]}), .a ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, Midori_rounds_sub_ResultXORkey[20]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_22_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, Midori_rounds_SR_Result[22]}), .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, Midori_rounds_sub_ResultXORkey[22]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_24_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, Midori_rounds_SR_Result[24]}), .a ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, Midori_rounds_sub_ResultXORkey[24]}), .c ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_26_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, Midori_rounds_SR_Result[26]}), .a ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, Midori_rounds_sub_ResultXORkey[26]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_28_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, Midori_rounds_SR_Result[28]}), .a ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, Midori_rounds_sub_ResultXORkey[28]}), .c ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_30_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2883, new_AGEMA_signal_2882, Midori_rounds_SR_Result[30]}), .a ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, Midori_rounds_sub_ResultXORkey[30]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_32_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, Midori_rounds_SR_Result[32]}), .a ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, Midori_rounds_sub_ResultXORkey[32]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_34_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, Midori_rounds_SR_Result[34]}), .a ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, Midori_rounds_sub_ResultXORkey[34]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_36_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, Midori_rounds_SR_Result[36]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, Midori_rounds_sub_ResultXORkey[36]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_38_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, Midori_rounds_SR_Result[38]}), .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, Midori_rounds_sub_ResultXORkey[38]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_40_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, Midori_rounds_SR_Result[40]}), .a ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, Midori_rounds_sub_ResultXORkey[40]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_42_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, Midori_rounds_SR_Result[42]}), .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, Midori_rounds_sub_ResultXORkey[42]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_44_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, Midori_rounds_SR_Result[44]}), .a ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, Midori_rounds_sub_ResultXORkey[44]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_46_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, Midori_rounds_SR_Result[46]}), .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, Midori_rounds_sub_ResultXORkey[46]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_48_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2839, new_AGEMA_signal_2838, Midori_rounds_SR_Result[48]}), .a ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, Midori_rounds_sub_ResultXORkey[48]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_50_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, Midori_rounds_SR_Result[50]}), .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, Midori_rounds_sub_ResultXORkey[50]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_52_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2919, new_AGEMA_signal_2918, Midori_rounds_SR_Result[52]}), .a ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, Midori_rounds_sub_ResultXORkey[52]}), .c ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_54_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, Midori_rounds_SR_Result[54]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, Midori_rounds_sub_ResultXORkey[54]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_56_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, Midori_rounds_SR_Result[56]}), .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, Midori_rounds_sub_ResultXORkey[56]}), .c ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_58_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, Midori_rounds_SR_Result[58]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, Midori_rounds_sub_ResultXORkey[58]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_60_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, Midori_rounds_SR_Result[60]}), .a ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, Midori_rounds_sub_ResultXORkey[60]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_62_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, Midori_rounds_SR_Result[62]}), .a ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, Midori_rounds_sub_ResultXORkey[62]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U23 ( .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U21 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U19 ( .a ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U16 ( .a ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U15 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, Midori_rounds_mul_MC1_n5}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U11 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, Midori_rounds_mul_input[58]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U8 ( .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U7 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, Midori_rounds_mul_input[48]}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, Midori_rounds_mul_MC1_n7}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U4 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U3 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, Midori_rounds_mul_input[54]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, Midori_rounds_mul_MC1_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U2 ( .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC1_U1 ( .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, Midori_rounds_mul_input[56]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, Midori_rounds_mul_MC1_n3}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U23 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U21 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U19 ( .a ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U16 ( .a ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U15 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, Midori_rounds_mul_MC2_n5}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U11 ( .a ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, Midori_rounds_mul_input[42]}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U8 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}), .b ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U7 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, Midori_rounds_mul_input[32]}), .c ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, Midori_rounds_mul_MC2_n7}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U4 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U3 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, Midori_rounds_mul_input[38]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, Midori_rounds_mul_MC2_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U2 ( .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC2_U1 ( .a ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, Midori_rounds_mul_input[40]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, Midori_rounds_mul_MC2_n3}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U23 ( .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U21 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U19 ( .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U16 ( .a ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U15 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, Midori_rounds_mul_MC3_n5}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U11 ( .a ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, Midori_rounds_mul_input[26]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U8 ( .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}), .b ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U7 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, Midori_rounds_mul_input[16]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, Midori_rounds_mul_MC3_n7}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U4 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U3 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, Midori_rounds_mul_input[22]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, Midori_rounds_mul_MC3_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U2 ( .a ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC3_U1 ( .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, Midori_rounds_mul_input[24]}), .c ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, Midori_rounds_mul_MC3_n3}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U23 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U21 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U19 ( .a ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U16 ( .a ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U15 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, Midori_rounds_mul_MC4_n5}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U11 ( .a ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, Midori_rounds_mul_input[10]}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U8 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}), .b ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U7 ( .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, Midori_rounds_mul_input[0]}), .c ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, Midori_rounds_mul_MC4_n7}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U4 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U3 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, Midori_rounds_mul_input[6]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, Midori_rounds_mul_MC4_n1}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U2 ( .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}) ) ;
    xnor_HPC3 #(.security_order(2), .pipeline(1)) Midori_rounds_mul_MC4_U1 ( .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Midori_rounds_mul_input[8]}), .c ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, Midori_rounds_mul_MC4_n3}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_0_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, Midori_rounds_mul_ResultXORkey[0]}), .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, Midori_rounds_SR_Inv_Result[0]}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, Midori_rounds_round_Result[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_2_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, Midori_rounds_mul_ResultXORkey[2]}), .a ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, Midori_rounds_round_Result[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_4_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, Midori_rounds_mul_ResultXORkey[4]}), .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, Midori_rounds_SR_Inv_Result[4]}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, Midori_rounds_round_Result[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_6_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, Midori_rounds_mul_ResultXORkey[6]}), .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, Midori_rounds_round_Result[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_8_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, Midori_rounds_mul_ResultXORkey[8]}), .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, Midori_rounds_SR_Inv_Result[8]}), .c ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, Midori_rounds_round_Result[8]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_10_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, Midori_rounds_mul_ResultXORkey[10]}), .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, Midori_rounds_round_Result[10]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_12_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, Midori_rounds_mul_ResultXORkey[12]}), .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, Midori_rounds_SR_Inv_Result[12]}), .c ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, Midori_rounds_round_Result[12]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_14_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, Midori_rounds_mul_ResultXORkey[14]}), .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, Midori_rounds_round_Result[14]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_16_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, Midori_rounds_mul_ResultXORkey[16]}), .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, Midori_rounds_SR_Inv_Result[16]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, Midori_rounds_round_Result[16]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_18_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, Midori_rounds_mul_ResultXORkey[18]}), .a ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, Midori_rounds_round_Result[18]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_20_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, Midori_rounds_mul_ResultXORkey[20]}), .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, Midori_rounds_SR_Inv_Result[20]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, Midori_rounds_round_Result[20]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_22_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, Midori_rounds_mul_ResultXORkey[22]}), .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, Midori_rounds_round_Result[22]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_24_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, Midori_rounds_mul_ResultXORkey[24]}), .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, Midori_rounds_SR_Inv_Result[24]}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, Midori_rounds_round_Result[24]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_26_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, Midori_rounds_mul_ResultXORkey[26]}), .a ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, Midori_rounds_round_Result[26]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_28_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, Midori_rounds_mul_ResultXORkey[28]}), .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, Midori_rounds_SR_Inv_Result[28]}), .c ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, Midori_rounds_round_Result[28]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_30_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, Midori_rounds_mul_ResultXORkey[30]}), .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, Midori_rounds_round_Result[30]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_32_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, Midori_rounds_mul_ResultXORkey[32]}), .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, Midori_rounds_SR_Inv_Result[32]}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, Midori_rounds_round_Result[32]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_34_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, Midori_rounds_mul_ResultXORkey[34]}), .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, Midori_rounds_round_Result[34]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_36_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, Midori_rounds_mul_ResultXORkey[36]}), .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, Midori_rounds_SR_Inv_Result[36]}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, Midori_rounds_round_Result[36]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_38_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, Midori_rounds_mul_ResultXORkey[38]}), .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, Midori_rounds_round_Result[38]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_40_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, Midori_rounds_mul_ResultXORkey[40]}), .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, Midori_rounds_SR_Inv_Result[40]}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, Midori_rounds_round_Result[40]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_42_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, Midori_rounds_mul_ResultXORkey[42]}), .a ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, Midori_rounds_round_Result[42]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_44_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, Midori_rounds_mul_ResultXORkey[44]}), .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, Midori_rounds_SR_Inv_Result[44]}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, Midori_rounds_round_Result[44]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_46_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, Midori_rounds_mul_ResultXORkey[46]}), .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, Midori_rounds_round_Result[46]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_48_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, Midori_rounds_mul_ResultXORkey[48]}), .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, Midori_rounds_SR_Inv_Result[48]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, Midori_rounds_round_Result[48]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_50_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, Midori_rounds_mul_ResultXORkey[50]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, Midori_rounds_round_Result[50]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_52_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, Midori_rounds_mul_ResultXORkey[52]}), .a ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, Midori_rounds_SR_Inv_Result[52]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, Midori_rounds_round_Result[52]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_54_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, Midori_rounds_mul_ResultXORkey[54]}), .a ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, Midori_rounds_round_Result[54]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_56_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, Midori_rounds_mul_ResultXORkey[56]}), .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, Midori_rounds_SR_Inv_Result[56]}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, Midori_rounds_round_Result[56]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_58_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, Midori_rounds_mul_ResultXORkey[58]}), .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, Midori_rounds_round_Result[58]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_60_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, Midori_rounds_mul_ResultXORkey[60]}), .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, Midori_rounds_SR_Inv_Result[60]}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, Midori_rounds_round_Result[60]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_62_U1 ( .s (new_AGEMA_signal_8091), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, Midori_rounds_mul_ResultXORkey[62]}), .a ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, Midori_rounds_round_Result[62]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (DataOut_s0[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (new_AGEMA_signal_5489), .Q (DataOut_s0[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (DataOut_s0[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (DataOut_s0[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (DataOut_s0[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_5493), .Q (DataOut_s0[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (DataOut_s0[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (new_AGEMA_signal_5495), .Q (DataOut_s0[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (DataOut_s0[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (DataOut_s0[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (DataOut_s0[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (DataOut_s0[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (DataOut_s0[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_5501), .Q (DataOut_s0[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (DataOut_s0[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (DataOut_s0[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (DataOut_s0[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_5505), .Q (DataOut_s0[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (DataOut_s0[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (DataOut_s0[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (DataOut_s0[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_5509), .Q (DataOut_s0[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_5510), .Q (DataOut_s0[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (DataOut_s0[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (DataOut_s0[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_5513), .Q (DataOut_s0[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_5514), .Q (DataOut_s0[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (DataOut_s0[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (DataOut_s0[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (DataOut_s0[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (DataOut_s0[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (DataOut_s0[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (done) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (DataOut_s1[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_5525), .Q (DataOut_s2[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (DataOut_s1[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (DataOut_s2[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (DataOut_s1[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_5529), .Q (DataOut_s2[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_5530), .Q (DataOut_s1[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (new_AGEMA_signal_5531), .Q (DataOut_s2[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (DataOut_s1[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (DataOut_s2[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (DataOut_s1[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (DataOut_s2[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (DataOut_s1[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_5537), .Q (DataOut_s2[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_5538), .Q (DataOut_s1[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (DataOut_s2[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (DataOut_s1[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (DataOut_s2[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (DataOut_s1[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (DataOut_s2[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (DataOut_s1[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_5545), .Q (DataOut_s2[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_5546), .Q (DataOut_s1[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_5547), .Q (DataOut_s2[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (DataOut_s1[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_5549), .Q (DataOut_s2[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_5550), .Q (DataOut_s1[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (DataOut_s2[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (DataOut_s1[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (DataOut_s2[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_5554), .Q (DataOut_s1[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (new_AGEMA_signal_5555), .Q (DataOut_s2[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (DataOut_s1[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_5557), .Q (DataOut_s2[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (DataOut_s1[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (DataOut_s2[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (DataOut_s1[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_5561), .Q (DataOut_s2[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (DataOut_s1[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (DataOut_s2[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (DataOut_s1[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_5565), .Q (DataOut_s2[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_5566), .Q (DataOut_s1[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_5567), .Q (DataOut_s2[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (DataOut_s1[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_5569), .Q (DataOut_s2[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_5570), .Q (DataOut_s1[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (DataOut_s2[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (DataOut_s1[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_5573), .Q (DataOut_s2[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_5574), .Q (DataOut_s1[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (DataOut_s2[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (DataOut_s1[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_5577), .Q (DataOut_s2[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (DataOut_s1[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (DataOut_s2[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (DataOut_s1[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (DataOut_s2[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (DataOut_s1[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (DataOut_s2[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (DataOut_s1[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_5585), .Q (DataOut_s2[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_5586), .Q (DataOut_s1[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (DataOut_s2[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_6796), .Q (new_AGEMA_signal_6797) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_6800), .Q (new_AGEMA_signal_6801) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_6804), .Q (new_AGEMA_signal_6805) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_6808), .Q (new_AGEMA_signal_6809) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_6812), .Q (new_AGEMA_signal_6813) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_6816), .Q (new_AGEMA_signal_6817) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_6820), .Q (new_AGEMA_signal_6821) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_6824), .Q (new_AGEMA_signal_6825) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_6829) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_6832), .Q (new_AGEMA_signal_6833) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_6836), .Q (new_AGEMA_signal_6837) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_6840), .Q (new_AGEMA_signal_6841) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_6844), .Q (new_AGEMA_signal_6845) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_6848), .Q (new_AGEMA_signal_6849) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_6852), .Q (new_AGEMA_signal_6853) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_6856), .Q (new_AGEMA_signal_6857) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_6860), .Q (new_AGEMA_signal_6861) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_6865) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_6868), .Q (new_AGEMA_signal_6869) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_6872), .Q (new_AGEMA_signal_6873) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_6876), .Q (new_AGEMA_signal_6877) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_6880), .Q (new_AGEMA_signal_6881) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_6884), .Q (new_AGEMA_signal_6885) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_6888), .Q (new_AGEMA_signal_6889) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_6892), .Q (new_AGEMA_signal_6893) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_6896), .Q (new_AGEMA_signal_6897) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_6900), .Q (new_AGEMA_signal_6901) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_6904), .Q (new_AGEMA_signal_6905) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_6908), .Q (new_AGEMA_signal_6909) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_6912), .Q (new_AGEMA_signal_6913) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_6916), .Q (new_AGEMA_signal_6917) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_6920), .Q (new_AGEMA_signal_6921) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_6924), .Q (new_AGEMA_signal_6925) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_6928), .Q (new_AGEMA_signal_6929) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_6932), .Q (new_AGEMA_signal_6933) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_6936), .Q (new_AGEMA_signal_6937) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_6940), .Q (new_AGEMA_signal_6941) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_6944), .Q (new_AGEMA_signal_6945) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_6948), .Q (new_AGEMA_signal_6949) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_6952), .Q (new_AGEMA_signal_6953) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_6956), .Q (new_AGEMA_signal_6957) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_6960), .Q (new_AGEMA_signal_6961) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_6964), .Q (new_AGEMA_signal_6965) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_6968), .Q (new_AGEMA_signal_6969) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_6972), .Q (new_AGEMA_signal_6973) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_6976), .Q (new_AGEMA_signal_6977) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_6980), .Q (new_AGEMA_signal_6981) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_6984), .Q (new_AGEMA_signal_6985) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_6988), .Q (new_AGEMA_signal_6989) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_6992), .Q (new_AGEMA_signal_6993) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_6996), .Q (new_AGEMA_signal_6997) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_7000), .Q (new_AGEMA_signal_7001) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_7004), .Q (new_AGEMA_signal_7005) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_7008), .Q (new_AGEMA_signal_7009) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_7012), .Q (new_AGEMA_signal_7013) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_7016), .Q (new_AGEMA_signal_7017) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_7020), .Q (new_AGEMA_signal_7021) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_7024), .Q (new_AGEMA_signal_7025) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_7028), .Q (new_AGEMA_signal_7029) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_7032), .Q (new_AGEMA_signal_7033) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_7036), .Q (new_AGEMA_signal_7037) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_7040), .Q (new_AGEMA_signal_7041) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_7044), .Q (new_AGEMA_signal_7045) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_7048), .Q (new_AGEMA_signal_7049) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_7052), .Q (new_AGEMA_signal_7053) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_7056), .Q (new_AGEMA_signal_7057) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_7060), .Q (new_AGEMA_signal_7061) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_7064), .Q (new_AGEMA_signal_7065) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_7068), .Q (new_AGEMA_signal_7069) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_7072), .Q (new_AGEMA_signal_7073) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_7076), .Q (new_AGEMA_signal_7077) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_7080), .Q (new_AGEMA_signal_7081) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_7084), .Q (new_AGEMA_signal_7085) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_7088), .Q (new_AGEMA_signal_7089) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_7092), .Q (new_AGEMA_signal_7093) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_7096), .Q (new_AGEMA_signal_7097) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_7100), .Q (new_AGEMA_signal_7101) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_7104), .Q (new_AGEMA_signal_7105) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_7108), .Q (new_AGEMA_signal_7109) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_7112), .Q (new_AGEMA_signal_7113) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_7116), .Q (new_AGEMA_signal_7117) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_7120), .Q (new_AGEMA_signal_7121) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_7124), .Q (new_AGEMA_signal_7125) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_7128), .Q (new_AGEMA_signal_7129) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_7132), .Q (new_AGEMA_signal_7133) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_7136), .Q (new_AGEMA_signal_7137) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_7140), .Q (new_AGEMA_signal_7141) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_7144), .Q (new_AGEMA_signal_7145) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_7148), .Q (new_AGEMA_signal_7149) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_7152), .Q (new_AGEMA_signal_7153) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_7156), .Q (new_AGEMA_signal_7157) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_7160), .Q (new_AGEMA_signal_7161) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_7164), .Q (new_AGEMA_signal_7165) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_7168), .Q (new_AGEMA_signal_7169) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_7173) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_7176), .Q (new_AGEMA_signal_7177) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_7180), .Q (new_AGEMA_signal_7181) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_7184), .Q (new_AGEMA_signal_7185) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_7188), .Q (new_AGEMA_signal_7189) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_7192), .Q (new_AGEMA_signal_7193) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_7196), .Q (new_AGEMA_signal_7197) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_7200), .Q (new_AGEMA_signal_7201) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_7204), .Q (new_AGEMA_signal_7205) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_7208), .Q (new_AGEMA_signal_7209) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_7212), .Q (new_AGEMA_signal_7213) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_7216), .Q (new_AGEMA_signal_7217) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_7220), .Q (new_AGEMA_signal_7221) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_7224), .Q (new_AGEMA_signal_7225) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_7228), .Q (new_AGEMA_signal_7229) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_7232), .Q (new_AGEMA_signal_7233) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_7236), .Q (new_AGEMA_signal_7237) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_7240), .Q (new_AGEMA_signal_7241) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_7244), .Q (new_AGEMA_signal_7245) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_7248), .Q (new_AGEMA_signal_7249) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_7252), .Q (new_AGEMA_signal_7253) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_7256), .Q (new_AGEMA_signal_7257) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_7260), .Q (new_AGEMA_signal_7261) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_7264), .Q (new_AGEMA_signal_7265) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_7268), .Q (new_AGEMA_signal_7269) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_7272), .Q (new_AGEMA_signal_7273) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_7276), .Q (new_AGEMA_signal_7277) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_7280), .Q (new_AGEMA_signal_7281) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_7284), .Q (new_AGEMA_signal_7285) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_7288), .Q (new_AGEMA_signal_7289) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_7292), .Q (new_AGEMA_signal_7293) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_7296), .Q (new_AGEMA_signal_7297) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_7300), .Q (new_AGEMA_signal_7301) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_7304), .Q (new_AGEMA_signal_7305) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_7308), .Q (new_AGEMA_signal_7309) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_7312), .Q (new_AGEMA_signal_7313) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_7316), .Q (new_AGEMA_signal_7317) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_7320), .Q (new_AGEMA_signal_7321) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_7324), .Q (new_AGEMA_signal_7325) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_7328), .Q (new_AGEMA_signal_7329) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_7332), .Q (new_AGEMA_signal_7333) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_7336), .Q (new_AGEMA_signal_7337) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_7340), .Q (new_AGEMA_signal_7341) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_7344), .Q (new_AGEMA_signal_7345) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_7348), .Q (new_AGEMA_signal_7349) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_7352), .Q (new_AGEMA_signal_7353) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_7356), .Q (new_AGEMA_signal_7357) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_7360), .Q (new_AGEMA_signal_7361) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_7364), .Q (new_AGEMA_signal_7365) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_7368), .Q (new_AGEMA_signal_7369) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_7372), .Q (new_AGEMA_signal_7373) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_7376), .Q (new_AGEMA_signal_7377) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_7380), .Q (new_AGEMA_signal_7381) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_7384), .Q (new_AGEMA_signal_7385) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_7388), .Q (new_AGEMA_signal_7389) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_7392), .Q (new_AGEMA_signal_7393) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_7396), .Q (new_AGEMA_signal_7397) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_7400), .Q (new_AGEMA_signal_7401) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_7404), .Q (new_AGEMA_signal_7405) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_7408), .Q (new_AGEMA_signal_7409) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_7412), .Q (new_AGEMA_signal_7413) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_7416), .Q (new_AGEMA_signal_7417) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_7420), .Q (new_AGEMA_signal_7421) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_7424), .Q (new_AGEMA_signal_7425) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_7428), .Q (new_AGEMA_signal_7429) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_7432), .Q (new_AGEMA_signal_7433) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_7436), .Q (new_AGEMA_signal_7437) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_7440), .Q (new_AGEMA_signal_7441) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_7445) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_7449) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_7453) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_7457) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_7461) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_7465) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_7469) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_7472), .Q (new_AGEMA_signal_7473) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_7477) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_7480), .Q (new_AGEMA_signal_7481) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_7485) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_7489) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_7493) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_7497) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_7501) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_7504), .Q (new_AGEMA_signal_7505) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_7509) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_7512), .Q (new_AGEMA_signal_7513) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_7517) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_7520), .Q (new_AGEMA_signal_7521) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_7524), .Q (new_AGEMA_signal_7525) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_7529) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_7532), .Q (new_AGEMA_signal_7533) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_7537) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_7540), .Q (new_AGEMA_signal_7541) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_7544), .Q (new_AGEMA_signal_7545) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_7548), .Q (new_AGEMA_signal_7549) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_7552), .Q (new_AGEMA_signal_7553) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_7556), .Q (new_AGEMA_signal_7557) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_7560), .Q (new_AGEMA_signal_7561) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_7562) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_7565), .Q (new_AGEMA_signal_7566) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_7569), .Q (new_AGEMA_signal_7570) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_7573), .Q (new_AGEMA_signal_7574) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_7577), .Q (new_AGEMA_signal_7578) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_7581), .Q (new_AGEMA_signal_7582) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_7585), .Q (new_AGEMA_signal_7586) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_7589), .Q (new_AGEMA_signal_7590) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_7593), .Q (new_AGEMA_signal_7594) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_7597), .Q (new_AGEMA_signal_7598) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_7601), .Q (new_AGEMA_signal_7602) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_7605), .Q (new_AGEMA_signal_7606) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_7609), .Q (new_AGEMA_signal_7610) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_7613), .Q (new_AGEMA_signal_7614) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_7617), .Q (new_AGEMA_signal_7618) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_7621), .Q (new_AGEMA_signal_7622) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_7625), .Q (new_AGEMA_signal_7626) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_7629), .Q (new_AGEMA_signal_7630) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_7633), .Q (new_AGEMA_signal_7634) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_7637), .Q (new_AGEMA_signal_7638) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_7641), .Q (new_AGEMA_signal_7642) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_7645), .Q (new_AGEMA_signal_7646) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_7649), .Q (new_AGEMA_signal_7650) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_7653), .Q (new_AGEMA_signal_7654) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_7657), .Q (new_AGEMA_signal_7658) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_7661), .Q (new_AGEMA_signal_7662) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_7665), .Q (new_AGEMA_signal_7666) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_7669), .Q (new_AGEMA_signal_7670) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_7673), .Q (new_AGEMA_signal_7674) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_7677), .Q (new_AGEMA_signal_7678) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_7681), .Q (new_AGEMA_signal_7682) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_7685), .Q (new_AGEMA_signal_7686) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_7689), .Q (new_AGEMA_signal_7690) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_7693), .Q (new_AGEMA_signal_7694) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_7697), .Q (new_AGEMA_signal_7698) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_7701), .Q (new_AGEMA_signal_7702) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_7705), .Q (new_AGEMA_signal_7706) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_7709), .Q (new_AGEMA_signal_7710) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_7713), .Q (new_AGEMA_signal_7714) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_7717), .Q (new_AGEMA_signal_7718) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_7721), .Q (new_AGEMA_signal_7722) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_7725), .Q (new_AGEMA_signal_7726) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_7729), .Q (new_AGEMA_signal_7730) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (clk), .D (new_AGEMA_signal_7733), .Q (new_AGEMA_signal_7734) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_7737), .Q (new_AGEMA_signal_7738) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_7741), .Q (new_AGEMA_signal_7742) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_7745), .Q (new_AGEMA_signal_7746) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_7749), .Q (new_AGEMA_signal_7750) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_7753), .Q (new_AGEMA_signal_7754) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_7757), .Q (new_AGEMA_signal_7758) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_7761), .Q (new_AGEMA_signal_7762) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_7765), .Q (new_AGEMA_signal_7766) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (clk), .D (new_AGEMA_signal_7769), .Q (new_AGEMA_signal_7770) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_7773), .Q (new_AGEMA_signal_7774) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_7777), .Q (new_AGEMA_signal_7778) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_7781), .Q (new_AGEMA_signal_7782) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_7785), .Q (new_AGEMA_signal_7786) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_7789), .Q (new_AGEMA_signal_7790) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_7793), .Q (new_AGEMA_signal_7794) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_7797), .Q (new_AGEMA_signal_7798) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_7801), .Q (new_AGEMA_signal_7802) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (clk), .D (new_AGEMA_signal_7805), .Q (new_AGEMA_signal_7806) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_7809), .Q (new_AGEMA_signal_7810) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_7813), .Q (new_AGEMA_signal_7814) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (clk), .D (new_AGEMA_signal_7817), .Q (new_AGEMA_signal_7818) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_7821), .Q (new_AGEMA_signal_7822) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_7825), .Q (new_AGEMA_signal_7826) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_7829), .Q (new_AGEMA_signal_7830) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_7833), .Q (new_AGEMA_signal_7834) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_7837), .Q (new_AGEMA_signal_7838) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (clk), .D (new_AGEMA_signal_7841), .Q (new_AGEMA_signal_7842) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_7845), .Q (new_AGEMA_signal_7846) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_7849), .Q (new_AGEMA_signal_7850) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (clk), .D (new_AGEMA_signal_7853), .Q (new_AGEMA_signal_7854) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_7857), .Q (new_AGEMA_signal_7858) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_7861), .Q (new_AGEMA_signal_7862) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_7865), .Q (new_AGEMA_signal_7866) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_7869), .Q (new_AGEMA_signal_7870) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (new_AGEMA_signal_7873), .Q (new_AGEMA_signal_7874) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (new_AGEMA_signal_7877), .Q (new_AGEMA_signal_7878) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_7881), .Q (new_AGEMA_signal_7882) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_7885), .Q (new_AGEMA_signal_7886) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_7889), .Q (new_AGEMA_signal_7890) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_7893), .Q (new_AGEMA_signal_7894) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (new_AGEMA_signal_7897), .Q (new_AGEMA_signal_7898) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (clk), .D (new_AGEMA_signal_7901), .Q (new_AGEMA_signal_7902) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_7905), .Q (new_AGEMA_signal_7906) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_7909), .Q (new_AGEMA_signal_7910) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (clk), .D (new_AGEMA_signal_7913), .Q (new_AGEMA_signal_7914) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (new_AGEMA_signal_7917), .Q (new_AGEMA_signal_7918) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (clk), .D (new_AGEMA_signal_7921), .Q (new_AGEMA_signal_7922) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (clk), .D (new_AGEMA_signal_7925), .Q (new_AGEMA_signal_7926) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_7929), .Q (new_AGEMA_signal_7930) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_7933), .Q (new_AGEMA_signal_7934) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (new_AGEMA_signal_7937), .Q (new_AGEMA_signal_7938) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (clk), .D (new_AGEMA_signal_7941), .Q (new_AGEMA_signal_7942) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_7945), .Q (new_AGEMA_signal_7946) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_6793), .Q (new_AGEMA_signal_8091) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_8094), .Q (new_AGEMA_signal_8095) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_8098), .Q (new_AGEMA_signal_8099) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_8102), .Q (new_AGEMA_signal_8103) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_8106), .Q (new_AGEMA_signal_8107) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_1_DQ), .Q (new_AGEMA_signal_8108) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_3674), .Q (new_AGEMA_signal_8109) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_3675), .Q (new_AGEMA_signal_8110) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_3_DQ), .Q (new_AGEMA_signal_8111) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_8112) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_8113) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_5_DQ), .Q (new_AGEMA_signal_8114) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_8115) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_8116) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_7_DQ), .Q (new_AGEMA_signal_8117) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_8118) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_8119) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_9_DQ), .Q (new_AGEMA_signal_8120) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_3686), .Q (new_AGEMA_signal_8121) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_3687), .Q (new_AGEMA_signal_8122) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_11_DQ), .Q (new_AGEMA_signal_8123) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_3690), .Q (new_AGEMA_signal_8124) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_3691), .Q (new_AGEMA_signal_8125) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_13_DQ), .Q (new_AGEMA_signal_8126) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_8127) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_3693), .Q (new_AGEMA_signal_8128) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_15_DQ), .Q (new_AGEMA_signal_8129) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_8130) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_8131) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_17_DQ), .Q (new_AGEMA_signal_8132) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_3698), .Q (new_AGEMA_signal_8133) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_3699), .Q (new_AGEMA_signal_8134) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_19_DQ), .Q (new_AGEMA_signal_8135) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_3702), .Q (new_AGEMA_signal_8136) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_3703), .Q (new_AGEMA_signal_8137) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_21_DQ), .Q (new_AGEMA_signal_8138) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_8139) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_3705), .Q (new_AGEMA_signal_8140) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_23_DQ), .Q (new_AGEMA_signal_8141) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_8142) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_8143) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_25_DQ), .Q (new_AGEMA_signal_8144) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_3710), .Q (new_AGEMA_signal_8145) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C (clk), .D (new_AGEMA_signal_3711), .Q (new_AGEMA_signal_8146) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_27_DQ), .Q (new_AGEMA_signal_8147) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_3714), .Q (new_AGEMA_signal_8148) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_3715), .Q (new_AGEMA_signal_8149) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_29_DQ), .Q (new_AGEMA_signal_8150) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_8151) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_3717), .Q (new_AGEMA_signal_8152) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_31_DQ), .Q (new_AGEMA_signal_8153) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_8154) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_8155) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_33_DQ), .Q (new_AGEMA_signal_8156) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_3722), .Q (new_AGEMA_signal_8157) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_3723), .Q (new_AGEMA_signal_8158) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_35_DQ), .Q (new_AGEMA_signal_8159) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_3726), .Q (new_AGEMA_signal_8160) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_8161) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_37_DQ), .Q (new_AGEMA_signal_8162) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_8163) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_8164) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_39_DQ), .Q (new_AGEMA_signal_8165) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_8166) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_8167) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_41_DQ), .Q (new_AGEMA_signal_8168) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_3734), .Q (new_AGEMA_signal_8169) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_3735), .Q (new_AGEMA_signal_8170) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_43_DQ), .Q (new_AGEMA_signal_8171) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_3738), .Q (new_AGEMA_signal_8172) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_8173) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_45_DQ), .Q (new_AGEMA_signal_8174) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_8175) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_8176) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_47_DQ), .Q (new_AGEMA_signal_8177) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_8178) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_8179) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_49_DQ), .Q (new_AGEMA_signal_8180) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_3746), .Q (new_AGEMA_signal_8181) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_3747), .Q (new_AGEMA_signal_8182) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_51_DQ), .Q (new_AGEMA_signal_8183) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_8184) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_8185) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_53_DQ), .Q (new_AGEMA_signal_8186) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_8187) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_8188) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_55_DQ), .Q (new_AGEMA_signal_8189) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_8190) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_8191) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_57_DQ), .Q (new_AGEMA_signal_8192) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_3758), .Q (new_AGEMA_signal_8193) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C (clk), .D (new_AGEMA_signal_3759), .Q (new_AGEMA_signal_8194) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_59_DQ), .Q (new_AGEMA_signal_8195) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_3762), .Q (new_AGEMA_signal_8196) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_3763), .Q (new_AGEMA_signal_8197) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_61_DQ), .Q (new_AGEMA_signal_8198) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_8199) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_3765), .Q (new_AGEMA_signal_8200) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_63_DQ), .Q (new_AGEMA_signal_8201) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_8202) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_8203) ) ;

    /* register cells */
    DFF_X1 controller_roundCounter_count_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8095), .Q (round_Signal[0]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8099), .Q (round_Signal[1]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8103), .Q (round_Signal[2]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_8107), .Q (round_Signal[3]), .QN () ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, Midori_rounds_roundResult_Reg_SFF_0_DQ}), .Q ({new_AGEMA_signal_1867, new_AGEMA_signal_1866, Midori_rounds_roundReg_out[0]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8110, new_AGEMA_signal_8109, new_AGEMA_signal_8108}), .Q ({new_AGEMA_signal_2673, new_AGEMA_signal_2672, Midori_rounds_roundReg_out[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, Midori_rounds_roundResult_Reg_SFF_2_DQ}), .Q ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, Midori_rounds_roundReg_out[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8113, new_AGEMA_signal_8112, new_AGEMA_signal_8111}), .Q ({new_AGEMA_signal_1869, new_AGEMA_signal_1868, Midori_rounds_roundReg_out[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, Midori_rounds_roundResult_Reg_SFF_4_DQ}), .Q ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, Midori_rounds_roundReg_out[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8116, new_AGEMA_signal_8115, new_AGEMA_signal_8114}), .Q ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, Midori_rounds_roundReg_out[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, Midori_rounds_roundResult_Reg_SFF_6_DQ}), .Q ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, Midori_rounds_roundReg_out[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8119, new_AGEMA_signal_8118, new_AGEMA_signal_8117}), .Q ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, Midori_rounds_roundReg_out[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_8_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, Midori_rounds_roundResult_Reg_SFF_8_DQ}), .Q ({new_AGEMA_signal_1899, new_AGEMA_signal_1898, Midori_rounds_roundReg_out[8]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_9_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8122, new_AGEMA_signal_8121, new_AGEMA_signal_8120}), .Q ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, Midori_rounds_roundReg_out[9]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_10_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, Midori_rounds_roundResult_Reg_SFF_10_DQ}), .Q ({new_AGEMA_signal_1905, new_AGEMA_signal_1904, Midori_rounds_roundReg_out[10]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_11_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8125, new_AGEMA_signal_8124, new_AGEMA_signal_8123}), .Q ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, Midori_rounds_roundReg_out[11]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_12_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, Midori_rounds_roundResult_Reg_SFF_12_DQ}), .Q ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, Midori_rounds_roundReg_out[12]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_13_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8128, new_AGEMA_signal_8127, new_AGEMA_signal_8126}), .Q ({new_AGEMA_signal_2703, new_AGEMA_signal_2702, Midori_rounds_roundReg_out[13]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_14_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, Midori_rounds_roundResult_Reg_SFF_14_DQ}), .Q ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, Midori_rounds_roundReg_out[14]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_15_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8131, new_AGEMA_signal_8130, new_AGEMA_signal_8129}), .Q ({new_AGEMA_signal_1917, new_AGEMA_signal_1916, Midori_rounds_roundReg_out[15]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_16_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, Midori_rounds_roundResult_Reg_SFF_16_DQ}), .Q ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, Midori_rounds_roundReg_out[16]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_17_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8134, new_AGEMA_signal_8133, new_AGEMA_signal_8132}), .Q ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, Midori_rounds_roundReg_out[17]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_18_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, Midori_rounds_roundResult_Reg_SFF_18_DQ}), .Q ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, Midori_rounds_roundReg_out[18]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_19_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8137, new_AGEMA_signal_8136, new_AGEMA_signal_8135}), .Q ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, Midori_rounds_roundReg_out[19]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_20_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, Midori_rounds_roundResult_Reg_SFF_20_DQ}), .Q ({new_AGEMA_signal_1947, new_AGEMA_signal_1946, Midori_rounds_roundReg_out[20]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_21_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8140, new_AGEMA_signal_8139, new_AGEMA_signal_8138}), .Q ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, Midori_rounds_roundReg_out[21]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_22_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, Midori_rounds_roundResult_Reg_SFF_22_DQ}), .Q ({new_AGEMA_signal_1953, new_AGEMA_signal_1952, Midori_rounds_roundReg_out[22]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_23_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8143, new_AGEMA_signal_8142, new_AGEMA_signal_8141}), .Q ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, Midori_rounds_roundReg_out[23]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_24_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, Midori_rounds_roundResult_Reg_SFF_24_DQ}), .Q ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, Midori_rounds_roundReg_out[24]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_25_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8146, new_AGEMA_signal_8145, new_AGEMA_signal_8144}), .Q ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, Midori_rounds_roundReg_out[25]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_26_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, Midori_rounds_roundResult_Reg_SFF_26_DQ}), .Q ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, Midori_rounds_roundReg_out[26]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_27_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8149, new_AGEMA_signal_8148, new_AGEMA_signal_8147}), .Q ({new_AGEMA_signal_1965, new_AGEMA_signal_1964, Midori_rounds_roundReg_out[27]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_28_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, Midori_rounds_roundResult_Reg_SFF_28_DQ}), .Q ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, Midori_rounds_roundReg_out[28]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_29_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8152, new_AGEMA_signal_8151, new_AGEMA_signal_8150}), .Q ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, Midori_rounds_roundReg_out[29]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_30_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, Midori_rounds_roundResult_Reg_SFF_30_DQ}), .Q ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, Midori_rounds_roundReg_out[30]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_31_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8155, new_AGEMA_signal_8154, new_AGEMA_signal_8153}), .Q ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, Midori_rounds_roundReg_out[31]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_32_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, Midori_rounds_roundResult_Reg_SFF_32_DQ}), .Q ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, Midori_rounds_roundReg_out[32]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_33_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8158, new_AGEMA_signal_8157, new_AGEMA_signal_8156}), .Q ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, Midori_rounds_roundReg_out[33]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_34_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, Midori_rounds_roundResult_Reg_SFF_34_DQ}), .Q ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, Midori_rounds_roundReg_out[34]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_35_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8161, new_AGEMA_signal_8160, new_AGEMA_signal_8159}), .Q ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, Midori_rounds_roundReg_out[35]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_36_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, Midori_rounds_roundResult_Reg_SFF_36_DQ}), .Q ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, Midori_rounds_roundReg_out[36]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_37_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8164, new_AGEMA_signal_8163, new_AGEMA_signal_8162}), .Q ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, Midori_rounds_roundReg_out[37]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_38_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, Midori_rounds_roundResult_Reg_SFF_38_DQ}), .Q ({new_AGEMA_signal_2017, new_AGEMA_signal_2016, Midori_rounds_roundReg_out[38]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_39_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8167, new_AGEMA_signal_8166, new_AGEMA_signal_8165}), .Q ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, Midori_rounds_roundReg_out[39]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_40_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, Midori_rounds_roundResult_Reg_SFF_40_DQ}), .Q ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, Midori_rounds_roundReg_out[40]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_41_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8170, new_AGEMA_signal_8169, new_AGEMA_signal_8168}), .Q ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, Midori_rounds_roundReg_out[41]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_42_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, Midori_rounds_roundResult_Reg_SFF_42_DQ}), .Q ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, Midori_rounds_roundReg_out[42]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_43_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8173, new_AGEMA_signal_8172, new_AGEMA_signal_8171}), .Q ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, Midori_rounds_roundReg_out[43]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_44_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, Midori_rounds_roundResult_Reg_SFF_44_DQ}), .Q ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, Midori_rounds_roundReg_out[44]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_45_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8176, new_AGEMA_signal_8175, new_AGEMA_signal_8174}), .Q ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, Midori_rounds_roundReg_out[45]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_46_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, Midori_rounds_roundResult_Reg_SFF_46_DQ}), .Q ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, Midori_rounds_roundReg_out[46]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_47_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8179, new_AGEMA_signal_8178, new_AGEMA_signal_8177}), .Q ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, Midori_rounds_roundReg_out[47]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_48_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, Midori_rounds_roundResult_Reg_SFF_48_DQ}), .Q ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, Midori_rounds_roundReg_out[48]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_49_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8182, new_AGEMA_signal_8181, new_AGEMA_signal_8180}), .Q ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, Midori_rounds_roundReg_out[49]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_50_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, Midori_rounds_roundResult_Reg_SFF_50_DQ}), .Q ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, Midori_rounds_roundReg_out[50]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_51_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8185, new_AGEMA_signal_8184, new_AGEMA_signal_8183}), .Q ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, Midori_rounds_roundReg_out[51]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_52_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, Midori_rounds_roundResult_Reg_SFF_52_DQ}), .Q ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, Midori_rounds_roundReg_out[52]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_53_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8188, new_AGEMA_signal_8187, new_AGEMA_signal_8186}), .Q ({new_AGEMA_signal_2803, new_AGEMA_signal_2802, Midori_rounds_roundReg_out[53]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_54_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, Midori_rounds_roundResult_Reg_SFF_54_DQ}), .Q ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, Midori_rounds_roundReg_out[54]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_55_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8191, new_AGEMA_signal_8190, new_AGEMA_signal_8189}), .Q ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, Midori_rounds_roundReg_out[55]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_56_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, Midori_rounds_roundResult_Reg_SFF_56_DQ}), .Q ({new_AGEMA_signal_2091, new_AGEMA_signal_2090, Midori_rounds_roundReg_out[56]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_57_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8194, new_AGEMA_signal_8193, new_AGEMA_signal_8192}), .Q ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, Midori_rounds_roundReg_out[57]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_58_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Midori_rounds_roundResult_Reg_SFF_58_DQ}), .Q ({new_AGEMA_signal_2097, new_AGEMA_signal_2096, Midori_rounds_roundReg_out[58]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_59_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8197, new_AGEMA_signal_8196, new_AGEMA_signal_8195}), .Q ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, Midori_rounds_roundReg_out[59]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_60_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, Midori_rounds_roundResult_Reg_SFF_60_DQ}), .Q ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, Midori_rounds_roundReg_out[60]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_61_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8200, new_AGEMA_signal_8199, new_AGEMA_signal_8198}), .Q ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, Midori_rounds_roundReg_out[61]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_62_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Midori_rounds_roundResult_Reg_SFF_62_DQ}), .Q ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, Midori_rounds_roundReg_out[62]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_63_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_8203, new_AGEMA_signal_8202, new_AGEMA_signal_8201}), .Q ({new_AGEMA_signal_2109, new_AGEMA_signal_2108, Midori_rounds_roundReg_out[63]}) ) ;
endmodule
