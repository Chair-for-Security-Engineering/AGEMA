/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_BDDcudd_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [706:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;

    /* cells in depth 0 */

    /* cells in depth 1 */
    buf_clk cell_891 ( .C ( clk ), .D ( X_s0[0] ), .Q ( signal_2337 ) ) ;
    buf_clk cell_893 ( .C ( clk ), .D ( X_s1[0] ), .Q ( signal_2339 ) ) ;
    buf_clk cell_895 ( .C ( clk ), .D ( X_s0[5] ), .Q ( signal_2341 ) ) ;
    buf_clk cell_897 ( .C ( clk ), .D ( X_s1[5] ), .Q ( signal_2343 ) ) ;
    buf_clk cell_919 ( .C ( clk ), .D ( X_s0[2] ), .Q ( signal_2365 ) ) ;
    buf_clk cell_923 ( .C ( clk ), .D ( X_s1[2] ), .Q ( signal_2369 ) ) ;
    buf_clk cell_1051 ( .C ( clk ), .D ( X_s0[3] ), .Q ( signal_2497 ) ) ;
    buf_clk cell_1057 ( .C ( clk ), .D ( X_s1[3] ), .Q ( signal_2503 ) ) ;
    buf_clk cell_1131 ( .C ( clk ), .D ( X_s0[6] ), .Q ( signal_2577 ) ) ;
    buf_clk cell_1141 ( .C ( clk ), .D ( X_s1[6] ), .Q ( signal_2587 ) ) ;
    buf_clk cell_1155 ( .C ( clk ), .D ( X_s0[4] ), .Q ( signal_2601 ) ) ;
    buf_clk cell_1167 ( .C ( clk ), .D ( X_s1[4] ), .Q ( signal_2613 ) ) ;
    buf_clk cell_1179 ( .C ( clk ), .D ( X_s0[7] ), .Q ( signal_2625 ) ) ;
    buf_clk cell_1193 ( .C ( clk ), .D ( X_s1[7] ), .Q ( signal_2639 ) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_176 ( .s ({X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_900, signal_192}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_177 ( .s ({X_s1[0], X_s0[0]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_901, signal_193}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_178 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_903, signal_194}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .s ({X_s1[1], X_s0[1]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_904, signal_195}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .s ({X_s1[5], X_s0[5]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_906, signal_196}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .s ({X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_907, signal_197}) ) ;
    buf_clk cell_892 ( .C ( clk ), .D ( signal_2337 ), .Q ( signal_2338 ) ) ;
    buf_clk cell_894 ( .C ( clk ), .D ( signal_2339 ), .Q ( signal_2340 ) ) ;
    buf_clk cell_896 ( .C ( clk ), .D ( signal_2341 ), .Q ( signal_2342 ) ) ;
    buf_clk cell_898 ( .C ( clk ), .D ( signal_2343 ), .Q ( signal_2344 ) ) ;
    buf_clk cell_920 ( .C ( clk ), .D ( signal_2365 ), .Q ( signal_2366 ) ) ;
    buf_clk cell_924 ( .C ( clk ), .D ( signal_2369 ), .Q ( signal_2370 ) ) ;
    buf_clk cell_1052 ( .C ( clk ), .D ( signal_2497 ), .Q ( signal_2498 ) ) ;
    buf_clk cell_1058 ( .C ( clk ), .D ( signal_2503 ), .Q ( signal_2504 ) ) ;
    buf_clk cell_1132 ( .C ( clk ), .D ( signal_2577 ), .Q ( signal_2578 ) ) ;
    buf_clk cell_1142 ( .C ( clk ), .D ( signal_2587 ), .Q ( signal_2588 ) ) ;
    buf_clk cell_1156 ( .C ( clk ), .D ( signal_2601 ), .Q ( signal_2602 ) ) ;
    buf_clk cell_1168 ( .C ( clk ), .D ( signal_2613 ), .Q ( signal_2614 ) ) ;
    buf_clk cell_1180 ( .C ( clk ), .D ( signal_2625 ), .Q ( signal_2626 ) ) ;
    buf_clk cell_1194 ( .C ( clk ), .D ( signal_2639 ), .Q ( signal_2640 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_899 ( .C ( clk ), .D ( signal_2342 ), .Q ( signal_2345 ) ) ;
    buf_clk cell_901 ( .C ( clk ), .D ( signal_2344 ), .Q ( signal_2347 ) ) ;
    buf_clk cell_903 ( .C ( clk ), .D ( signal_194 ), .Q ( signal_2349 ) ) ;
    buf_clk cell_905 ( .C ( clk ), .D ( signal_903 ), .Q ( signal_2351 ) ) ;
    buf_clk cell_907 ( .C ( clk ), .D ( signal_192 ), .Q ( signal_2353 ) ) ;
    buf_clk cell_909 ( .C ( clk ), .D ( signal_900 ), .Q ( signal_2355 ) ) ;
    buf_clk cell_911 ( .C ( clk ), .D ( signal_193 ), .Q ( signal_2357 ) ) ;
    buf_clk cell_913 ( .C ( clk ), .D ( signal_901 ), .Q ( signal_2359 ) ) ;
    buf_clk cell_915 ( .C ( clk ), .D ( signal_195 ), .Q ( signal_2361 ) ) ;
    buf_clk cell_917 ( .C ( clk ), .D ( signal_904 ), .Q ( signal_2363 ) ) ;
    buf_clk cell_921 ( .C ( clk ), .D ( signal_2366 ), .Q ( signal_2367 ) ) ;
    buf_clk cell_925 ( .C ( clk ), .D ( signal_2370 ), .Q ( signal_2371 ) ) ;
    buf_clk cell_927 ( .C ( clk ), .D ( signal_196 ), .Q ( signal_2373 ) ) ;
    buf_clk cell_929 ( .C ( clk ), .D ( signal_906 ), .Q ( signal_2375 ) ) ;
    buf_clk cell_1053 ( .C ( clk ), .D ( signal_2498 ), .Q ( signal_2499 ) ) ;
    buf_clk cell_1059 ( .C ( clk ), .D ( signal_2504 ), .Q ( signal_2505 ) ) ;
    buf_clk cell_1075 ( .C ( clk ), .D ( signal_197 ), .Q ( signal_2521 ) ) ;
    buf_clk cell_1079 ( .C ( clk ), .D ( signal_907 ), .Q ( signal_2525 ) ) ;
    buf_clk cell_1133 ( .C ( clk ), .D ( signal_2578 ), .Q ( signal_2579 ) ) ;
    buf_clk cell_1143 ( .C ( clk ), .D ( signal_2588 ), .Q ( signal_2589 ) ) ;
    buf_clk cell_1157 ( .C ( clk ), .D ( signal_2602 ), .Q ( signal_2603 ) ) ;
    buf_clk cell_1169 ( .C ( clk ), .D ( signal_2614 ), .Q ( signal_2615 ) ) ;
    buf_clk cell_1181 ( .C ( clk ), .D ( signal_2626 ), .Q ( signal_2627 ) ) ;
    buf_clk cell_1195 ( .C ( clk ), .D ( signal_2640 ), .Q ( signal_2641 ) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .s ({signal_2340, signal_2338}), .b ({1'b0, 1'b0}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_908, signal_198}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_183 ( .s ({signal_2340, signal_2338}), .b ({signal_904, signal_195}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_909, signal_199}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .s ({signal_2340, signal_2338}), .b ({signal_903, signal_194}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_910, signal_200}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b1}), .a ({signal_901, signal_193}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_911, signal_201}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .s ({signal_2344, signal_2342}), .b ({signal_903, signal_194}), .a ({signal_900, signal_192}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_912, signal_202}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_187 ( .s ({signal_2340, signal_2338}), .b ({1'b0, 1'b1}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_913, signal_203}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_188 ( .s ({signal_2344, signal_2342}), .b ({signal_901, signal_193}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_914, signal_204}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_189 ( .s ({signal_2344, signal_2342}), .b ({signal_901, signal_193}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_915, signal_205}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_190 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b1}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_916, signal_206}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_191 ( .s ({signal_2344, signal_2342}), .b ({signal_900, signal_192}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_917, signal_207}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_192 ( .s ({signal_2340, signal_2338}), .b ({1'b0, 1'b0}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_918, signal_208}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_193 ( .s ({signal_2344, signal_2342}), .b ({signal_904, signal_195}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[17] ), .c ({signal_919, signal_209}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_194 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b1}), .a ({signal_900, signal_192}), .clk ( clk ), .r ( Fresh[18] ), .c ({signal_920, signal_210}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_195 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b0}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[19] ), .c ({signal_921, signal_211}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_196 ( .s ({signal_2344, signal_2342}), .b ({signal_904, signal_195}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[20] ), .c ({signal_922, signal_212}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_197 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b1}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[21] ), .c ({signal_923, signal_213}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_198 ( .s ({signal_2344, signal_2342}), .b ({signal_900, signal_192}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[22] ), .c ({signal_924, signal_214}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_199 ( .s ({signal_2344, signal_2342}), .b ({signal_901, signal_193}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[23] ), .c ({signal_925, signal_215}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_200 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b0}), .a ({signal_901, signal_193}), .clk ( clk ), .r ( Fresh[24] ), .c ({signal_926, signal_216}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_201 ( .s ({signal_2340, signal_2338}), .b ({signal_904, signal_195}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[25] ), .c ({signal_927, signal_217}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_202 ( .s ({signal_2344, signal_2342}), .b ({signal_900, signal_192}), .a ({signal_901, signal_193}), .clk ( clk ), .r ( Fresh[26] ), .c ({signal_928, signal_218}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_203 ( .s ({signal_2344, signal_2342}), .b ({signal_903, signal_194}), .a ({signal_901, signal_193}), .clk ( clk ), .r ( Fresh[27] ), .c ({signal_929, signal_219}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_204 ( .s ({signal_2344, signal_2342}), .b ({1'b0, 1'b0}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[28] ), .c ({signal_930, signal_220}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_205 ( .s ({signal_2344, signal_2342}), .b ({signal_900, signal_192}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[29] ), .c ({signal_931, signal_221}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_206 ( .s ({signal_2340, signal_2338}), .b ({signal_903, signal_194}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[30] ), .c ({signal_932, signal_222}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_207 ( .s ({signal_2340, signal_2338}), .b ({signal_903, signal_194}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[31] ), .c ({signal_933, signal_223}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_208 ( .s ({signal_2340, signal_2338}), .b ({1'b0, 1'b1}), .a ({signal_904, signal_195}), .clk ( clk ), .r ( Fresh[32] ), .c ({signal_934, signal_224}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_209 ( .s ({signal_2340, signal_2338}), .b ({signal_904, signal_195}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[33] ), .c ({signal_935, signal_225}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_210 ( .s ({signal_2344, signal_2342}), .b ({signal_904, signal_195}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[34] ), .c ({signal_936, signal_226}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_211 ( .s ({signal_2344, signal_2342}), .b ({signal_904, signal_195}), .a ({signal_900, signal_192}), .clk ( clk ), .r ( Fresh[35] ), .c ({signal_937, signal_227}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_212 ( .s ({signal_2344, signal_2342}), .b ({signal_901, signal_193}), .a ({signal_900, signal_192}), .clk ( clk ), .r ( Fresh[36] ), .c ({signal_938, signal_228}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_213 ( .s ({signal_2344, signal_2342}), .b ({signal_900, signal_192}), .a ({signal_903, signal_194}), .clk ( clk ), .r ( Fresh[37] ), .c ({signal_939, signal_229}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_214 ( .s ({signal_2344, signal_2342}), .b ({signal_903, signal_194}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[38] ), .c ({signal_940, signal_230}) ) ;
    buf_clk cell_900 ( .C ( clk ), .D ( signal_2345 ), .Q ( signal_2346 ) ) ;
    buf_clk cell_902 ( .C ( clk ), .D ( signal_2347 ), .Q ( signal_2348 ) ) ;
    buf_clk cell_904 ( .C ( clk ), .D ( signal_2349 ), .Q ( signal_2350 ) ) ;
    buf_clk cell_906 ( .C ( clk ), .D ( signal_2351 ), .Q ( signal_2352 ) ) ;
    buf_clk cell_908 ( .C ( clk ), .D ( signal_2353 ), .Q ( signal_2354 ) ) ;
    buf_clk cell_910 ( .C ( clk ), .D ( signal_2355 ), .Q ( signal_2356 ) ) ;
    buf_clk cell_912 ( .C ( clk ), .D ( signal_2357 ), .Q ( signal_2358 ) ) ;
    buf_clk cell_914 ( .C ( clk ), .D ( signal_2359 ), .Q ( signal_2360 ) ) ;
    buf_clk cell_916 ( .C ( clk ), .D ( signal_2361 ), .Q ( signal_2362 ) ) ;
    buf_clk cell_918 ( .C ( clk ), .D ( signal_2363 ), .Q ( signal_2364 ) ) ;
    buf_clk cell_922 ( .C ( clk ), .D ( signal_2367 ), .Q ( signal_2368 ) ) ;
    buf_clk cell_926 ( .C ( clk ), .D ( signal_2371 ), .Q ( signal_2372 ) ) ;
    buf_clk cell_928 ( .C ( clk ), .D ( signal_2373 ), .Q ( signal_2374 ) ) ;
    buf_clk cell_930 ( .C ( clk ), .D ( signal_2375 ), .Q ( signal_2376 ) ) ;
    buf_clk cell_1054 ( .C ( clk ), .D ( signal_2499 ), .Q ( signal_2500 ) ) ;
    buf_clk cell_1060 ( .C ( clk ), .D ( signal_2505 ), .Q ( signal_2506 ) ) ;
    buf_clk cell_1076 ( .C ( clk ), .D ( signal_2521 ), .Q ( signal_2522 ) ) ;
    buf_clk cell_1080 ( .C ( clk ), .D ( signal_2525 ), .Q ( signal_2526 ) ) ;
    buf_clk cell_1134 ( .C ( clk ), .D ( signal_2579 ), .Q ( signal_2580 ) ) ;
    buf_clk cell_1144 ( .C ( clk ), .D ( signal_2589 ), .Q ( signal_2590 ) ) ;
    buf_clk cell_1158 ( .C ( clk ), .D ( signal_2603 ), .Q ( signal_2604 ) ) ;
    buf_clk cell_1170 ( .C ( clk ), .D ( signal_2615 ), .Q ( signal_2616 ) ) ;
    buf_clk cell_1182 ( .C ( clk ), .D ( signal_2627 ), .Q ( signal_2628 ) ) ;
    buf_clk cell_1196 ( .C ( clk ), .D ( signal_2641 ), .Q ( signal_2642 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_931 ( .C ( clk ), .D ( signal_2368 ), .Q ( signal_2377 ) ) ;
    buf_clk cell_933 ( .C ( clk ), .D ( signal_2372 ), .Q ( signal_2379 ) ) ;
    buf_clk cell_935 ( .C ( clk ), .D ( signal_198 ), .Q ( signal_2381 ) ) ;
    buf_clk cell_937 ( .C ( clk ), .D ( signal_908 ), .Q ( signal_2383 ) ) ;
    buf_clk cell_939 ( .C ( clk ), .D ( signal_203 ), .Q ( signal_2385 ) ) ;
    buf_clk cell_941 ( .C ( clk ), .D ( signal_913 ), .Q ( signal_2387 ) ) ;
    buf_clk cell_943 ( .C ( clk ), .D ( signal_2374 ), .Q ( signal_2389 ) ) ;
    buf_clk cell_945 ( .C ( clk ), .D ( signal_2376 ), .Q ( signal_2391 ) ) ;
    buf_clk cell_947 ( .C ( clk ), .D ( signal_204 ), .Q ( signal_2393 ) ) ;
    buf_clk cell_949 ( .C ( clk ), .D ( signal_914 ), .Q ( signal_2395 ) ) ;
    buf_clk cell_951 ( .C ( clk ), .D ( signal_229 ), .Q ( signal_2397 ) ) ;
    buf_clk cell_953 ( .C ( clk ), .D ( signal_939 ), .Q ( signal_2399 ) ) ;
    buf_clk cell_955 ( .C ( clk ), .D ( signal_215 ), .Q ( signal_2401 ) ) ;
    buf_clk cell_957 ( .C ( clk ), .D ( signal_925 ), .Q ( signal_2403 ) ) ;
    buf_clk cell_959 ( .C ( clk ), .D ( signal_202 ), .Q ( signal_2405 ) ) ;
    buf_clk cell_961 ( .C ( clk ), .D ( signal_912 ), .Q ( signal_2407 ) ) ;
    buf_clk cell_963 ( .C ( clk ), .D ( signal_206 ), .Q ( signal_2409 ) ) ;
    buf_clk cell_965 ( .C ( clk ), .D ( signal_916 ), .Q ( signal_2411 ) ) ;
    buf_clk cell_967 ( .C ( clk ), .D ( signal_199 ), .Q ( signal_2413 ) ) ;
    buf_clk cell_969 ( .C ( clk ), .D ( signal_909 ), .Q ( signal_2415 ) ) ;
    buf_clk cell_971 ( .C ( clk ), .D ( signal_2358 ), .Q ( signal_2417 ) ) ;
    buf_clk cell_973 ( .C ( clk ), .D ( signal_2360 ), .Q ( signal_2419 ) ) ;
    buf_clk cell_975 ( .C ( clk ), .D ( signal_227 ), .Q ( signal_2421 ) ) ;
    buf_clk cell_977 ( .C ( clk ), .D ( signal_937 ), .Q ( signal_2423 ) ) ;
    buf_clk cell_979 ( .C ( clk ), .D ( signal_201 ), .Q ( signal_2425 ) ) ;
    buf_clk cell_981 ( .C ( clk ), .D ( signal_911 ), .Q ( signal_2427 ) ) ;
    buf_clk cell_983 ( .C ( clk ), .D ( signal_216 ), .Q ( signal_2429 ) ) ;
    buf_clk cell_985 ( .C ( clk ), .D ( signal_926 ), .Q ( signal_2431 ) ) ;
    buf_clk cell_987 ( .C ( clk ), .D ( signal_200 ), .Q ( signal_2433 ) ) ;
    buf_clk cell_989 ( .C ( clk ), .D ( signal_910 ), .Q ( signal_2435 ) ) ;
    buf_clk cell_991 ( .C ( clk ), .D ( signal_230 ), .Q ( signal_2437 ) ) ;
    buf_clk cell_993 ( .C ( clk ), .D ( signal_940 ), .Q ( signal_2439 ) ) ;
    buf_clk cell_995 ( .C ( clk ), .D ( signal_219 ), .Q ( signal_2441 ) ) ;
    buf_clk cell_997 ( .C ( clk ), .D ( signal_929 ), .Q ( signal_2443 ) ) ;
    buf_clk cell_999 ( .C ( clk ), .D ( signal_210 ), .Q ( signal_2445 ) ) ;
    buf_clk cell_1001 ( .C ( clk ), .D ( signal_920 ), .Q ( signal_2447 ) ) ;
    buf_clk cell_1003 ( .C ( clk ), .D ( signal_2354 ), .Q ( signal_2449 ) ) ;
    buf_clk cell_1005 ( .C ( clk ), .D ( signal_2356 ), .Q ( signal_2451 ) ) ;
    buf_clk cell_1007 ( .C ( clk ), .D ( signal_223 ), .Q ( signal_2453 ) ) ;
    buf_clk cell_1009 ( .C ( clk ), .D ( signal_933 ), .Q ( signal_2455 ) ) ;
    buf_clk cell_1011 ( .C ( clk ), .D ( signal_209 ), .Q ( signal_2457 ) ) ;
    buf_clk cell_1013 ( .C ( clk ), .D ( signal_919 ), .Q ( signal_2459 ) ) ;
    buf_clk cell_1015 ( .C ( clk ), .D ( signal_217 ), .Q ( signal_2461 ) ) ;
    buf_clk cell_1017 ( .C ( clk ), .D ( signal_927 ), .Q ( signal_2463 ) ) ;
    buf_clk cell_1019 ( .C ( clk ), .D ( signal_226 ), .Q ( signal_2465 ) ) ;
    buf_clk cell_1021 ( .C ( clk ), .D ( signal_936 ), .Q ( signal_2467 ) ) ;
    buf_clk cell_1023 ( .C ( clk ), .D ( signal_228 ), .Q ( signal_2469 ) ) ;
    buf_clk cell_1025 ( .C ( clk ), .D ( signal_938 ), .Q ( signal_2471 ) ) ;
    buf_clk cell_1027 ( .C ( clk ), .D ( signal_207 ), .Q ( signal_2473 ) ) ;
    buf_clk cell_1029 ( .C ( clk ), .D ( signal_917 ), .Q ( signal_2475 ) ) ;
    buf_clk cell_1031 ( .C ( clk ), .D ( signal_214 ), .Q ( signal_2477 ) ) ;
    buf_clk cell_1033 ( .C ( clk ), .D ( signal_924 ), .Q ( signal_2479 ) ) ;
    buf_clk cell_1035 ( .C ( clk ), .D ( signal_212 ), .Q ( signal_2481 ) ) ;
    buf_clk cell_1037 ( .C ( clk ), .D ( signal_922 ), .Q ( signal_2483 ) ) ;
    buf_clk cell_1039 ( .C ( clk ), .D ( signal_208 ), .Q ( signal_2485 ) ) ;
    buf_clk cell_1041 ( .C ( clk ), .D ( signal_918 ), .Q ( signal_2487 ) ) ;
    buf_clk cell_1043 ( .C ( clk ), .D ( signal_220 ), .Q ( signal_2489 ) ) ;
    buf_clk cell_1045 ( .C ( clk ), .D ( signal_930 ), .Q ( signal_2491 ) ) ;
    buf_clk cell_1047 ( .C ( clk ), .D ( signal_222 ), .Q ( signal_2493 ) ) ;
    buf_clk cell_1049 ( .C ( clk ), .D ( signal_932 ), .Q ( signal_2495 ) ) ;
    buf_clk cell_1055 ( .C ( clk ), .D ( signal_2500 ), .Q ( signal_2501 ) ) ;
    buf_clk cell_1061 ( .C ( clk ), .D ( signal_2506 ), .Q ( signal_2507 ) ) ;
    buf_clk cell_1063 ( .C ( clk ), .D ( signal_211 ), .Q ( signal_2509 ) ) ;
    buf_clk cell_1065 ( .C ( clk ), .D ( signal_921 ), .Q ( signal_2511 ) ) ;
    buf_clk cell_1067 ( .C ( clk ), .D ( signal_213 ), .Q ( signal_2513 ) ) ;
    buf_clk cell_1069 ( .C ( clk ), .D ( signal_923 ), .Q ( signal_2515 ) ) ;
    buf_clk cell_1071 ( .C ( clk ), .D ( signal_205 ), .Q ( signal_2517 ) ) ;
    buf_clk cell_1073 ( .C ( clk ), .D ( signal_915 ), .Q ( signal_2519 ) ) ;
    buf_clk cell_1077 ( .C ( clk ), .D ( signal_2522 ), .Q ( signal_2523 ) ) ;
    buf_clk cell_1081 ( .C ( clk ), .D ( signal_2526 ), .Q ( signal_2527 ) ) ;
    buf_clk cell_1083 ( .C ( clk ), .D ( signal_218 ), .Q ( signal_2529 ) ) ;
    buf_clk cell_1085 ( .C ( clk ), .D ( signal_928 ), .Q ( signal_2531 ) ) ;
    buf_clk cell_1087 ( .C ( clk ), .D ( signal_221 ), .Q ( signal_2533 ) ) ;
    buf_clk cell_1089 ( .C ( clk ), .D ( signal_931 ), .Q ( signal_2535 ) ) ;
    buf_clk cell_1135 ( .C ( clk ), .D ( signal_2580 ), .Q ( signal_2581 ) ) ;
    buf_clk cell_1145 ( .C ( clk ), .D ( signal_2590 ), .Q ( signal_2591 ) ) ;
    buf_clk cell_1159 ( .C ( clk ), .D ( signal_2604 ), .Q ( signal_2605 ) ) ;
    buf_clk cell_1171 ( .C ( clk ), .D ( signal_2616 ), .Q ( signal_2617 ) ) ;
    buf_clk cell_1183 ( .C ( clk ), .D ( signal_2628 ), .Q ( signal_2629 ) ) ;
    buf_clk cell_1197 ( .C ( clk ), .D ( signal_2642 ), .Q ( signal_2643 ) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_215 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[39] ), .c ({signal_941, signal_231}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_216 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[40] ), .c ({signal_942, signal_232}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_217 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[41] ), .c ({signal_943, signal_233}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_218 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[42] ), .c ({signal_944, signal_234}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_219 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[43] ), .c ({signal_945, signal_235}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_220 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[44] ), .c ({signal_946, signal_236}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_221 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[45] ), .c ({signal_947, signal_237}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_222 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[46] ), .c ({signal_948, signal_238}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_223 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[47] ), .c ({signal_949, signal_239}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_224 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[48] ), .c ({signal_950, signal_240}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_225 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[49] ), .c ({signal_951, signal_241}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_226 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[50] ), .c ({signal_952, signal_242}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_227 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[51] ), .c ({signal_953, signal_243}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_228 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[52] ), .c ({signal_954, signal_244}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_229 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[53] ), .c ({signal_955, signal_245}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_230 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[54] ), .c ({signal_956, signal_246}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_231 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[55] ), .c ({signal_957, signal_247}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_232 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[56] ), .c ({signal_958, signal_248}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_233 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[57] ), .c ({signal_959, signal_249}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_234 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[58] ), .c ({signal_960, signal_250}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[59] ), .c ({signal_961, signal_251}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[60] ), .c ({signal_962, signal_252}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[61] ), .c ({signal_963, signal_253}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[62] ), .c ({signal_964, signal_254}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[63] ), .c ({signal_965, signal_255}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[64] ), .c ({signal_966, signal_256}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[65] ), .c ({signal_967, signal_257}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[66] ), .c ({signal_968, signal_258}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[67] ), .c ({signal_969, signal_259}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[68] ), .c ({signal_970, signal_260}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[69] ), .c ({signal_971, signal_261}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[70] ), .c ({signal_972, signal_262}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[71] ), .c ({signal_973, signal_263}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[72] ), .c ({signal_974, signal_264}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[73] ), .c ({signal_975, signal_265}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[74] ), .c ({signal_976, signal_266}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[75] ), .c ({signal_977, signal_267}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[76] ), .c ({signal_978, signal_268}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[77] ), .c ({signal_979, signal_269}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[78] ), .c ({signal_980, signal_270}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[79] ), .c ({signal_981, signal_271}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[80] ), .c ({signal_982, signal_272}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_257 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[81] ), .c ({signal_983, signal_273}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[82] ), .c ({signal_984, signal_274}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[83] ), .c ({signal_985, signal_275}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[84] ), .c ({signal_986, signal_276}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[85] ), .c ({signal_987, signal_277}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[86] ), .c ({signal_988, signal_278}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[87] ), .c ({signal_989, signal_279}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[88] ), .c ({signal_990, signal_280}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[89] ), .c ({signal_991, signal_281}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[90] ), .c ({signal_992, signal_282}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_267 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[91] ), .c ({signal_993, signal_283}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_268 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[92] ), .c ({signal_994, signal_284}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[93] ), .c ({signal_995, signal_285}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[94] ), .c ({signal_996, signal_286}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[95] ), .c ({signal_997, signal_287}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[96] ), .c ({signal_998, signal_288}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[97] ), .c ({signal_999, signal_289}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[98] ), .c ({signal_1000, signal_290}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[99] ), .c ({signal_1001, signal_291}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[100] ), .c ({signal_1002, signal_292}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[101] ), .c ({signal_1003, signal_293}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[102] ), .c ({signal_1004, signal_294}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .s ({signal_2372, signal_2368}), .b ({signal_925, signal_215}), .a ({signal_938, signal_228}), .clk ( clk ), .r ( Fresh[103] ), .c ({signal_1006, signal_295}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_280 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[104] ), .c ({signal_1007, signal_296}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_281 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[105] ), .c ({signal_1008, signal_297}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_282 ( .s ({signal_2372, signal_2368}), .b ({signal_918, signal_208}), .a ({signal_914, signal_204}), .clk ( clk ), .r ( Fresh[106] ), .c ({signal_1009, signal_298}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_283 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[107] ), .c ({signal_1010, signal_299}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_284 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[108] ), .c ({signal_1011, signal_300}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_285 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[109] ), .c ({signal_1012, signal_301}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_286 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[110] ), .c ({signal_1013, signal_302}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_287 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[111] ), .c ({signal_1014, signal_303}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_288 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[112] ), .c ({signal_1015, signal_304}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_289 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[113] ), .c ({signal_1016, signal_305}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_290 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[114] ), .c ({signal_1017, signal_306}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_291 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[115] ), .c ({signal_1018, signal_307}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_292 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[116] ), .c ({signal_1019, signal_308}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_293 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[117] ), .c ({signal_1020, signal_309}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_294 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[118] ), .c ({signal_1021, signal_310}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_295 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[119] ), .c ({signal_1022, signal_311}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_296 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[120] ), .c ({signal_1023, signal_312}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_297 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[121] ), .c ({signal_1024, signal_313}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_298 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[122] ), .c ({signal_1025, signal_314}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_299 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[123] ), .c ({signal_1026, signal_315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_300 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[124] ), .c ({signal_1027, signal_316}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_301 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[125] ), .c ({signal_1028, signal_317}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_302 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[126] ), .c ({signal_1029, signal_318}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_303 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[127] ), .c ({signal_1030, signal_319}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_304 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[128] ), .c ({signal_1031, signal_320}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_305 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[129] ), .c ({signal_1032, signal_321}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_306 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[130] ), .c ({signal_1033, signal_322}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_307 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[131] ), .c ({signal_1034, signal_323}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_308 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[132] ), .c ({signal_1035, signal_324}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_309 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[133] ), .c ({signal_1036, signal_325}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_310 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[134] ), .c ({signal_1037, signal_326}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_311 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[135] ), .c ({signal_1038, signal_327}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_312 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[136] ), .c ({signal_1039, signal_328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_313 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[137] ), .c ({signal_1040, signal_329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_314 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[138] ), .c ({signal_1041, signal_330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_315 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[139] ), .c ({signal_1042, signal_331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_316 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[140] ), .c ({signal_1043, signal_332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_317 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[141] ), .c ({signal_1044, signal_333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_318 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[142] ), .c ({signal_1045, signal_334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_319 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[143] ), .c ({signal_1046, signal_335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_320 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[144] ), .c ({signal_1047, signal_336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_321 ( .s ({signal_2372, signal_2368}), .b ({signal_936, signal_226}), .a ({signal_2376, signal_2374}), .clk ( clk ), .r ( Fresh[145] ), .c ({signal_1048, signal_337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_322 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[146] ), .c ({signal_1049, signal_338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_323 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[147] ), .c ({signal_1050, signal_339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_324 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[148] ), .c ({signal_1051, signal_340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_325 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[149] ), .c ({signal_1052, signal_341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_326 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[150] ), .c ({signal_1053, signal_342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_327 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[151] ), .c ({signal_1054, signal_343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_328 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[152] ), .c ({signal_1055, signal_344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_329 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[153] ), .c ({signal_1056, signal_345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_330 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[154] ), .c ({signal_1057, signal_346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_331 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[155] ), .c ({signal_1058, signal_347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_332 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[156] ), .c ({signal_1059, signal_348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_333 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[157] ), .c ({signal_1060, signal_349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_334 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[158] ), .c ({signal_1061, signal_350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_335 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_2352, signal_2350}), .clk ( clk ), .r ( Fresh[159] ), .c ({signal_1062, signal_351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_336 ( .s ({signal_2372, signal_2368}), .b ({signal_933, signal_223}), .a ({signal_937, signal_227}), .clk ( clk ), .r ( Fresh[160] ), .c ({signal_1063, signal_352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_337 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[161] ), .c ({signal_1064, signal_353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_338 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[162] ), .c ({signal_1065, signal_354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_339 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[163] ), .c ({signal_1066, signal_355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_340 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[164] ), .c ({signal_1067, signal_356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_341 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[165] ), .c ({signal_1068, signal_357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_342 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[166] ), .c ({signal_1069, signal_358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_343 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[167] ), .c ({signal_1070, signal_359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_344 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[168] ), .c ({signal_1071, signal_360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_345 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[169] ), .c ({signal_1072, signal_361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_346 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[170] ), .c ({signal_1073, signal_362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_347 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_934, signal_224}), .clk ( clk ), .r ( Fresh[171] ), .c ({signal_1074, signal_363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_348 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[172] ), .c ({signal_1075, signal_364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_349 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[173] ), .c ({signal_1076, signal_365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_350 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[174] ), .c ({signal_1077, signal_366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_351 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[175] ), .c ({signal_1078, signal_367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_352 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[176] ), .c ({signal_1079, signal_368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_353 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[177] ), .c ({signal_1080, signal_369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_354 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[178] ), .c ({signal_1081, signal_370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_355 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[179] ), .c ({signal_1082, signal_371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_356 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[180] ), .c ({signal_1083, signal_372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_357 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[181] ), .c ({signal_1084, signal_373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_358 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[182] ), .c ({signal_1085, signal_374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_359 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[183] ), .c ({signal_1086, signal_375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_360 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[184] ), .c ({signal_1087, signal_376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_361 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[185] ), .c ({signal_1088, signal_377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_362 ( .s ({signal_2348, signal_2346}), .b ({signal_2364, signal_2362}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[186] ), .c ({signal_1089, signal_378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_363 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[187] ), .c ({signal_1090, signal_379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_364 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[188] ), .c ({signal_1091, signal_380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_365 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_2356, signal_2354}), .clk ( clk ), .r ( Fresh[189] ), .c ({signal_1092, signal_381}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_366 ( .s ({signal_2372, signal_2368}), .b ({signal_915, signal_205}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[190] ), .c ({signal_1093, signal_382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_367 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b0}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[191] ), .c ({signal_1094, signal_383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_368 ( .s ({signal_2372, signal_2368}), .b ({signal_918, signal_208}), .a ({signal_2364, signal_2362}), .clk ( clk ), .r ( Fresh[192] ), .c ({signal_1095, signal_384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_369 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[193] ), .c ({signal_1096, signal_385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_370 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[194] ), .c ({signal_1097, signal_386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_371 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[195] ), .c ({signal_1098, signal_387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_372 ( .s ({signal_2348, signal_2346}), .b ({1'b0, 1'b1}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[196] ), .c ({signal_1099, signal_388}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_373 ( .s ({signal_2348, signal_2346}), .b ({signal_927, signal_217}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[197] ), .c ({signal_1100, signal_389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_374 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[198] ), .c ({signal_1101, signal_390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_375 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_909, signal_199}), .clk ( clk ), .r ( Fresh[199] ), .c ({signal_1102, signal_391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_376 ( .s ({signal_2372, signal_2368}), .b ({signal_934, signal_224}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[200] ), .c ({signal_1103, signal_392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_377 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[201] ), .c ({signal_1104, signal_393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_378 ( .s ({signal_2348, signal_2346}), .b ({signal_2356, signal_2354}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[202] ), .c ({signal_1105, signal_394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_379 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[203] ), .c ({signal_1106, signal_395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_380 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[204] ), .c ({signal_1107, signal_396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_381 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({1'b0, 1'b1}), .clk ( clk ), .r ( Fresh[205] ), .c ({signal_1108, signal_397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_382 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[206] ), .c ({signal_1109, signal_398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_383 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[207] ), .c ({signal_1110, signal_399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_384 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[208] ), .c ({signal_1111, signal_400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_385 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[209] ), .c ({signal_1112, signal_401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_386 ( .s ({signal_2348, signal_2346}), .b ({signal_918, signal_208}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[210] ), .c ({signal_1113, signal_402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_387 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_935, signal_225}), .clk ( clk ), .r ( Fresh[211] ), .c ({signal_1114, signal_403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_388 ( .s ({signal_2348, signal_2346}), .b ({signal_932, signal_222}), .a ({1'b0, 1'b0}), .clk ( clk ), .r ( Fresh[212] ), .c ({signal_1115, signal_404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_389 ( .s ({signal_2348, signal_2346}), .b ({signal_934, signal_224}), .a ({signal_933, signal_223}), .clk ( clk ), .r ( Fresh[213] ), .c ({signal_1116, signal_405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_390 ( .s ({signal_2348, signal_2346}), .b ({signal_2360, signal_2358}), .a ({signal_927, signal_217}), .clk ( clk ), .r ( Fresh[214] ), .c ({signal_1117, signal_406}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_391 ( .s ({signal_2348, signal_2346}), .b ({signal_910, signal_200}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[215] ), .c ({signal_1118, signal_407}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_392 ( .s ({signal_2348, signal_2346}), .b ({signal_933, signal_223}), .a ({signal_910, signal_200}), .clk ( clk ), .r ( Fresh[216] ), .c ({signal_1119, signal_408}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_393 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_913, signal_203}), .clk ( clk ), .r ( Fresh[217] ), .c ({signal_1120, signal_409}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_394 ( .s ({signal_2348, signal_2346}), .b ({signal_2352, signal_2350}), .a ({signal_932, signal_222}), .clk ( clk ), .r ( Fresh[218] ), .c ({signal_1121, signal_410}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_395 ( .s ({signal_2348, signal_2346}), .b ({signal_935, signal_225}), .a ({signal_908, signal_198}), .clk ( clk ), .r ( Fresh[219] ), .c ({signal_1122, signal_411}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_396 ( .s ({signal_2348, signal_2346}), .b ({signal_908, signal_198}), .a ({signal_918, signal_208}), .clk ( clk ), .r ( Fresh[220] ), .c ({signal_1123, signal_412}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_397 ( .s ({signal_2372, signal_2368}), .b ({signal_936, signal_226}), .a ({signal_916, signal_206}), .clk ( clk ), .r ( Fresh[221] ), .c ({signal_1124, signal_413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_398 ( .s ({signal_2348, signal_2346}), .b ({signal_909, signal_199}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[222] ), .c ({signal_1125, signal_414}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_399 ( .s ({signal_2348, signal_2346}), .b ({signal_913, signal_203}), .a ({signal_2360, signal_2358}), .clk ( clk ), .r ( Fresh[223] ), .c ({signal_1126, signal_415}) ) ;
    buf_clk cell_932 ( .C ( clk ), .D ( signal_2377 ), .Q ( signal_2378 ) ) ;
    buf_clk cell_934 ( .C ( clk ), .D ( signal_2379 ), .Q ( signal_2380 ) ) ;
    buf_clk cell_936 ( .C ( clk ), .D ( signal_2381 ), .Q ( signal_2382 ) ) ;
    buf_clk cell_938 ( .C ( clk ), .D ( signal_2383 ), .Q ( signal_2384 ) ) ;
    buf_clk cell_940 ( .C ( clk ), .D ( signal_2385 ), .Q ( signal_2386 ) ) ;
    buf_clk cell_942 ( .C ( clk ), .D ( signal_2387 ), .Q ( signal_2388 ) ) ;
    buf_clk cell_944 ( .C ( clk ), .D ( signal_2389 ), .Q ( signal_2390 ) ) ;
    buf_clk cell_946 ( .C ( clk ), .D ( signal_2391 ), .Q ( signal_2392 ) ) ;
    buf_clk cell_948 ( .C ( clk ), .D ( signal_2393 ), .Q ( signal_2394 ) ) ;
    buf_clk cell_950 ( .C ( clk ), .D ( signal_2395 ), .Q ( signal_2396 ) ) ;
    buf_clk cell_952 ( .C ( clk ), .D ( signal_2397 ), .Q ( signal_2398 ) ) ;
    buf_clk cell_954 ( .C ( clk ), .D ( signal_2399 ), .Q ( signal_2400 ) ) ;
    buf_clk cell_956 ( .C ( clk ), .D ( signal_2401 ), .Q ( signal_2402 ) ) ;
    buf_clk cell_958 ( .C ( clk ), .D ( signal_2403 ), .Q ( signal_2404 ) ) ;
    buf_clk cell_960 ( .C ( clk ), .D ( signal_2405 ), .Q ( signal_2406 ) ) ;
    buf_clk cell_962 ( .C ( clk ), .D ( signal_2407 ), .Q ( signal_2408 ) ) ;
    buf_clk cell_964 ( .C ( clk ), .D ( signal_2409 ), .Q ( signal_2410 ) ) ;
    buf_clk cell_966 ( .C ( clk ), .D ( signal_2411 ), .Q ( signal_2412 ) ) ;
    buf_clk cell_968 ( .C ( clk ), .D ( signal_2413 ), .Q ( signal_2414 ) ) ;
    buf_clk cell_970 ( .C ( clk ), .D ( signal_2415 ), .Q ( signal_2416 ) ) ;
    buf_clk cell_972 ( .C ( clk ), .D ( signal_2417 ), .Q ( signal_2418 ) ) ;
    buf_clk cell_974 ( .C ( clk ), .D ( signal_2419 ), .Q ( signal_2420 ) ) ;
    buf_clk cell_976 ( .C ( clk ), .D ( signal_2421 ), .Q ( signal_2422 ) ) ;
    buf_clk cell_978 ( .C ( clk ), .D ( signal_2423 ), .Q ( signal_2424 ) ) ;
    buf_clk cell_980 ( .C ( clk ), .D ( signal_2425 ), .Q ( signal_2426 ) ) ;
    buf_clk cell_982 ( .C ( clk ), .D ( signal_2427 ), .Q ( signal_2428 ) ) ;
    buf_clk cell_984 ( .C ( clk ), .D ( signal_2429 ), .Q ( signal_2430 ) ) ;
    buf_clk cell_986 ( .C ( clk ), .D ( signal_2431 ), .Q ( signal_2432 ) ) ;
    buf_clk cell_988 ( .C ( clk ), .D ( signal_2433 ), .Q ( signal_2434 ) ) ;
    buf_clk cell_990 ( .C ( clk ), .D ( signal_2435 ), .Q ( signal_2436 ) ) ;
    buf_clk cell_992 ( .C ( clk ), .D ( signal_2437 ), .Q ( signal_2438 ) ) ;
    buf_clk cell_994 ( .C ( clk ), .D ( signal_2439 ), .Q ( signal_2440 ) ) ;
    buf_clk cell_996 ( .C ( clk ), .D ( signal_2441 ), .Q ( signal_2442 ) ) ;
    buf_clk cell_998 ( .C ( clk ), .D ( signal_2443 ), .Q ( signal_2444 ) ) ;
    buf_clk cell_1000 ( .C ( clk ), .D ( signal_2445 ), .Q ( signal_2446 ) ) ;
    buf_clk cell_1002 ( .C ( clk ), .D ( signal_2447 ), .Q ( signal_2448 ) ) ;
    buf_clk cell_1004 ( .C ( clk ), .D ( signal_2449 ), .Q ( signal_2450 ) ) ;
    buf_clk cell_1006 ( .C ( clk ), .D ( signal_2451 ), .Q ( signal_2452 ) ) ;
    buf_clk cell_1008 ( .C ( clk ), .D ( signal_2453 ), .Q ( signal_2454 ) ) ;
    buf_clk cell_1010 ( .C ( clk ), .D ( signal_2455 ), .Q ( signal_2456 ) ) ;
    buf_clk cell_1012 ( .C ( clk ), .D ( signal_2457 ), .Q ( signal_2458 ) ) ;
    buf_clk cell_1014 ( .C ( clk ), .D ( signal_2459 ), .Q ( signal_2460 ) ) ;
    buf_clk cell_1016 ( .C ( clk ), .D ( signal_2461 ), .Q ( signal_2462 ) ) ;
    buf_clk cell_1018 ( .C ( clk ), .D ( signal_2463 ), .Q ( signal_2464 ) ) ;
    buf_clk cell_1020 ( .C ( clk ), .D ( signal_2465 ), .Q ( signal_2466 ) ) ;
    buf_clk cell_1022 ( .C ( clk ), .D ( signal_2467 ), .Q ( signal_2468 ) ) ;
    buf_clk cell_1024 ( .C ( clk ), .D ( signal_2469 ), .Q ( signal_2470 ) ) ;
    buf_clk cell_1026 ( .C ( clk ), .D ( signal_2471 ), .Q ( signal_2472 ) ) ;
    buf_clk cell_1028 ( .C ( clk ), .D ( signal_2473 ), .Q ( signal_2474 ) ) ;
    buf_clk cell_1030 ( .C ( clk ), .D ( signal_2475 ), .Q ( signal_2476 ) ) ;
    buf_clk cell_1032 ( .C ( clk ), .D ( signal_2477 ), .Q ( signal_2478 ) ) ;
    buf_clk cell_1034 ( .C ( clk ), .D ( signal_2479 ), .Q ( signal_2480 ) ) ;
    buf_clk cell_1036 ( .C ( clk ), .D ( signal_2481 ), .Q ( signal_2482 ) ) ;
    buf_clk cell_1038 ( .C ( clk ), .D ( signal_2483 ), .Q ( signal_2484 ) ) ;
    buf_clk cell_1040 ( .C ( clk ), .D ( signal_2485 ), .Q ( signal_2486 ) ) ;
    buf_clk cell_1042 ( .C ( clk ), .D ( signal_2487 ), .Q ( signal_2488 ) ) ;
    buf_clk cell_1044 ( .C ( clk ), .D ( signal_2489 ), .Q ( signal_2490 ) ) ;
    buf_clk cell_1046 ( .C ( clk ), .D ( signal_2491 ), .Q ( signal_2492 ) ) ;
    buf_clk cell_1048 ( .C ( clk ), .D ( signal_2493 ), .Q ( signal_2494 ) ) ;
    buf_clk cell_1050 ( .C ( clk ), .D ( signal_2495 ), .Q ( signal_2496 ) ) ;
    buf_clk cell_1056 ( .C ( clk ), .D ( signal_2501 ), .Q ( signal_2502 ) ) ;
    buf_clk cell_1062 ( .C ( clk ), .D ( signal_2507 ), .Q ( signal_2508 ) ) ;
    buf_clk cell_1064 ( .C ( clk ), .D ( signal_2509 ), .Q ( signal_2510 ) ) ;
    buf_clk cell_1066 ( .C ( clk ), .D ( signal_2511 ), .Q ( signal_2512 ) ) ;
    buf_clk cell_1068 ( .C ( clk ), .D ( signal_2513 ), .Q ( signal_2514 ) ) ;
    buf_clk cell_1070 ( .C ( clk ), .D ( signal_2515 ), .Q ( signal_2516 ) ) ;
    buf_clk cell_1072 ( .C ( clk ), .D ( signal_2517 ), .Q ( signal_2518 ) ) ;
    buf_clk cell_1074 ( .C ( clk ), .D ( signal_2519 ), .Q ( signal_2520 ) ) ;
    buf_clk cell_1078 ( .C ( clk ), .D ( signal_2523 ), .Q ( signal_2524 ) ) ;
    buf_clk cell_1082 ( .C ( clk ), .D ( signal_2527 ), .Q ( signal_2528 ) ) ;
    buf_clk cell_1084 ( .C ( clk ), .D ( signal_2529 ), .Q ( signal_2530 ) ) ;
    buf_clk cell_1086 ( .C ( clk ), .D ( signal_2531 ), .Q ( signal_2532 ) ) ;
    buf_clk cell_1088 ( .C ( clk ), .D ( signal_2533 ), .Q ( signal_2534 ) ) ;
    buf_clk cell_1090 ( .C ( clk ), .D ( signal_2535 ), .Q ( signal_2536 ) ) ;
    buf_clk cell_1136 ( .C ( clk ), .D ( signal_2581 ), .Q ( signal_2582 ) ) ;
    buf_clk cell_1146 ( .C ( clk ), .D ( signal_2591 ), .Q ( signal_2592 ) ) ;
    buf_clk cell_1160 ( .C ( clk ), .D ( signal_2605 ), .Q ( signal_2606 ) ) ;
    buf_clk cell_1172 ( .C ( clk ), .D ( signal_2617 ), .Q ( signal_2618 ) ) ;
    buf_clk cell_1184 ( .C ( clk ), .D ( signal_2629 ), .Q ( signal_2630 ) ) ;
    buf_clk cell_1198 ( .C ( clk ), .D ( signal_2643 ), .Q ( signal_2644 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_1091 ( .C ( clk ), .D ( signal_2502 ), .Q ( signal_2537 ) ) ;
    buf_clk cell_1093 ( .C ( clk ), .D ( signal_2508 ), .Q ( signal_2539 ) ) ;
    buf_clk cell_1095 ( .C ( clk ), .D ( signal_413 ), .Q ( signal_2541 ) ) ;
    buf_clk cell_1097 ( .C ( clk ), .D ( signal_1124 ), .Q ( signal_2543 ) ) ;
    buf_clk cell_1099 ( .C ( clk ), .D ( signal_298 ), .Q ( signal_2545 ) ) ;
    buf_clk cell_1101 ( .C ( clk ), .D ( signal_1009 ), .Q ( signal_2547 ) ) ;
    buf_clk cell_1103 ( .C ( clk ), .D ( signal_382 ), .Q ( signal_2549 ) ) ;
    buf_clk cell_1105 ( .C ( clk ), .D ( signal_1093 ), .Q ( signal_2551 ) ) ;
    buf_clk cell_1107 ( .C ( clk ), .D ( signal_2454 ), .Q ( signal_2553 ) ) ;
    buf_clk cell_1109 ( .C ( clk ), .D ( signal_2456 ), .Q ( signal_2555 ) ) ;
    buf_clk cell_1111 ( .C ( clk ), .D ( signal_231 ), .Q ( signal_2557 ) ) ;
    buf_clk cell_1113 ( .C ( clk ), .D ( signal_941 ), .Q ( signal_2559 ) ) ;
    buf_clk cell_1115 ( .C ( clk ), .D ( signal_384 ), .Q ( signal_2561 ) ) ;
    buf_clk cell_1117 ( .C ( clk ), .D ( signal_1095 ), .Q ( signal_2563 ) ) ;
    buf_clk cell_1119 ( .C ( clk ), .D ( signal_321 ), .Q ( signal_2565 ) ) ;
    buf_clk cell_1121 ( .C ( clk ), .D ( signal_1032 ), .Q ( signal_2567 ) ) ;
    buf_clk cell_1123 ( .C ( clk ), .D ( signal_295 ), .Q ( signal_2569 ) ) ;
    buf_clk cell_1125 ( .C ( clk ), .D ( signal_1006 ), .Q ( signal_2571 ) ) ;
    buf_clk cell_1127 ( .C ( clk ), .D ( signal_352 ), .Q ( signal_2573 ) ) ;
    buf_clk cell_1129 ( .C ( clk ), .D ( signal_1063 ), .Q ( signal_2575 ) ) ;
    buf_clk cell_1137 ( .C ( clk ), .D ( signal_2582 ), .Q ( signal_2583 ) ) ;
    buf_clk cell_1147 ( .C ( clk ), .D ( signal_2592 ), .Q ( signal_2593 ) ) ;
    buf_clk cell_1161 ( .C ( clk ), .D ( signal_2606 ), .Q ( signal_2607 ) ) ;
    buf_clk cell_1173 ( .C ( clk ), .D ( signal_2618 ), .Q ( signal_2619 ) ) ;
    buf_clk cell_1185 ( .C ( clk ), .D ( signal_2630 ), .Q ( signal_2631 ) ) ;
    buf_clk cell_1199 ( .C ( clk ), .D ( signal_2644 ), .Q ( signal_2645 ) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_400 ( .s ({signal_2380, signal_2378}), .b ({signal_1026, signal_315}), .a ({signal_963, signal_253}), .clk ( clk ), .r ( Fresh[224] ), .c ({signal_1127, signal_416}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_401 ( .s ({signal_2380, signal_2378}), .b ({signal_1097, signal_386}), .a ({signal_1064, signal_353}), .clk ( clk ), .r ( Fresh[225] ), .c ({signal_1128, signal_417}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_402 ( .s ({signal_2380, signal_2378}), .b ({signal_1123, signal_412}), .a ({signal_1044, signal_333}), .clk ( clk ), .r ( Fresh[226] ), .c ({signal_1129, signal_418}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_403 ( .s ({signal_2380, signal_2378}), .b ({signal_958, signal_248}), .a ({signal_946, signal_236}), .clk ( clk ), .r ( Fresh[227] ), .c ({signal_1130, signal_419}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_404 ( .s ({signal_2380, signal_2378}), .b ({signal_1032, signal_321}), .a ({signal_2384, signal_2382}), .clk ( clk ), .r ( Fresh[228] ), .c ({signal_1131, signal_420}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_405 ( .s ({signal_2380, signal_2378}), .b ({signal_2388, signal_2386}), .a ({signal_1096, signal_385}), .clk ( clk ), .r ( Fresh[229] ), .c ({signal_1132, signal_421}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_406 ( .s ({signal_2380, signal_2378}), .b ({signal_1102, signal_391}), .a ({signal_1053, signal_342}), .clk ( clk ), .r ( Fresh[230] ), .c ({signal_1133, signal_422}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_407 ( .s ({signal_2380, signal_2378}), .b ({signal_1092, signal_381}), .a ({signal_2392, signal_2390}), .clk ( clk ), .r ( Fresh[231] ), .c ({signal_1134, signal_423}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_408 ( .s ({signal_2380, signal_2378}), .b ({signal_1120, signal_409}), .a ({signal_1033, signal_322}), .clk ( clk ), .r ( Fresh[232] ), .c ({signal_1135, signal_424}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_409 ( .s ({signal_2380, signal_2378}), .b ({signal_2396, signal_2394}), .a ({signal_1041, signal_330}), .clk ( clk ), .r ( Fresh[233] ), .c ({signal_1136, signal_425}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_410 ( .s ({signal_2380, signal_2378}), .b ({signal_969, signal_259}), .a ({signal_1109, signal_398}), .clk ( clk ), .r ( Fresh[234] ), .c ({signal_1137, signal_426}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_411 ( .s ({signal_2380, signal_2378}), .b ({signal_2400, signal_2398}), .a ({signal_1067, signal_356}), .clk ( clk ), .r ( Fresh[235] ), .c ({signal_1138, signal_427}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_412 ( .s ({signal_2380, signal_2378}), .b ({signal_2404, signal_2402}), .a ({signal_1119, signal_408}), .clk ( clk ), .r ( Fresh[236] ), .c ({signal_1139, signal_428}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_413 ( .s ({signal_2380, signal_2378}), .b ({signal_965, signal_255}), .a ({signal_1037, signal_326}), .clk ( clk ), .r ( Fresh[237] ), .c ({signal_1140, signal_429}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_414 ( .s ({signal_2380, signal_2378}), .b ({signal_1086, signal_375}), .a ({signal_1004, signal_294}), .clk ( clk ), .r ( Fresh[238] ), .c ({signal_1141, signal_430}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_415 ( .s ({signal_2380, signal_2378}), .b ({signal_1119, signal_408}), .a ({signal_1121, signal_410}), .clk ( clk ), .r ( Fresh[239] ), .c ({signal_1142, signal_431}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_416 ( .s ({signal_2380, signal_2378}), .b ({signal_2408, signal_2406}), .a ({signal_985, signal_275}), .clk ( clk ), .r ( Fresh[240] ), .c ({signal_1143, signal_432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_417 ( .s ({signal_2380, signal_2378}), .b ({signal_948, signal_238}), .a ({signal_1012, signal_301}), .clk ( clk ), .r ( Fresh[241] ), .c ({signal_1144, signal_433}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_418 ( .s ({signal_2380, signal_2378}), .b ({signal_1080, signal_369}), .a ({signal_2392, signal_2390}), .clk ( clk ), .r ( Fresh[242] ), .c ({signal_1145, signal_434}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_419 ( .s ({signal_2380, signal_2378}), .b ({signal_998, signal_288}), .a ({signal_1096, signal_385}), .clk ( clk ), .r ( Fresh[243] ), .c ({signal_1146, signal_435}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_420 ( .s ({signal_2380, signal_2378}), .b ({signal_1068, signal_357}), .a ({signal_2412, signal_2410}), .clk ( clk ), .r ( Fresh[244] ), .c ({signal_1147, signal_436}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_421 ( .s ({signal_2380, signal_2378}), .b ({signal_1096, signal_385}), .a ({signal_1119, signal_408}), .clk ( clk ), .r ( Fresh[245] ), .c ({signal_1148, signal_437}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_422 ( .s ({signal_2380, signal_2378}), .b ({signal_982, signal_272}), .a ({signal_2416, signal_2414}), .clk ( clk ), .r ( Fresh[246] ), .c ({signal_1149, signal_438}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_423 ( .s ({signal_2380, signal_2378}), .b ({signal_957, signal_247}), .a ({signal_979, signal_269}), .clk ( clk ), .r ( Fresh[247] ), .c ({signal_1150, signal_439}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_424 ( .s ({signal_2380, signal_2378}), .b ({signal_1036, signal_325}), .a ({signal_978, signal_268}), .clk ( clk ), .r ( Fresh[248] ), .c ({signal_1151, signal_440}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_425 ( .s ({signal_2380, signal_2378}), .b ({signal_1079, signal_368}), .a ({signal_1059, signal_348}), .clk ( clk ), .r ( Fresh[249] ), .c ({signal_1152, signal_441}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_426 ( .s ({signal_2380, signal_2378}), .b ({signal_1125, signal_414}), .a ({signal_1087, signal_376}), .clk ( clk ), .r ( Fresh[250] ), .c ({signal_1153, signal_442}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_427 ( .s ({signal_2380, signal_2378}), .b ({signal_2420, signal_2418}), .a ({signal_997, signal_287}), .clk ( clk ), .r ( Fresh[251] ), .c ({signal_1154, signal_443}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_428 ( .s ({signal_2380, signal_2378}), .b ({signal_1100, signal_389}), .a ({signal_1003, signal_293}), .clk ( clk ), .r ( Fresh[252] ), .c ({signal_1155, signal_444}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_429 ( .s ({signal_2380, signal_2378}), .b ({signal_1102, signal_391}), .a ({signal_1042, signal_331}), .clk ( clk ), .r ( Fresh[253] ), .c ({signal_1156, signal_445}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_430 ( .s ({signal_2380, signal_2378}), .b ({signal_1007, signal_296}), .a ({signal_2424, signal_2422}), .clk ( clk ), .r ( Fresh[254] ), .c ({signal_1157, signal_446}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_431 ( .s ({signal_2380, signal_2378}), .b ({signal_1118, signal_407}), .a ({signal_1112, signal_401}), .clk ( clk ), .r ( Fresh[255] ), .c ({signal_1158, signal_447}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_432 ( .s ({signal_2380, signal_2378}), .b ({signal_1067, signal_356}), .a ({signal_2428, signal_2426}), .clk ( clk ), .r ( Fresh[256] ), .c ({signal_1159, signal_448}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_433 ( .s ({signal_2380, signal_2378}), .b ({signal_1109, signal_398}), .a ({signal_978, signal_268}), .clk ( clk ), .r ( Fresh[257] ), .c ({signal_1160, signal_449}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_434 ( .s ({signal_2380, signal_2378}), .b ({signal_989, signal_279}), .a ({signal_1092, signal_381}), .clk ( clk ), .r ( Fresh[258] ), .c ({signal_1161, signal_450}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_435 ( .s ({signal_2380, signal_2378}), .b ({signal_1050, signal_339}), .a ({signal_1041, signal_330}), .clk ( clk ), .r ( Fresh[259] ), .c ({signal_1162, signal_451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_436 ( .s ({signal_2380, signal_2378}), .b ({signal_2428, signal_2426}), .a ({signal_1068, signal_357}), .clk ( clk ), .r ( Fresh[260] ), .c ({signal_1163, signal_452}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_437 ( .s ({signal_2380, signal_2378}), .b ({signal_1123, signal_412}), .a ({signal_1003, signal_293}), .clk ( clk ), .r ( Fresh[261] ), .c ({signal_1164, signal_453}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_438 ( .s ({signal_2380, signal_2378}), .b ({signal_1003, signal_293}), .a ({signal_1039, signal_328}), .clk ( clk ), .r ( Fresh[262] ), .c ({signal_1165, signal_454}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_439 ( .s ({signal_2380, signal_2378}), .b ({signal_1076, signal_365}), .a ({signal_1008, signal_297}), .clk ( clk ), .r ( Fresh[263] ), .c ({signal_1166, signal_455}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_440 ( .s ({signal_2380, signal_2378}), .b ({signal_1107, signal_396}), .a ({signal_1088, signal_377}), .clk ( clk ), .r ( Fresh[264] ), .c ({signal_1167, signal_456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_441 ( .s ({signal_2380, signal_2378}), .b ({signal_2384, signal_2382}), .a ({signal_982, signal_272}), .clk ( clk ), .r ( Fresh[265] ), .c ({signal_1168, signal_457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_442 ( .s ({signal_2380, signal_2378}), .b ({signal_1018, signal_307}), .a ({signal_995, signal_285}), .clk ( clk ), .r ( Fresh[266] ), .c ({signal_1169, signal_458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_443 ( .s ({signal_2380, signal_2378}), .b ({signal_1035, signal_324}), .a ({signal_1106, signal_395}), .clk ( clk ), .r ( Fresh[267] ), .c ({signal_1170, signal_459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_444 ( .s ({signal_2380, signal_2378}), .b ({signal_1053, signal_342}), .a ({signal_982, signal_272}), .clk ( clk ), .r ( Fresh[268] ), .c ({signal_1171, signal_460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_445 ( .s ({signal_2380, signal_2378}), .b ({signal_1091, signal_380}), .a ({signal_2432, signal_2430}), .clk ( clk ), .r ( Fresh[269] ), .c ({signal_1172, signal_461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_446 ( .s ({signal_2380, signal_2378}), .b ({signal_968, signal_258}), .a ({signal_961, signal_251}), .clk ( clk ), .r ( Fresh[270] ), .c ({signal_1173, signal_462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_447 ( .s ({signal_2380, signal_2378}), .b ({signal_1105, signal_394}), .a ({signal_1047, signal_336}), .clk ( clk ), .r ( Fresh[271] ), .c ({signal_1174, signal_463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_448 ( .s ({signal_2380, signal_2378}), .b ({1'b0, 1'b1}), .a ({signal_955, signal_245}), .clk ( clk ), .r ( Fresh[272] ), .c ({signal_1175, signal_464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_449 ( .s ({signal_2380, signal_2378}), .b ({signal_964, signal_254}), .a ({signal_1033, signal_322}), .clk ( clk ), .r ( Fresh[273] ), .c ({signal_1176, signal_465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_450 ( .s ({signal_2380, signal_2378}), .b ({signal_955, signal_245}), .a ({signal_1050, signal_339}), .clk ( clk ), .r ( Fresh[274] ), .c ({signal_1177, signal_466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_451 ( .s ({signal_2380, signal_2378}), .b ({signal_953, signal_243}), .a ({signal_1084, signal_373}), .clk ( clk ), .r ( Fresh[275] ), .c ({signal_1178, signal_467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_452 ( .s ({signal_2380, signal_2378}), .b ({signal_2424, signal_2422}), .a ({signal_1038, signal_327}), .clk ( clk ), .r ( Fresh[276] ), .c ({signal_1179, signal_468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_453 ( .s ({signal_2380, signal_2378}), .b ({signal_1039, signal_328}), .a ({signal_947, signal_237}), .clk ( clk ), .r ( Fresh[277] ), .c ({signal_1180, signal_469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_454 ( .s ({signal_2380, signal_2378}), .b ({signal_1073, signal_362}), .a ({signal_2388, signal_2386}), .clk ( clk ), .r ( Fresh[278] ), .c ({signal_1181, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_455 ( .s ({signal_2380, signal_2378}), .b ({signal_1066, signal_355}), .a ({signal_988, signal_278}), .clk ( clk ), .r ( Fresh[279] ), .c ({signal_1182, signal_471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_456 ( .s ({signal_2380, signal_2378}), .b ({signal_1007, signal_296}), .a ({signal_1126, signal_415}), .clk ( clk ), .r ( Fresh[280] ), .c ({signal_1183, signal_472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_457 ( .s ({signal_2380, signal_2378}), .b ({1'b0, 1'b1}), .a ({signal_1071, signal_360}), .clk ( clk ), .r ( Fresh[281] ), .c ({signal_1184, signal_473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_458 ( .s ({signal_2380, signal_2378}), .b ({signal_974, signal_264}), .a ({signal_996, signal_286}), .clk ( clk ), .r ( Fresh[282] ), .c ({signal_1185, signal_474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_459 ( .s ({signal_2380, signal_2378}), .b ({signal_1115, signal_404}), .a ({signal_2436, signal_2434}), .clk ( clk ), .r ( Fresh[283] ), .c ({signal_1186, signal_475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_460 ( .s ({signal_2380, signal_2378}), .b ({signal_1112, signal_401}), .a ({signal_1028, signal_317}), .clk ( clk ), .r ( Fresh[284] ), .c ({signal_1187, signal_476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_461 ( .s ({signal_2380, signal_2378}), .b ({signal_947, signal_237}), .a ({signal_985, signal_275}), .clk ( clk ), .r ( Fresh[285] ), .c ({signal_1188, signal_477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_462 ( .s ({signal_2380, signal_2378}), .b ({signal_986, signal_276}), .a ({signal_1116, signal_405}), .clk ( clk ), .r ( Fresh[286] ), .c ({signal_1189, signal_478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_463 ( .s ({signal_2380, signal_2378}), .b ({signal_1043, signal_332}), .a ({signal_964, signal_254}), .clk ( clk ), .r ( Fresh[287] ), .c ({signal_1190, signal_479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_464 ( .s ({signal_2380, signal_2378}), .b ({signal_1050, signal_339}), .a ({signal_978, signal_268}), .clk ( clk ), .r ( Fresh[288] ), .c ({signal_1191, signal_480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_465 ( .s ({signal_2380, signal_2378}), .b ({signal_1116, signal_405}), .a ({signal_968, signal_258}), .clk ( clk ), .r ( Fresh[289] ), .c ({signal_1192, signal_481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_466 ( .s ({signal_2380, signal_2378}), .b ({signal_1021, signal_310}), .a ({signal_2440, signal_2438}), .clk ( clk ), .r ( Fresh[290] ), .c ({signal_1193, signal_482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_467 ( .s ({signal_2380, signal_2378}), .b ({signal_977, signal_267}), .a ({signal_980, signal_270}), .clk ( clk ), .r ( Fresh[291] ), .c ({signal_1194, signal_483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_468 ( .s ({signal_2380, signal_2378}), .b ({signal_953, signal_243}), .a ({signal_1050, signal_339}), .clk ( clk ), .r ( Fresh[292] ), .c ({signal_1195, signal_484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_469 ( .s ({signal_2380, signal_2378}), .b ({signal_951, signal_241}), .a ({signal_1069, signal_358}), .clk ( clk ), .r ( Fresh[293] ), .c ({signal_1196, signal_485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_470 ( .s ({signal_2380, signal_2378}), .b ({signal_1040, signal_329}), .a ({signal_2444, signal_2442}), .clk ( clk ), .r ( Fresh[294] ), .c ({signal_1197, signal_486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_471 ( .s ({signal_2380, signal_2378}), .b ({signal_1113, signal_402}), .a ({signal_1089, signal_378}), .clk ( clk ), .r ( Fresh[295] ), .c ({signal_1198, signal_487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_472 ( .s ({signal_2380, signal_2378}), .b ({signal_2412, signal_2410}), .a ({signal_1071, signal_360}), .clk ( clk ), .r ( Fresh[296] ), .c ({signal_1199, signal_488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_473 ( .s ({signal_2380, signal_2378}), .b ({signal_1098, signal_387}), .a ({signal_996, signal_286}), .clk ( clk ), .r ( Fresh[297] ), .c ({signal_1200, signal_489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_474 ( .s ({signal_2380, signal_2378}), .b ({signal_944, signal_234}), .a ({signal_1064, signal_353}), .clk ( clk ), .r ( Fresh[298] ), .c ({signal_1201, signal_490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_475 ( .s ({signal_2380, signal_2378}), .b ({signal_1098, signal_387}), .a ({signal_1052, signal_341}), .clk ( clk ), .r ( Fresh[299] ), .c ({signal_1202, signal_491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_476 ( .s ({signal_2380, signal_2378}), .b ({signal_1109, signal_398}), .a ({signal_2448, signal_2446}), .clk ( clk ), .r ( Fresh[300] ), .c ({signal_1203, signal_492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_477 ( .s ({signal_2380, signal_2378}), .b ({signal_1022, signal_311}), .a ({signal_1077, signal_366}), .clk ( clk ), .r ( Fresh[301] ), .c ({signal_1204, signal_493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_478 ( .s ({signal_2380, signal_2378}), .b ({signal_960, signal_250}), .a ({signal_1114, signal_403}), .clk ( clk ), .r ( Fresh[302] ), .c ({signal_1205, signal_494}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_479 ( .s ({signal_2380, signal_2378}), .b ({signal_1057, signal_346}), .a ({signal_1041, signal_330}), .clk ( clk ), .r ( Fresh[303] ), .c ({signal_1206, signal_495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_480 ( .s ({signal_2380, signal_2378}), .b ({signal_1002, signal_292}), .a ({signal_978, signal_268}), .clk ( clk ), .r ( Fresh[304] ), .c ({signal_1207, signal_496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_481 ( .s ({signal_2380, signal_2378}), .b ({signal_1087, signal_376}), .a ({signal_1028, signal_317}), .clk ( clk ), .r ( Fresh[305] ), .c ({signal_1208, signal_497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_482 ( .s ({signal_2380, signal_2378}), .b ({signal_1098, signal_387}), .a ({signal_984, signal_274}), .clk ( clk ), .r ( Fresh[306] ), .c ({signal_1209, signal_498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_483 ( .s ({signal_2380, signal_2378}), .b ({signal_1031, signal_320}), .a ({signal_1030, signal_319}), .clk ( clk ), .r ( Fresh[307] ), .c ({signal_1210, signal_499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_484 ( .s ({signal_2380, signal_2378}), .b ({signal_1041, signal_330}), .a ({signal_988, signal_278}), .clk ( clk ), .r ( Fresh[308] ), .c ({signal_1211, signal_500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_485 ( .s ({signal_2380, signal_2378}), .b ({signal_1092, signal_381}), .a ({signal_1111, signal_400}), .clk ( clk ), .r ( Fresh[309] ), .c ({signal_1212, signal_501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_486 ( .s ({signal_2380, signal_2378}), .b ({signal_950, signal_240}), .a ({signal_1052, signal_341}), .clk ( clk ), .r ( Fresh[310] ), .c ({signal_1213, signal_502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_487 ( .s ({signal_2380, signal_2378}), .b ({signal_1015, signal_304}), .a ({signal_996, signal_286}), .clk ( clk ), .r ( Fresh[311] ), .c ({signal_1214, signal_503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_488 ( .s ({signal_2380, signal_2378}), .b ({signal_1072, signal_361}), .a ({signal_1071, signal_360}), .clk ( clk ), .r ( Fresh[312] ), .c ({signal_1215, signal_504}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_489 ( .s ({signal_2380, signal_2378}), .b ({signal_970, signal_260}), .a ({signal_977, signal_267}), .clk ( clk ), .r ( Fresh[313] ), .c ({signal_1216, signal_505}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_490 ( .s ({signal_2380, signal_2378}), .b ({signal_1115, signal_404}), .a ({signal_1117, signal_406}), .clk ( clk ), .r ( Fresh[314] ), .c ({signal_1217, signal_506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_491 ( .s ({signal_2380, signal_2378}), .b ({signal_1056, signal_345}), .a ({signal_1061, signal_350}), .clk ( clk ), .r ( Fresh[315] ), .c ({signal_1218, signal_507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_492 ( .s ({signal_2380, signal_2378}), .b ({signal_1091, signal_380}), .a ({signal_955, signal_245}), .clk ( clk ), .r ( Fresh[316] ), .c ({signal_1219, signal_508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_493 ( .s ({signal_2380, signal_2378}), .b ({signal_2452, signal_2450}), .a ({signal_1099, signal_388}), .clk ( clk ), .r ( Fresh[317] ), .c ({signal_1220, signal_509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_494 ( .s ({signal_2380, signal_2378}), .b ({signal_954, signal_244}), .a ({signal_1053, signal_342}), .clk ( clk ), .r ( Fresh[318] ), .c ({signal_1221, signal_510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_495 ( .s ({signal_2380, signal_2378}), .b ({signal_1010, signal_299}), .a ({signal_1115, signal_404}), .clk ( clk ), .r ( Fresh[319] ), .c ({signal_1222, signal_511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_496 ( .s ({signal_2380, signal_2378}), .b ({signal_1044, signal_333}), .a ({signal_960, signal_250}), .clk ( clk ), .r ( Fresh[320] ), .c ({signal_1223, signal_512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_497 ( .s ({signal_2380, signal_2378}), .b ({signal_982, signal_272}), .a ({signal_974, signal_264}), .clk ( clk ), .r ( Fresh[321] ), .c ({signal_1224, signal_513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_498 ( .s ({signal_2380, signal_2378}), .b ({signal_942, signal_232}), .a ({signal_1039, signal_328}), .clk ( clk ), .r ( Fresh[322] ), .c ({signal_1225, signal_514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_499 ( .s ({signal_2380, signal_2378}), .b ({signal_2456, signal_2454}), .a ({signal_1012, signal_301}), .clk ( clk ), .r ( Fresh[323] ), .c ({signal_1226, signal_515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_500 ( .s ({signal_2380, signal_2378}), .b ({signal_1055, signal_344}), .a ({signal_1083, signal_372}), .clk ( clk ), .r ( Fresh[324] ), .c ({signal_1227, signal_516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_501 ( .s ({signal_2380, signal_2378}), .b ({signal_1030, signal_319}), .a ({signal_956, signal_246}), .clk ( clk ), .r ( Fresh[325] ), .c ({signal_1228, signal_517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_502 ( .s ({signal_2380, signal_2378}), .b ({signal_1057, signal_346}), .a ({signal_943, signal_233}), .clk ( clk ), .r ( Fresh[326] ), .c ({signal_1229, signal_518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_503 ( .s ({signal_2380, signal_2378}), .b ({signal_1049, signal_338}), .a ({signal_1104, signal_393}), .clk ( clk ), .r ( Fresh[327] ), .c ({signal_1230, signal_519}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_504 ( .s ({signal_2380, signal_2378}), .b ({signal_1001, signal_291}), .a ({signal_1076, signal_365}), .clk ( clk ), .r ( Fresh[328] ), .c ({signal_1231, signal_520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_505 ( .s ({signal_2380, signal_2378}), .b ({signal_958, signal_248}), .a ({signal_2460, signal_2458}), .clk ( clk ), .r ( Fresh[329] ), .c ({signal_1232, signal_521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_506 ( .s ({signal_2380, signal_2378}), .b ({signal_1065, signal_354}), .a ({signal_1111, signal_400}), .clk ( clk ), .r ( Fresh[330] ), .c ({signal_1233, signal_522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_507 ( .s ({signal_2380, signal_2378}), .b ({signal_2464, signal_2462}), .a ({signal_953, signal_243}), .clk ( clk ), .r ( Fresh[331] ), .c ({signal_1234, signal_523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_508 ( .s ({signal_2380, signal_2378}), .b ({signal_983, signal_273}), .a ({signal_1020, signal_309}), .clk ( clk ), .r ( Fresh[332] ), .c ({signal_1235, signal_524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_509 ( .s ({signal_2380, signal_2378}), .b ({signal_949, signal_239}), .a ({signal_1041, signal_330}), .clk ( clk ), .r ( Fresh[333] ), .c ({signal_1236, signal_525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_510 ( .s ({signal_2380, signal_2378}), .b ({signal_1119, signal_408}), .a ({signal_2408, signal_2406}), .clk ( clk ), .r ( Fresh[334] ), .c ({signal_1237, signal_526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_511 ( .s ({signal_2380, signal_2378}), .b ({signal_1035, signal_324}), .a ({signal_1058, signal_347}), .clk ( clk ), .r ( Fresh[335] ), .c ({signal_1238, signal_527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_512 ( .s ({signal_2380, signal_2378}), .b ({signal_945, signal_235}), .a ({signal_1083, signal_372}), .clk ( clk ), .r ( Fresh[336] ), .c ({signal_1239, signal_528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_513 ( .s ({signal_2380, signal_2378}), .b ({signal_999, signal_289}), .a ({signal_1085, signal_374}), .clk ( clk ), .r ( Fresh[337] ), .c ({signal_1240, signal_529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_514 ( .s ({signal_2380, signal_2378}), .b ({signal_1013, signal_302}), .a ({signal_1061, signal_350}), .clk ( clk ), .r ( Fresh[338] ), .c ({signal_1241, signal_530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_515 ( .s ({signal_2380, signal_2378}), .b ({signal_1037, signal_326}), .a ({signal_1021, signal_310}), .clk ( clk ), .r ( Fresh[339] ), .c ({signal_1242, signal_531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_516 ( .s ({signal_2380, signal_2378}), .b ({signal_1049, signal_338}), .a ({signal_1037, signal_326}), .clk ( clk ), .r ( Fresh[340] ), .c ({signal_1243, signal_532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_517 ( .s ({signal_2380, signal_2378}), .b ({signal_957, signal_247}), .a ({signal_941, signal_231}), .clk ( clk ), .r ( Fresh[341] ), .c ({signal_1244, signal_533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_518 ( .s ({signal_2380, signal_2378}), .b ({signal_1067, signal_356}), .a ({signal_1120, signal_409}), .clk ( clk ), .r ( Fresh[342] ), .c ({signal_1245, signal_534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_519 ( .s ({signal_2380, signal_2378}), .b ({signal_959, signal_249}), .a ({signal_2384, signal_2382}), .clk ( clk ), .r ( Fresh[343] ), .c ({signal_1246, signal_535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_520 ( .s ({signal_2380, signal_2378}), .b ({1'b0, 1'b0}), .a ({signal_1016, signal_305}), .clk ( clk ), .r ( Fresh[344] ), .c ({signal_1247, signal_536}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_521 ( .s ({signal_2380, signal_2378}), .b ({signal_2468, signal_2466}), .a ({signal_1020, signal_309}), .clk ( clk ), .r ( Fresh[345] ), .c ({signal_1248, signal_537}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_522 ( .s ({signal_2380, signal_2378}), .b ({signal_1035, signal_324}), .a ({signal_2456, signal_2454}), .clk ( clk ), .r ( Fresh[346] ), .c ({signal_1249, signal_538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_523 ( .s ({signal_2380, signal_2378}), .b ({signal_2440, signal_2438}), .a ({signal_1062, signal_351}), .clk ( clk ), .r ( Fresh[347] ), .c ({signal_1250, signal_539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_524 ( .s ({signal_2380, signal_2378}), .b ({signal_985, signal_275}), .a ({signal_2392, signal_2390}), .clk ( clk ), .r ( Fresh[348] ), .c ({signal_1251, signal_540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_525 ( .s ({signal_2380, signal_2378}), .b ({signal_966, signal_256}), .a ({signal_985, signal_275}), .clk ( clk ), .r ( Fresh[349] ), .c ({signal_1252, signal_541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_526 ( .s ({signal_2380, signal_2378}), .b ({signal_1037, signal_326}), .a ({signal_1017, signal_306}), .clk ( clk ), .r ( Fresh[350] ), .c ({signal_1253, signal_542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_527 ( .s ({signal_2380, signal_2378}), .b ({signal_1068, signal_357}), .a ({signal_947, signal_237}), .clk ( clk ), .r ( Fresh[351] ), .c ({signal_1254, signal_543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_528 ( .s ({signal_2380, signal_2378}), .b ({signal_1019, signal_308}), .a ({signal_1036, signal_325}), .clk ( clk ), .r ( Fresh[352] ), .c ({signal_1255, signal_544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_529 ( .s ({signal_2380, signal_2378}), .b ({signal_998, signal_288}), .a ({signal_988, signal_278}), .clk ( clk ), .r ( Fresh[353] ), .c ({signal_1256, signal_545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_530 ( .s ({signal_2380, signal_2378}), .b ({signal_1088, signal_377}), .a ({signal_1064, signal_353}), .clk ( clk ), .r ( Fresh[354] ), .c ({signal_1257, signal_546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_531 ( .s ({signal_2380, signal_2378}), .b ({signal_1027, signal_316}), .a ({signal_1074, signal_363}), .clk ( clk ), .r ( Fresh[355] ), .c ({signal_1258, signal_547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_532 ( .s ({signal_2380, signal_2378}), .b ({signal_1100, signal_389}), .a ({signal_1060, signal_349}), .clk ( clk ), .r ( Fresh[356] ), .c ({signal_1259, signal_548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_533 ( .s ({signal_2380, signal_2378}), .b ({signal_1004, signal_294}), .a ({signal_2460, signal_2458}), .clk ( clk ), .r ( Fresh[357] ), .c ({signal_1260, signal_549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_534 ( .s ({signal_2380, signal_2378}), .b ({signal_1091, signal_380}), .a ({signal_1053, signal_342}), .clk ( clk ), .r ( Fresh[358] ), .c ({signal_1261, signal_550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_535 ( .s ({signal_2380, signal_2378}), .b ({signal_1110, signal_399}), .a ({signal_2472, signal_2470}), .clk ( clk ), .r ( Fresh[359] ), .c ({signal_1262, signal_551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_536 ( .s ({signal_2380, signal_2378}), .b ({signal_995, signal_285}), .a ({signal_2436, signal_2434}), .clk ( clk ), .r ( Fresh[360] ), .c ({signal_1263, signal_552}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_537 ( .s ({signal_2380, signal_2378}), .b ({signal_1014, signal_303}), .a ({signal_1015, signal_304}), .clk ( clk ), .r ( Fresh[361] ), .c ({signal_1264, signal_553}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_538 ( .s ({signal_2380, signal_2378}), .b ({signal_1047, signal_336}), .a ({signal_1065, signal_354}), .clk ( clk ), .r ( Fresh[362] ), .c ({signal_1265, signal_554}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_539 ( .s ({signal_2380, signal_2378}), .b ({signal_951, signal_241}), .a ({signal_1084, signal_373}), .clk ( clk ), .r ( Fresh[363] ), .c ({signal_1266, signal_555}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_540 ( .s ({signal_2380, signal_2378}), .b ({signal_1092, signal_381}), .a ({signal_1066, signal_355}), .clk ( clk ), .r ( Fresh[364] ), .c ({signal_1267, signal_556}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_541 ( .s ({signal_2380, signal_2378}), .b ({signal_2476, signal_2474}), .a ({signal_1029, signal_318}), .clk ( clk ), .r ( Fresh[365] ), .c ({signal_1268, signal_557}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_542 ( .s ({signal_2380, signal_2378}), .b ({signal_994, signal_284}), .a ({signal_1021, signal_310}), .clk ( clk ), .r ( Fresh[366] ), .c ({signal_1269, signal_558}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_543 ( .s ({signal_2380, signal_2378}), .b ({signal_1013, signal_302}), .a ({signal_1027, signal_316}), .clk ( clk ), .r ( Fresh[367] ), .c ({signal_1270, signal_559}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_544 ( .s ({signal_2380, signal_2378}), .b ({signal_952, signal_242}), .a ({signal_962, signal_252}), .clk ( clk ), .r ( Fresh[368] ), .c ({signal_1271, signal_560}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_545 ( .s ({signal_2380, signal_2378}), .b ({signal_1060, signal_349}), .a ({signal_1121, signal_410}), .clk ( clk ), .r ( Fresh[369] ), .c ({signal_1272, signal_561}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_546 ( .s ({signal_2380, signal_2378}), .b ({signal_1102, signal_391}), .a ({signal_1115, signal_404}), .clk ( clk ), .r ( Fresh[370] ), .c ({signal_1273, signal_562}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_547 ( .s ({signal_2380, signal_2378}), .b ({signal_1081, signal_370}), .a ({signal_1015, signal_304}), .clk ( clk ), .r ( Fresh[371] ), .c ({signal_1274, signal_563}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_548 ( .s ({signal_2380, signal_2378}), .b ({signal_1045, signal_334}), .a ({signal_1108, signal_397}), .clk ( clk ), .r ( Fresh[372] ), .c ({signal_1275, signal_564}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_549 ( .s ({signal_2380, signal_2378}), .b ({signal_984, signal_274}), .a ({signal_1092, signal_381}), .clk ( clk ), .r ( Fresh[373] ), .c ({signal_1276, signal_565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_550 ( .s ({signal_2380, signal_2378}), .b ({signal_1037, signal_326}), .a ({signal_1024, signal_313}), .clk ( clk ), .r ( Fresh[374] ), .c ({signal_1277, signal_566}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_551 ( .s ({signal_2380, signal_2378}), .b ({signal_1056, signal_345}), .a ({signal_1062, signal_351}), .clk ( clk ), .r ( Fresh[375] ), .c ({signal_1278, signal_567}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_552 ( .s ({signal_2380, signal_2378}), .b ({signal_1000, signal_290}), .a ({signal_948, signal_238}), .clk ( clk ), .r ( Fresh[376] ), .c ({signal_1279, signal_568}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_553 ( .s ({signal_2380, signal_2378}), .b ({signal_1105, signal_394}), .a ({signal_975, signal_265}), .clk ( clk ), .r ( Fresh[377] ), .c ({signal_1280, signal_569}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_554 ( .s ({signal_2380, signal_2378}), .b ({signal_1066, signal_355}), .a ({signal_971, signal_261}), .clk ( clk ), .r ( Fresh[378] ), .c ({signal_1281, signal_570}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_555 ( .s ({signal_2380, signal_2378}), .b ({signal_994, signal_284}), .a ({signal_2480, signal_2478}), .clk ( clk ), .r ( Fresh[379] ), .c ({signal_1282, signal_571}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_556 ( .s ({signal_2380, signal_2378}), .b ({signal_1073, signal_362}), .a ({signal_1003, signal_293}), .clk ( clk ), .r ( Fresh[380] ), .c ({signal_1283, signal_572}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_557 ( .s ({signal_2380, signal_2378}), .b ({signal_1062, signal_351}), .a ({signal_2484, signal_2482}), .clk ( clk ), .r ( Fresh[381] ), .c ({signal_1284, signal_573}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_558 ( .s ({signal_2380, signal_2378}), .b ({signal_954, signal_244}), .a ({signal_980, signal_270}), .clk ( clk ), .r ( Fresh[382] ), .c ({signal_1285, signal_574}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_559 ( .s ({signal_2380, signal_2378}), .b ({signal_1041, signal_330}), .a ({signal_2488, signal_2486}), .clk ( clk ), .r ( Fresh[383] ), .c ({signal_1286, signal_575}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_560 ( .s ({signal_2380, signal_2378}), .b ({signal_999, signal_289}), .a ({signal_976, signal_266}), .clk ( clk ), .r ( Fresh[384] ), .c ({signal_1287, signal_576}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_561 ( .s ({signal_2380, signal_2378}), .b ({signal_1097, signal_386}), .a ({signal_1011, signal_300}), .clk ( clk ), .r ( Fresh[385] ), .c ({signal_1288, signal_577}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_562 ( .s ({signal_2380, signal_2378}), .b ({signal_2492, signal_2490}), .a ({signal_1108, signal_397}), .clk ( clk ), .r ( Fresh[386] ), .c ({signal_1289, signal_578}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_563 ( .s ({signal_2380, signal_2378}), .b ({signal_1094, signal_383}), .a ({signal_1083, signal_372}), .clk ( clk ), .r ( Fresh[387] ), .c ({signal_1290, signal_579}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_564 ( .s ({signal_2380, signal_2378}), .b ({signal_965, signal_255}), .a ({signal_2488, signal_2486}), .clk ( clk ), .r ( Fresh[388] ), .c ({signal_1291, signal_580}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_565 ( .s ({signal_2380, signal_2378}), .b ({signal_989, signal_279}), .a ({signal_1086, signal_375}), .clk ( clk ), .r ( Fresh[389] ), .c ({signal_1292, signal_581}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_566 ( .s ({signal_2380, signal_2378}), .b ({signal_2452, signal_2450}), .a ({signal_1030, signal_319}), .clk ( clk ), .r ( Fresh[390] ), .c ({signal_1293, signal_582}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_567 ( .s ({signal_2380, signal_2378}), .b ({signal_1076, signal_365}), .a ({signal_1028, signal_317}), .clk ( clk ), .r ( Fresh[391] ), .c ({signal_1294, signal_583}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_568 ( .s ({signal_2380, signal_2378}), .b ({signal_1047, signal_336}), .a ({signal_1087, signal_376}), .clk ( clk ), .r ( Fresh[392] ), .c ({signal_1295, signal_584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_569 ( .s ({signal_2380, signal_2378}), .b ({signal_1120, signal_409}), .a ({signal_1042, signal_331}), .clk ( clk ), .r ( Fresh[393] ), .c ({signal_1296, signal_585}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_570 ( .s ({signal_2380, signal_2378}), .b ({signal_951, signal_241}), .a ({signal_973, signal_263}), .clk ( clk ), .r ( Fresh[394] ), .c ({signal_1297, signal_586}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_571 ( .s ({signal_2380, signal_2378}), .b ({signal_979, signal_269}), .a ({signal_1061, signal_350}), .clk ( clk ), .r ( Fresh[395] ), .c ({signal_1298, signal_587}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_572 ( .s ({signal_2380, signal_2378}), .b ({signal_1049, signal_338}), .a ({signal_1085, signal_374}), .clk ( clk ), .r ( Fresh[396] ), .c ({signal_1299, signal_588}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_573 ( .s ({signal_2380, signal_2378}), .b ({signal_1045, signal_334}), .a ({signal_963, signal_253}), .clk ( clk ), .r ( Fresh[397] ), .c ({signal_1300, signal_589}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_574 ( .s ({signal_2380, signal_2378}), .b ({signal_1118, signal_407}), .a ({signal_1081, signal_370}), .clk ( clk ), .r ( Fresh[398] ), .c ({signal_1301, signal_590}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_575 ( .s ({signal_2380, signal_2378}), .b ({signal_997, signal_287}), .a ({signal_992, signal_282}), .clk ( clk ), .r ( Fresh[399] ), .c ({signal_1302, signal_591}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_576 ( .s ({signal_2380, signal_2378}), .b ({signal_2448, signal_2446}), .a ({signal_1050, signal_339}), .clk ( clk ), .r ( Fresh[400] ), .c ({signal_1303, signal_592}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_577 ( .s ({signal_2380, signal_2378}), .b ({signal_1117, signal_406}), .a ({signal_987, signal_277}), .clk ( clk ), .r ( Fresh[401] ), .c ({signal_1304, signal_593}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_578 ( .s ({signal_2380, signal_2378}), .b ({signal_1101, signal_390}), .a ({signal_1061, signal_350}), .clk ( clk ), .r ( Fresh[402] ), .c ({signal_1305, signal_594}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_579 ( .s ({signal_2380, signal_2378}), .b ({signal_1046, signal_335}), .a ({signal_1059, signal_348}), .clk ( clk ), .r ( Fresh[403] ), .c ({signal_1306, signal_595}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_580 ( .s ({signal_2380, signal_2378}), .b ({signal_972, signal_262}), .a ({signal_2428, signal_2426}), .clk ( clk ), .r ( Fresh[404] ), .c ({signal_1307, signal_596}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_581 ( .s ({signal_2380, signal_2378}), .b ({signal_2424, signal_2422}), .a ({signal_1031, signal_320}), .clk ( clk ), .r ( Fresh[405] ), .c ({signal_1308, signal_597}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_582 ( .s ({signal_2380, signal_2378}), .b ({signal_1070, signal_359}), .a ({signal_2496, signal_2494}), .clk ( clk ), .r ( Fresh[406] ), .c ({signal_1309, signal_598}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_583 ( .s ({signal_2380, signal_2378}), .b ({signal_1107, signal_396}), .a ({signal_1037, signal_326}), .clk ( clk ), .r ( Fresh[407] ), .c ({signal_1310, signal_599}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_584 ( .s ({signal_2380, signal_2378}), .b ({signal_1024, signal_313}), .a ({signal_1062, signal_351}), .clk ( clk ), .r ( Fresh[408] ), .c ({signal_1311, signal_600}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_585 ( .s ({signal_2380, signal_2378}), .b ({signal_1084, signal_373}), .a ({signal_1027, signal_316}), .clk ( clk ), .r ( Fresh[409] ), .c ({signal_1312, signal_601}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_586 ( .s ({signal_2380, signal_2378}), .b ({signal_995, signal_285}), .a ({signal_1122, signal_411}), .clk ( clk ), .r ( Fresh[410] ), .c ({signal_1313, signal_602}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_587 ( .s ({signal_2380, signal_2378}), .b ({signal_2384, signal_2382}), .a ({signal_991, signal_281}), .clk ( clk ), .r ( Fresh[411] ), .c ({signal_1314, signal_603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_588 ( .s ({signal_2380, signal_2378}), .b ({signal_1025, signal_314}), .a ({signal_2484, signal_2482}), .clk ( clk ), .r ( Fresh[412] ), .c ({signal_1315, signal_604}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_589 ( .s ({signal_2508, signal_2502}), .b ({signal_1103, signal_392}), .a ({signal_1048, signal_337}), .clk ( clk ), .r ( Fresh[413] ), .c ({signal_1317, signal_605}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_590 ( .s ({signal_2380, signal_2378}), .b ({signal_944, signal_234}), .a ({signal_2424, signal_2422}), .clk ( clk ), .r ( Fresh[414] ), .c ({signal_1318, signal_606}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_591 ( .s ({signal_2380, signal_2378}), .b ({signal_971, signal_261}), .a ({signal_947, signal_237}), .clk ( clk ), .r ( Fresh[415] ), .c ({signal_1319, signal_607}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_592 ( .s ({signal_2380, signal_2378}), .b ({signal_982, signal_272}), .a ({signal_1117, signal_406}), .clk ( clk ), .r ( Fresh[416] ), .c ({signal_1320, signal_608}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_593 ( .s ({signal_2380, signal_2378}), .b ({signal_2412, signal_2410}), .a ({signal_1044, signal_333}), .clk ( clk ), .r ( Fresh[417] ), .c ({signal_1321, signal_609}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_594 ( .s ({signal_2380, signal_2378}), .b ({signal_1108, signal_397}), .a ({signal_995, signal_285}), .clk ( clk ), .r ( Fresh[418] ), .c ({signal_1322, signal_610}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_595 ( .s ({signal_2380, signal_2378}), .b ({signal_950, signal_240}), .a ({signal_999, signal_289}), .clk ( clk ), .r ( Fresh[419] ), .c ({signal_1323, signal_611}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_596 ( .s ({signal_2380, signal_2378}), .b ({signal_976, signal_266}), .a ({signal_1000, signal_290}), .clk ( clk ), .r ( Fresh[420] ), .c ({signal_1324, signal_612}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_597 ( .s ({signal_2380, signal_2378}), .b ({signal_1068, signal_357}), .a ({signal_1026, signal_315}), .clk ( clk ), .r ( Fresh[421] ), .c ({signal_1325, signal_613}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_598 ( .s ({signal_2380, signal_2378}), .b ({signal_2408, signal_2406}), .a ({signal_1082, signal_371}), .clk ( clk ), .r ( Fresh[422] ), .c ({signal_1326, signal_614}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_599 ( .s ({signal_2380, signal_2378}), .b ({signal_948, signal_238}), .a ({signal_2460, signal_2458}), .clk ( clk ), .r ( Fresh[423] ), .c ({signal_1327, signal_615}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_600 ( .s ({signal_2380, signal_2378}), .b ({signal_2472, signal_2470}), .a ({signal_972, signal_262}), .clk ( clk ), .r ( Fresh[424] ), .c ({signal_1328, signal_616}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_601 ( .s ({signal_2380, signal_2378}), .b ({signal_958, signal_248}), .a ({signal_1035, signal_324}), .clk ( clk ), .r ( Fresh[425] ), .c ({signal_1329, signal_617}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_602 ( .s ({signal_2380, signal_2378}), .b ({signal_974, signal_264}), .a ({signal_982, signal_272}), .clk ( clk ), .r ( Fresh[426] ), .c ({signal_1330, signal_618}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_603 ( .s ({signal_2380, signal_2378}), .b ({signal_1081, signal_370}), .a ({signal_2512, signal_2510}), .clk ( clk ), .r ( Fresh[427] ), .c ({signal_1331, signal_619}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_604 ( .s ({signal_2380, signal_2378}), .b ({signal_2516, signal_2514}), .a ({signal_1078, signal_367}), .clk ( clk ), .r ( Fresh[428] ), .c ({signal_1332, signal_620}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_605 ( .s ({signal_2380, signal_2378}), .b ({signal_1051, signal_340}), .a ({signal_954, signal_244}), .clk ( clk ), .r ( Fresh[429] ), .c ({signal_1333, signal_621}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_606 ( .s ({signal_2380, signal_2378}), .b ({signal_983, signal_273}), .a ({signal_958, signal_248}), .clk ( clk ), .r ( Fresh[430] ), .c ({signal_1334, signal_622}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_607 ( .s ({signal_2380, signal_2378}), .b ({signal_1068, signal_357}), .a ({signal_1126, signal_415}), .clk ( clk ), .r ( Fresh[431] ), .c ({signal_1335, signal_623}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_608 ( .s ({signal_2380, signal_2378}), .b ({signal_2520, signal_2518}), .a ({signal_1014, signal_303}), .clk ( clk ), .r ( Fresh[432] ), .c ({signal_1336, signal_624}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_609 ( .s ({signal_2380, signal_2378}), .b ({signal_1029, signal_318}), .a ({signal_977, signal_267}), .clk ( clk ), .r ( Fresh[433] ), .c ({signal_1337, signal_625}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_610 ( .s ({signal_2380, signal_2378}), .b ({signal_1042, signal_331}), .a ({signal_1037, signal_326}), .clk ( clk ), .r ( Fresh[434] ), .c ({signal_1338, signal_626}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_611 ( .s ({signal_2380, signal_2378}), .b ({signal_1038, signal_327}), .a ({signal_1057, signal_346}), .clk ( clk ), .r ( Fresh[435] ), .c ({signal_1339, signal_627}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_612 ( .s ({signal_2380, signal_2378}), .b ({signal_995, signal_285}), .a ({signal_973, signal_263}), .clk ( clk ), .r ( Fresh[436] ), .c ({signal_1340, signal_628}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_613 ( .s ({signal_2380, signal_2378}), .b ({signal_1099, signal_388}), .a ({signal_946, signal_236}), .clk ( clk ), .r ( Fresh[437] ), .c ({signal_1341, signal_629}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_614 ( .s ({signal_2380, signal_2378}), .b ({signal_990, signal_280}), .a ({signal_966, signal_256}), .clk ( clk ), .r ( Fresh[438] ), .c ({signal_1342, signal_630}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_615 ( .s ({signal_2380, signal_2378}), .b ({signal_1077, signal_366}), .a ({signal_1126, signal_415}), .clk ( clk ), .r ( Fresh[439] ), .c ({signal_1343, signal_631}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_616 ( .s ({signal_2380, signal_2378}), .b ({signal_1091, signal_380}), .a ({signal_981, signal_271}), .clk ( clk ), .r ( Fresh[440] ), .c ({signal_1344, signal_632}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_617 ( .s ({signal_2380, signal_2378}), .b ({signal_1013, signal_302}), .a ({signal_944, signal_234}), .clk ( clk ), .r ( Fresh[441] ), .c ({signal_1345, signal_633}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_618 ( .s ({signal_2380, signal_2378}), .b ({signal_1057, signal_346}), .a ({signal_1060, signal_349}), .clk ( clk ), .r ( Fresh[442] ), .c ({signal_1346, signal_634}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_619 ( .s ({signal_2380, signal_2378}), .b ({signal_1026, signal_315}), .a ({signal_977, signal_267}), .clk ( clk ), .r ( Fresh[443] ), .c ({signal_1347, signal_635}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_620 ( .s ({signal_2380, signal_2378}), .b ({signal_1107, signal_396}), .a ({signal_1018, signal_307}), .clk ( clk ), .r ( Fresh[444] ), .c ({signal_1348, signal_636}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_621 ( .s ({signal_2380, signal_2378}), .b ({signal_2412, signal_2410}), .a ({signal_1114, signal_403}), .clk ( clk ), .r ( Fresh[445] ), .c ({signal_1349, signal_637}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_622 ( .s ({signal_2380, signal_2378}), .b ({signal_943, signal_233}), .a ({signal_942, signal_232}), .clk ( clk ), .r ( Fresh[446] ), .c ({signal_1350, signal_638}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_623 ( .s ({signal_2380, signal_2378}), .b ({signal_1089, signal_378}), .a ({signal_2528, signal_2524}), .clk ( clk ), .r ( Fresh[447] ), .c ({signal_1351, signal_639}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_624 ( .s ({signal_2380, signal_2378}), .b ({signal_1075, signal_364}), .a ({signal_967, signal_257}), .clk ( clk ), .r ( Fresh[448] ), .c ({signal_1352, signal_640}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_625 ( .s ({signal_2380, signal_2378}), .b ({signal_1023, signal_312}), .a ({signal_989, signal_279}), .clk ( clk ), .r ( Fresh[449] ), .c ({signal_1353, signal_641}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_626 ( .s ({signal_2380, signal_2378}), .b ({signal_2532, signal_2530}), .a ({signal_1019, signal_308}), .clk ( clk ), .r ( Fresh[450] ), .c ({signal_1354, signal_642}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_627 ( .s ({signal_2380, signal_2378}), .b ({signal_1090, signal_379}), .a ({signal_953, signal_243}), .clk ( clk ), .r ( Fresh[451] ), .c ({signal_1355, signal_643}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_628 ( .s ({signal_2380, signal_2378}), .b ({signal_1070, signal_359}), .a ({signal_947, signal_237}), .clk ( clk ), .r ( Fresh[452] ), .c ({signal_1356, signal_644}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_629 ( .s ({signal_2380, signal_2378}), .b ({signal_958, signal_248}), .a ({signal_1054, signal_343}), .clk ( clk ), .r ( Fresh[453] ), .c ({signal_1357, signal_645}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_630 ( .s ({signal_2380, signal_2378}), .b ({signal_977, signal_267}), .a ({signal_2464, signal_2462}), .clk ( clk ), .r ( Fresh[454] ), .c ({signal_1358, signal_646}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_631 ( .s ({signal_2380, signal_2378}), .b ({signal_1064, signal_353}), .a ({signal_1033, signal_322}), .clk ( clk ), .r ( Fresh[455] ), .c ({signal_1359, signal_647}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_632 ( .s ({signal_2380, signal_2378}), .b ({signal_993, signal_283}), .a ({signal_1002, signal_292}), .clk ( clk ), .r ( Fresh[456] ), .c ({signal_1360, signal_648}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_633 ( .s ({signal_2380, signal_2378}), .b ({signal_1071, signal_360}), .a ({signal_1068, signal_357}), .clk ( clk ), .r ( Fresh[457] ), .c ({signal_1361, signal_649}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_634 ( .s ({signal_2380, signal_2378}), .b ({signal_2452, signal_2450}), .a ({signal_958, signal_248}), .clk ( clk ), .r ( Fresh[458] ), .c ({signal_1362, signal_650}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_635 ( .s ({signal_2380, signal_2378}), .b ({signal_2536, signal_2534}), .a ({signal_1079, signal_368}), .clk ( clk ), .r ( Fresh[459] ), .c ({signal_1363, signal_651}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_636 ( .s ({signal_2380, signal_2378}), .b ({signal_1008, signal_297}), .a ({signal_1050, signal_339}), .clk ( clk ), .r ( Fresh[460] ), .c ({signal_1364, signal_652}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_637 ( .s ({signal_2380, signal_2378}), .b ({signal_1090, signal_379}), .a ({signal_962, signal_252}), .clk ( clk ), .r ( Fresh[461] ), .c ({signal_1365, signal_653}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_638 ( .s ({signal_2380, signal_2378}), .b ({signal_950, signal_240}), .a ({signal_995, signal_285}), .clk ( clk ), .r ( Fresh[462] ), .c ({signal_1366, signal_654}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_639 ( .s ({signal_2380, signal_2378}), .b ({signal_1034, signal_323}), .a ({signal_1025, signal_314}), .clk ( clk ), .r ( Fresh[463] ), .c ({signal_1367, signal_655}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_640 ( .s ({signal_2380, signal_2378}), .b ({signal_945, signal_235}), .a ({signal_1101, signal_390}), .clk ( clk ), .r ( Fresh[464] ), .c ({signal_1368, signal_656}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_641 ( .s ({signal_2380, signal_2378}), .b ({signal_1115, signal_404}), .a ({signal_984, signal_274}), .clk ( clk ), .r ( Fresh[465] ), .c ({signal_1369, signal_657}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_642 ( .s ({signal_2380, signal_2378}), .b ({signal_1086, signal_375}), .a ({signal_1027, signal_316}), .clk ( clk ), .r ( Fresh[466] ), .c ({signal_1370, signal_658}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_643 ( .s ({signal_2380, signal_2378}), .b ({signal_1116, signal_405}), .a ({signal_1071, signal_360}), .clk ( clk ), .r ( Fresh[467] ), .c ({signal_1371, signal_659}) ) ;
    buf_clk cell_1092 ( .C ( clk ), .D ( signal_2537 ), .Q ( signal_2538 ) ) ;
    buf_clk cell_1094 ( .C ( clk ), .D ( signal_2539 ), .Q ( signal_2540 ) ) ;
    buf_clk cell_1096 ( .C ( clk ), .D ( signal_2541 ), .Q ( signal_2542 ) ) ;
    buf_clk cell_1098 ( .C ( clk ), .D ( signal_2543 ), .Q ( signal_2544 ) ) ;
    buf_clk cell_1100 ( .C ( clk ), .D ( signal_2545 ), .Q ( signal_2546 ) ) ;
    buf_clk cell_1102 ( .C ( clk ), .D ( signal_2547 ), .Q ( signal_2548 ) ) ;
    buf_clk cell_1104 ( .C ( clk ), .D ( signal_2549 ), .Q ( signal_2550 ) ) ;
    buf_clk cell_1106 ( .C ( clk ), .D ( signal_2551 ), .Q ( signal_2552 ) ) ;
    buf_clk cell_1108 ( .C ( clk ), .D ( signal_2553 ), .Q ( signal_2554 ) ) ;
    buf_clk cell_1110 ( .C ( clk ), .D ( signal_2555 ), .Q ( signal_2556 ) ) ;
    buf_clk cell_1112 ( .C ( clk ), .D ( signal_2557 ), .Q ( signal_2558 ) ) ;
    buf_clk cell_1114 ( .C ( clk ), .D ( signal_2559 ), .Q ( signal_2560 ) ) ;
    buf_clk cell_1116 ( .C ( clk ), .D ( signal_2561 ), .Q ( signal_2562 ) ) ;
    buf_clk cell_1118 ( .C ( clk ), .D ( signal_2563 ), .Q ( signal_2564 ) ) ;
    buf_clk cell_1120 ( .C ( clk ), .D ( signal_2565 ), .Q ( signal_2566 ) ) ;
    buf_clk cell_1122 ( .C ( clk ), .D ( signal_2567 ), .Q ( signal_2568 ) ) ;
    buf_clk cell_1124 ( .C ( clk ), .D ( signal_2569 ), .Q ( signal_2570 ) ) ;
    buf_clk cell_1126 ( .C ( clk ), .D ( signal_2571 ), .Q ( signal_2572 ) ) ;
    buf_clk cell_1128 ( .C ( clk ), .D ( signal_2573 ), .Q ( signal_2574 ) ) ;
    buf_clk cell_1130 ( .C ( clk ), .D ( signal_2575 ), .Q ( signal_2576 ) ) ;
    buf_clk cell_1138 ( .C ( clk ), .D ( signal_2583 ), .Q ( signal_2584 ) ) ;
    buf_clk cell_1148 ( .C ( clk ), .D ( signal_2593 ), .Q ( signal_2594 ) ) ;
    buf_clk cell_1162 ( .C ( clk ), .D ( signal_2607 ), .Q ( signal_2608 ) ) ;
    buf_clk cell_1174 ( .C ( clk ), .D ( signal_2619 ), .Q ( signal_2620 ) ) ;
    buf_clk cell_1186 ( .C ( clk ), .D ( signal_2631 ), .Q ( signal_2632 ) ) ;
    buf_clk cell_1200 ( .C ( clk ), .D ( signal_2645 ), .Q ( signal_2646 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_1139 ( .C ( clk ), .D ( signal_2584 ), .Q ( signal_2585 ) ) ;
    buf_clk cell_1149 ( .C ( clk ), .D ( signal_2594 ), .Q ( signal_2595 ) ) ;
    buf_clk cell_1151 ( .C ( clk ), .D ( signal_605 ), .Q ( signal_2597 ) ) ;
    buf_clk cell_1153 ( .C ( clk ), .D ( signal_1317 ), .Q ( signal_2599 ) ) ;
    buf_clk cell_1163 ( .C ( clk ), .D ( signal_2608 ), .Q ( signal_2609 ) ) ;
    buf_clk cell_1175 ( .C ( clk ), .D ( signal_2620 ), .Q ( signal_2621 ) ) ;
    buf_clk cell_1187 ( .C ( clk ), .D ( signal_2632 ), .Q ( signal_2633 ) ) ;
    buf_clk cell_1201 ( .C ( clk ), .D ( signal_2646 ), .Q ( signal_2647 ) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_644 ( .s ({signal_2540, signal_2538}), .b ({signal_1189, signal_478}), .a ({signal_1351, signal_639}), .clk ( clk ), .r ( Fresh[468] ), .c ({signal_1372, signal_660}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_645 ( .s ({signal_2540, signal_2538}), .b ({signal_1325, signal_613}), .a ({signal_1172, signal_461}), .clk ( clk ), .r ( Fresh[469] ), .c ({signal_1373, signal_661}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_646 ( .s ({signal_2540, signal_2538}), .b ({signal_1275, signal_564}), .a ({signal_1281, signal_570}), .clk ( clk ), .r ( Fresh[470] ), .c ({signal_1374, signal_662}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_647 ( .s ({signal_2540, signal_2538}), .b ({signal_1332, signal_620}), .a ({signal_1319, signal_607}), .clk ( clk ), .r ( Fresh[471] ), .c ({signal_1375, signal_663}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_648 ( .s ({signal_2540, signal_2538}), .b ({signal_1369, signal_657}), .a ({signal_1150, signal_439}), .clk ( clk ), .r ( Fresh[472] ), .c ({signal_1376, signal_664}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_649 ( .s ({signal_2540, signal_2538}), .b ({signal_1344, signal_632}), .a ({signal_1349, signal_637}), .clk ( clk ), .r ( Fresh[473] ), .c ({signal_1377, signal_665}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_650 ( .s ({signal_2540, signal_2538}), .b ({signal_1304, signal_593}), .a ({signal_1353, signal_641}), .clk ( clk ), .r ( Fresh[474] ), .c ({signal_1378, signal_666}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_651 ( .s ({signal_2540, signal_2538}), .b ({signal_1146, signal_435}), .a ({signal_1162, signal_451}), .clk ( clk ), .r ( Fresh[475] ), .c ({signal_1379, signal_667}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_652 ( .s ({signal_2540, signal_2538}), .b ({signal_1132, signal_421}), .a ({signal_1203, signal_492}), .clk ( clk ), .r ( Fresh[476] ), .c ({signal_1380, signal_668}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_653 ( .s ({signal_2540, signal_2538}), .b ({signal_1302, signal_591}), .a ({signal_1241, signal_530}), .clk ( clk ), .r ( Fresh[477] ), .c ({signal_1381, signal_669}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_654 ( .s ({signal_2540, signal_2538}), .b ({signal_1171, signal_460}), .a ({signal_1274, signal_563}), .clk ( clk ), .r ( Fresh[478] ), .c ({signal_1382, signal_670}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_655 ( .s ({signal_2540, signal_2538}), .b ({signal_1228, signal_517}), .a ({signal_1321, signal_609}), .clk ( clk ), .r ( Fresh[479] ), .c ({signal_1383, signal_671}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_656 ( .s ({signal_2540, signal_2538}), .b ({signal_1254, signal_543}), .a ({signal_1295, signal_584}), .clk ( clk ), .r ( Fresh[480] ), .c ({signal_1384, signal_672}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_657 ( .s ({signal_2540, signal_2538}), .b ({signal_2544, signal_2542}), .a ({signal_1233, signal_522}), .clk ( clk ), .r ( Fresh[481] ), .c ({signal_1385, signal_673}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_658 ( .s ({signal_2540, signal_2538}), .b ({signal_1249, signal_538}), .a ({signal_2548, signal_2546}), .clk ( clk ), .r ( Fresh[482] ), .c ({signal_1386, signal_674}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_659 ( .s ({signal_2540, signal_2538}), .b ({signal_1149, signal_438}), .a ({signal_1318, signal_606}), .clk ( clk ), .r ( Fresh[483] ), .c ({signal_1387, signal_675}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_660 ( .s ({signal_2540, signal_2538}), .b ({signal_1131, signal_420}), .a ({signal_1306, signal_595}), .clk ( clk ), .r ( Fresh[484] ), .c ({signal_1388, signal_676}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_661 ( .s ({signal_2540, signal_2538}), .b ({signal_1139, signal_428}), .a ({signal_1242, signal_531}), .clk ( clk ), .r ( Fresh[485] ), .c ({signal_1389, signal_677}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_662 ( .s ({signal_2540, signal_2538}), .b ({signal_1362, signal_650}), .a ({signal_1348, signal_636}), .clk ( clk ), .r ( Fresh[486] ), .c ({signal_1390, signal_678}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_663 ( .s ({signal_2540, signal_2538}), .b ({signal_1268, signal_557}), .a ({signal_1160, signal_449}), .clk ( clk ), .r ( Fresh[487] ), .c ({signal_1391, signal_679}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_664 ( .s ({signal_2540, signal_2538}), .b ({signal_1220, signal_509}), .a ({signal_1310, signal_599}), .clk ( clk ), .r ( Fresh[488] ), .c ({signal_1392, signal_680}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_665 ( .s ({signal_2540, signal_2538}), .b ({signal_1230, signal_519}), .a ({signal_1350, signal_638}), .clk ( clk ), .r ( Fresh[489] ), .c ({signal_1393, signal_681}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_666 ( .s ({signal_2540, signal_2538}), .b ({signal_1128, signal_417}), .a ({signal_1130, signal_419}), .clk ( clk ), .r ( Fresh[490] ), .c ({signal_1394, signal_682}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_667 ( .s ({signal_2540, signal_2538}), .b ({signal_1328, signal_616}), .a ({signal_1298, signal_587}), .clk ( clk ), .r ( Fresh[491] ), .c ({signal_1395, signal_683}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_668 ( .s ({signal_2540, signal_2538}), .b ({signal_1193, signal_482}), .a ({signal_2552, signal_2550}), .clk ( clk ), .r ( Fresh[492] ), .c ({signal_1396, signal_684}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_669 ( .s ({signal_2540, signal_2538}), .b ({signal_1144, signal_433}), .a ({signal_1140, signal_429}), .clk ( clk ), .r ( Fresh[493] ), .c ({signal_1397, signal_685}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_670 ( .s ({signal_2540, signal_2538}), .b ({signal_1165, signal_454}), .a ({signal_1322, signal_610}), .clk ( clk ), .r ( Fresh[494] ), .c ({signal_1398, signal_686}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_671 ( .s ({signal_2540, signal_2538}), .b ({signal_1358, signal_646}), .a ({signal_1367, signal_655}), .clk ( clk ), .r ( Fresh[495] ), .c ({signal_1399, signal_687}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_672 ( .s ({signal_2540, signal_2538}), .b ({signal_1243, signal_532}), .a ({signal_1307, signal_596}), .clk ( clk ), .r ( Fresh[496] ), .c ({signal_1400, signal_688}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_673 ( .s ({signal_2540, signal_2538}), .b ({signal_1315, signal_604}), .a ({signal_1161, signal_450}), .clk ( clk ), .r ( Fresh[497] ), .c ({signal_1401, signal_689}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_674 ( .s ({signal_2540, signal_2538}), .b ({signal_1337, signal_625}), .a ({signal_1324, signal_612}), .clk ( clk ), .r ( Fresh[498] ), .c ({signal_1402, signal_690}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_675 ( .s ({signal_2540, signal_2538}), .b ({signal_1167, signal_456}), .a ({signal_1284, signal_573}), .clk ( clk ), .r ( Fresh[499] ), .c ({signal_1403, signal_691}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_676 ( .s ({signal_2540, signal_2538}), .b ({signal_1333, signal_621}), .a ({signal_1195, signal_484}), .clk ( clk ), .r ( Fresh[500] ), .c ({signal_1404, signal_692}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_677 ( .s ({signal_2540, signal_2538}), .b ({signal_1272, signal_561}), .a ({signal_1186, signal_475}), .clk ( clk ), .r ( Fresh[501] ), .c ({signal_1405, signal_693}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_678 ( .s ({signal_2540, signal_2538}), .b ({signal_1202, signal_491}), .a ({signal_1184, signal_473}), .clk ( clk ), .r ( Fresh[502] ), .c ({signal_1406, signal_694}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_679 ( .s ({signal_2540, signal_2538}), .b ({signal_1253, signal_542}), .a ({signal_1238, signal_527}), .clk ( clk ), .r ( Fresh[503] ), .c ({signal_1407, signal_695}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_680 ( .s ({signal_2540, signal_2538}), .b ({signal_1185, signal_474}), .a ({signal_2556, signal_2554}), .clk ( clk ), .r ( Fresh[504] ), .c ({signal_1408, signal_696}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_681 ( .s ({signal_2540, signal_2538}), .b ({signal_1354, signal_642}), .a ({signal_1261, signal_550}), .clk ( clk ), .r ( Fresh[505] ), .c ({signal_1409, signal_697}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_682 ( .s ({signal_2540, signal_2538}), .b ({signal_1276, signal_565}), .a ({signal_1188, signal_477}), .clk ( clk ), .r ( Fresh[506] ), .c ({signal_1410, signal_698}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_683 ( .s ({signal_2540, signal_2538}), .b ({signal_1216, signal_505}), .a ({signal_1226, signal_515}), .clk ( clk ), .r ( Fresh[507] ), .c ({signal_1411, signal_699}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_684 ( .s ({signal_2540, signal_2538}), .b ({signal_1287, signal_576}), .a ({signal_1313, signal_602}), .clk ( clk ), .r ( Fresh[508] ), .c ({signal_1412, signal_700}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_685 ( .s ({signal_2540, signal_2538}), .b ({signal_1232, signal_521}), .a ({signal_1135, signal_424}), .clk ( clk ), .r ( Fresh[509] ), .c ({signal_1413, signal_701}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_686 ( .s ({signal_2540, signal_2538}), .b ({signal_1326, signal_614}), .a ({signal_1280, signal_569}), .clk ( clk ), .r ( Fresh[510] ), .c ({signal_1414, signal_702}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_687 ( .s ({signal_2540, signal_2538}), .b ({signal_1365, signal_653}), .a ({signal_1368, signal_656}), .clk ( clk ), .r ( Fresh[511] ), .c ({signal_1415, signal_703}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_688 ( .s ({signal_2540, signal_2538}), .b ({signal_1215, signal_504}), .a ({signal_1266, signal_555}), .clk ( clk ), .r ( Fresh[512] ), .c ({signal_1416, signal_704}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_689 ( .s ({signal_2540, signal_2538}), .b ({signal_1156, signal_445}), .a ({signal_1252, signal_541}), .clk ( clk ), .r ( Fresh[513] ), .c ({signal_1417, signal_705}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_690 ( .s ({signal_2540, signal_2538}), .b ({signal_1177, signal_466}), .a ({signal_1197, signal_486}), .clk ( clk ), .r ( Fresh[514] ), .c ({signal_1418, signal_706}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_691 ( .s ({signal_2540, signal_2538}), .b ({signal_1297, signal_586}), .a ({signal_1323, signal_611}), .clk ( clk ), .r ( Fresh[515] ), .c ({signal_1419, signal_707}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_692 ( .s ({signal_2540, signal_2538}), .b ({signal_1179, signal_468}), .a ({signal_1255, signal_544}), .clk ( clk ), .r ( Fresh[516] ), .c ({signal_1420, signal_708}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_693 ( .s ({signal_2540, signal_2538}), .b ({signal_1314, signal_603}), .a ({signal_1163, signal_452}), .clk ( clk ), .r ( Fresh[517] ), .c ({signal_1421, signal_709}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_694 ( .s ({signal_2540, signal_2538}), .b ({signal_2560, signal_2558}), .a ({signal_1256, signal_545}), .clk ( clk ), .r ( Fresh[518] ), .c ({signal_1422, signal_710}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_695 ( .s ({signal_2540, signal_2538}), .b ({signal_1331, signal_619}), .a ({signal_1210, signal_499}), .clk ( clk ), .r ( Fresh[519] ), .c ({signal_1423, signal_711}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_696 ( .s ({signal_2540, signal_2538}), .b ({signal_1258, signal_547}), .a ({signal_1194, signal_483}), .clk ( clk ), .r ( Fresh[520] ), .c ({signal_1424, signal_712}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_697 ( .s ({signal_2540, signal_2538}), .b ({signal_1343, signal_631}), .a ({signal_1199, signal_488}), .clk ( clk ), .r ( Fresh[521] ), .c ({signal_1425, signal_713}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_698 ( .s ({signal_2540, signal_2538}), .b ({signal_1264, signal_553}), .a ({signal_1154, signal_443}), .clk ( clk ), .r ( Fresh[522] ), .c ({signal_1426, signal_714}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_699 ( .s ({signal_2540, signal_2538}), .b ({signal_1265, signal_554}), .a ({signal_1234, signal_523}), .clk ( clk ), .r ( Fresh[523] ), .c ({signal_1427, signal_715}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_700 ( .s ({signal_2540, signal_2538}), .b ({signal_1178, signal_467}), .a ({signal_1247, signal_536}), .clk ( clk ), .r ( Fresh[524] ), .c ({signal_1428, signal_716}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_701 ( .s ({signal_2540, signal_2538}), .b ({signal_1138, signal_427}), .a ({signal_1292, signal_581}), .clk ( clk ), .r ( Fresh[525] ), .c ({signal_1429, signal_717}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_702 ( .s ({signal_2540, signal_2538}), .b ({signal_1155, signal_444}), .a ({signal_1341, signal_629}), .clk ( clk ), .r ( Fresh[526] ), .c ({signal_1430, signal_718}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_703 ( .s ({signal_2540, signal_2538}), .b ({signal_1181, signal_470}), .a ({signal_1342, signal_630}), .clk ( clk ), .r ( Fresh[527] ), .c ({signal_1431, signal_719}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_704 ( .s ({signal_2540, signal_2538}), .b ({signal_1166, signal_455}), .a ({signal_1340, signal_628}), .clk ( clk ), .r ( Fresh[528] ), .c ({signal_1432, signal_720}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_705 ( .s ({signal_2540, signal_2538}), .b ({signal_1359, signal_647}), .a ({signal_1269, signal_558}), .clk ( clk ), .r ( Fresh[529] ), .c ({signal_1433, signal_721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_706 ( .s ({signal_2540, signal_2538}), .b ({signal_1148, signal_437}), .a ({signal_1339, signal_627}), .clk ( clk ), .r ( Fresh[530] ), .c ({signal_1434, signal_722}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_707 ( .s ({signal_2540, signal_2538}), .b ({signal_1201, signal_490}), .a ({signal_1237, signal_526}), .clk ( clk ), .r ( Fresh[531] ), .c ({signal_1435, signal_723}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_708 ( .s ({signal_2540, signal_2538}), .b ({signal_1227, signal_516}), .a ({signal_1320, signal_608}), .clk ( clk ), .r ( Fresh[532] ), .c ({signal_1436, signal_724}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_709 ( .s ({signal_2540, signal_2538}), .b ({signal_1225, signal_514}), .a ({signal_1366, signal_654}), .clk ( clk ), .r ( Fresh[533] ), .c ({signal_1437, signal_725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_710 ( .s ({signal_2540, signal_2538}), .b ({signal_1127, signal_416}), .a ({signal_1222, signal_511}), .clk ( clk ), .r ( Fresh[534] ), .c ({signal_1438, signal_726}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_711 ( .s ({signal_2540, signal_2538}), .b ({signal_1299, signal_588}), .a ({signal_1142, signal_431}), .clk ( clk ), .r ( Fresh[535] ), .c ({signal_1439, signal_727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_712 ( .s ({signal_2540, signal_2538}), .b ({signal_1240, signal_529}), .a ({signal_1190, signal_479}), .clk ( clk ), .r ( Fresh[536] ), .c ({signal_1440, signal_728}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_713 ( .s ({signal_2540, signal_2538}), .b ({signal_2564, signal_2562}), .a ({signal_1335, signal_623}), .clk ( clk ), .r ( Fresh[537] ), .c ({signal_1441, signal_729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_714 ( .s ({signal_2540, signal_2538}), .b ({signal_1278, signal_567}), .a ({signal_1279, signal_568}), .clk ( clk ), .r ( Fresh[538] ), .c ({signal_1442, signal_730}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_715 ( .s ({signal_2540, signal_2538}), .b ({signal_1257, signal_546}), .a ({signal_1357, signal_645}), .clk ( clk ), .r ( Fresh[539] ), .c ({signal_1443, signal_731}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_716 ( .s ({signal_2540, signal_2538}), .b ({signal_1204, signal_493}), .a ({signal_1219, signal_508}), .clk ( clk ), .r ( Fresh[540] ), .c ({signal_1444, signal_732}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_717 ( .s ({signal_2540, signal_2538}), .b ({signal_1277, signal_566}), .a ({signal_1136, signal_425}), .clk ( clk ), .r ( Fresh[541] ), .c ({signal_1445, signal_733}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_718 ( .s ({signal_2540, signal_2538}), .b ({signal_1206, signal_495}), .a ({signal_2568, signal_2566}), .clk ( clk ), .r ( Fresh[542] ), .c ({signal_1446, signal_734}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_719 ( .s ({signal_2540, signal_2538}), .b ({signal_1221, signal_510}), .a ({signal_1159, signal_448}), .clk ( clk ), .r ( Fresh[543] ), .c ({signal_1447, signal_735}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_720 ( .s ({signal_2540, signal_2538}), .b ({signal_1296, signal_585}), .a ({signal_1129, signal_418}), .clk ( clk ), .r ( Fresh[544] ), .c ({signal_1448, signal_736}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_721 ( .s ({signal_2540, signal_2538}), .b ({signal_2572, signal_2570}), .a ({signal_1180, signal_469}), .clk ( clk ), .r ( Fresh[545] ), .c ({signal_1449, signal_737}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_722 ( .s ({signal_2540, signal_2538}), .b ({signal_1134, signal_423}), .a ({signal_1198, signal_487}), .clk ( clk ), .r ( Fresh[546] ), .c ({signal_1450, signal_738}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_723 ( .s ({signal_2540, signal_2538}), .b ({signal_1345, signal_633}), .a ({signal_1288, signal_577}), .clk ( clk ), .r ( Fresh[547] ), .c ({signal_1451, signal_739}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_724 ( .s ({signal_2540, signal_2538}), .b ({signal_1229, signal_518}), .a ({signal_1363, signal_651}), .clk ( clk ), .r ( Fresh[548] ), .c ({signal_1452, signal_740}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_725 ( .s ({signal_2540, signal_2538}), .b ({signal_1289, signal_578}), .a ({signal_1267, signal_556}), .clk ( clk ), .r ( Fresh[549] ), .c ({signal_1453, signal_741}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_726 ( .s ({signal_2540, signal_2538}), .b ({signal_1244, signal_533}), .a ({signal_1151, signal_440}), .clk ( clk ), .r ( Fresh[550] ), .c ({signal_1454, signal_742}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_727 ( .s ({signal_2540, signal_2538}), .b ({signal_1183, signal_472}), .a ({signal_1371, signal_659}), .clk ( clk ), .r ( Fresh[551] ), .c ({signal_1455, signal_743}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_728 ( .s ({signal_2540, signal_2538}), .b ({signal_1308, signal_597}), .a ({signal_1294, signal_583}), .clk ( clk ), .r ( Fresh[552] ), .c ({signal_1456, signal_744}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_729 ( .s ({signal_2540, signal_2538}), .b ({signal_1212, signal_501}), .a ({signal_1152, signal_441}), .clk ( clk ), .r ( Fresh[553] ), .c ({signal_1457, signal_745}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_730 ( .s ({signal_2540, signal_2538}), .b ({signal_1334, signal_622}), .a ({signal_1263, signal_552}), .clk ( clk ), .r ( Fresh[554] ), .c ({signal_1458, signal_746}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_731 ( .s ({signal_2540, signal_2538}), .b ({signal_1231, signal_520}), .a ({signal_1137, signal_426}), .clk ( clk ), .r ( Fresh[555] ), .c ({signal_1459, signal_747}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_732 ( .s ({signal_2540, signal_2538}), .b ({signal_1217, signal_506}), .a ({signal_1291, signal_580}), .clk ( clk ), .r ( Fresh[556] ), .c ({signal_1460, signal_748}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_733 ( .s ({signal_2540, signal_2538}), .b ({signal_1207, signal_496}), .a ({signal_1157, signal_446}), .clk ( clk ), .r ( Fresh[557] ), .c ({signal_1461, signal_749}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_734 ( .s ({signal_2540, signal_2538}), .b ({signal_2576, signal_2574}), .a ({signal_1205, signal_494}), .clk ( clk ), .r ( Fresh[558] ), .c ({signal_1462, signal_750}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_735 ( .s ({signal_2540, signal_2538}), .b ({signal_1196, signal_485}), .a ({signal_1364, signal_652}), .clk ( clk ), .r ( Fresh[559] ), .c ({signal_1463, signal_751}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_736 ( .s ({signal_2540, signal_2538}), .b ({signal_1271, signal_560}), .a ({signal_1260, signal_549}), .clk ( clk ), .r ( Fresh[560] ), .c ({signal_1464, signal_752}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_737 ( .s ({signal_2540, signal_2538}), .b ({signal_1246, signal_535}), .a ({signal_1282, signal_571}), .clk ( clk ), .r ( Fresh[561] ), .c ({signal_1465, signal_753}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_738 ( .s ({signal_2540, signal_2538}), .b ({signal_1361, signal_649}), .a ({signal_1327, signal_615}), .clk ( clk ), .r ( Fresh[562] ), .c ({signal_1466, signal_754}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_739 ( .s ({signal_2540, signal_2538}), .b ({signal_1236, signal_525}), .a ({signal_1259, signal_548}), .clk ( clk ), .r ( Fresh[563] ), .c ({signal_1467, signal_755}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_740 ( .s ({signal_2540, signal_2538}), .b ({signal_1262, signal_551}), .a ({signal_1245, signal_534}), .clk ( clk ), .r ( Fresh[564] ), .c ({signal_1468, signal_756}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_741 ( .s ({signal_2540, signal_2538}), .b ({signal_1182, signal_471}), .a ({signal_1251, signal_540}), .clk ( clk ), .r ( Fresh[565] ), .c ({signal_1469, signal_757}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_742 ( .s ({signal_2540, signal_2538}), .b ({signal_1347, signal_635}), .a ({signal_1305, signal_594}), .clk ( clk ), .r ( Fresh[566] ), .c ({signal_1470, signal_758}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_743 ( .s ({signal_2540, signal_2538}), .b ({signal_1370, signal_658}), .a ({signal_1235, signal_524}), .clk ( clk ), .r ( Fresh[567] ), .c ({signal_1471, signal_759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_744 ( .s ({signal_2540, signal_2538}), .b ({signal_1158, signal_447}), .a ({signal_1175, signal_464}), .clk ( clk ), .r ( Fresh[568] ), .c ({signal_1472, signal_760}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_745 ( .s ({signal_2540, signal_2538}), .b ({signal_1286, signal_575}), .a ({signal_1270, signal_559}), .clk ( clk ), .r ( Fresh[569] ), .c ({signal_1473, signal_761}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_746 ( .s ({signal_2540, signal_2538}), .b ({signal_1262, signal_551}), .a ({signal_1330, signal_618}), .clk ( clk ), .r ( Fresh[570] ), .c ({signal_1474, signal_762}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_747 ( .s ({signal_2540, signal_2538}), .b ({signal_1192, signal_481}), .a ({signal_1250, signal_539}), .clk ( clk ), .r ( Fresh[571] ), .c ({signal_1475, signal_763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_748 ( .s ({signal_2540, signal_2538}), .b ({signal_1200, signal_489}), .a ({signal_1329, signal_617}), .clk ( clk ), .r ( Fresh[572] ), .c ({signal_1476, signal_764}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_749 ( .s ({signal_2540, signal_2538}), .b ({signal_1248, signal_537}), .a ({signal_1283, signal_572}), .clk ( clk ), .r ( Fresh[573] ), .c ({signal_1477, signal_765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_750 ( .s ({signal_2540, signal_2538}), .b ({signal_1356, signal_644}), .a ({signal_1174, signal_463}), .clk ( clk ), .r ( Fresh[574] ), .c ({signal_1478, signal_766}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_751 ( .s ({signal_2540, signal_2538}), .b ({signal_1164, signal_453}), .a ({signal_1192, signal_481}), .clk ( clk ), .r ( Fresh[575] ), .c ({signal_1479, signal_767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_752 ( .s ({signal_2540, signal_2538}), .b ({signal_1209, signal_498}), .a ({signal_1293, signal_582}), .clk ( clk ), .r ( Fresh[576] ), .c ({signal_1480, signal_768}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_753 ( .s ({signal_2540, signal_2538}), .b ({signal_1285, signal_574}), .a ({signal_1346, signal_634}), .clk ( clk ), .r ( Fresh[577] ), .c ({signal_1481, signal_769}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_754 ( .s ({signal_2540, signal_2538}), .b ({signal_1176, signal_465}), .a ({signal_1141, signal_430}), .clk ( clk ), .r ( Fresh[578] ), .c ({signal_1482, signal_770}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_755 ( .s ({signal_2540, signal_2538}), .b ({signal_1168, signal_457}), .a ({signal_1338, signal_626}), .clk ( clk ), .r ( Fresh[579] ), .c ({signal_1483, signal_771}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_756 ( .s ({signal_2540, signal_2538}), .b ({signal_1336, signal_624}), .a ({signal_1224, signal_513}), .clk ( clk ), .r ( Fresh[580] ), .c ({signal_1484, signal_772}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_757 ( .s ({signal_2540, signal_2538}), .b ({signal_1223, signal_512}), .a ({signal_1208, signal_497}), .clk ( clk ), .r ( Fresh[581] ), .c ({signal_1485, signal_773}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_758 ( .s ({signal_2540, signal_2538}), .b ({signal_1187, signal_476}), .a ({signal_1211, signal_500}), .clk ( clk ), .r ( Fresh[582] ), .c ({signal_1486, signal_774}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_759 ( .s ({signal_2540, signal_2538}), .b ({signal_1360, signal_648}), .a ({signal_1303, signal_592}), .clk ( clk ), .r ( Fresh[583] ), .c ({signal_1487, signal_775}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_760 ( .s ({signal_2540, signal_2538}), .b ({signal_1239, signal_528}), .a ({signal_1173, signal_462}), .clk ( clk ), .r ( Fresh[584] ), .c ({signal_1488, signal_776}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_761 ( .s ({signal_2540, signal_2538}), .b ({signal_1218, signal_507}), .a ({signal_1300, signal_589}), .clk ( clk ), .r ( Fresh[585] ), .c ({signal_1489, signal_777}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_762 ( .s ({signal_2540, signal_2538}), .b ({signal_1312, signal_601}), .a ({signal_1213, signal_502}), .clk ( clk ), .r ( Fresh[586] ), .c ({signal_1490, signal_778}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_763 ( .s ({signal_2540, signal_2538}), .b ({signal_1133, signal_422}), .a ({signal_1214, signal_503}), .clk ( clk ), .r ( Fresh[587] ), .c ({signal_1491, signal_779}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_764 ( .s ({signal_2540, signal_2538}), .b ({signal_1170, signal_459}), .a ({signal_1145, signal_434}), .clk ( clk ), .r ( Fresh[588] ), .c ({signal_1492, signal_780}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_765 ( .s ({signal_2540, signal_2538}), .b ({signal_1153, signal_442}), .a ({signal_1143, signal_432}), .clk ( clk ), .r ( Fresh[589] ), .c ({signal_1493, signal_781}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_766 ( .s ({signal_2540, signal_2538}), .b ({signal_1355, signal_643}), .a ({signal_1301, signal_590}), .clk ( clk ), .r ( Fresh[590] ), .c ({signal_1494, signal_782}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_767 ( .s ({signal_2540, signal_2538}), .b ({signal_1147, signal_436}), .a ({signal_1311, signal_600}), .clk ( clk ), .r ( Fresh[591] ), .c ({signal_1495, signal_783}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_768 ( .s ({signal_2540, signal_2538}), .b ({signal_1191, signal_480}), .a ({signal_1290, signal_579}), .clk ( clk ), .r ( Fresh[592] ), .c ({signal_1496, signal_784}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_769 ( .s ({signal_2540, signal_2538}), .b ({signal_1273, signal_562}), .a ({signal_1352, signal_640}), .clk ( clk ), .r ( Fresh[593] ), .c ({signal_1497, signal_785}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_770 ( .s ({signal_2540, signal_2538}), .b ({signal_1309, signal_598}), .a ({signal_1169, signal_458}), .clk ( clk ), .r ( Fresh[594] ), .c ({signal_1498, signal_786}) ) ;
    buf_clk cell_1140 ( .C ( clk ), .D ( signal_2585 ), .Q ( signal_2586 ) ) ;
    buf_clk cell_1150 ( .C ( clk ), .D ( signal_2595 ), .Q ( signal_2596 ) ) ;
    buf_clk cell_1152 ( .C ( clk ), .D ( signal_2597 ), .Q ( signal_2598 ) ) ;
    buf_clk cell_1154 ( .C ( clk ), .D ( signal_2599 ), .Q ( signal_2600 ) ) ;
    buf_clk cell_1164 ( .C ( clk ), .D ( signal_2609 ), .Q ( signal_2610 ) ) ;
    buf_clk cell_1176 ( .C ( clk ), .D ( signal_2621 ), .Q ( signal_2622 ) ) ;
    buf_clk cell_1188 ( .C ( clk ), .D ( signal_2633 ), .Q ( signal_2634 ) ) ;
    buf_clk cell_1202 ( .C ( clk ), .D ( signal_2647 ), .Q ( signal_2648 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_1165 ( .C ( clk ), .D ( signal_2610 ), .Q ( signal_2611 ) ) ;
    buf_clk cell_1177 ( .C ( clk ), .D ( signal_2622 ), .Q ( signal_2623 ) ) ;
    buf_clk cell_1189 ( .C ( clk ), .D ( signal_2634 ), .Q ( signal_2635 ) ) ;
    buf_clk cell_1203 ( .C ( clk ), .D ( signal_2648 ), .Q ( signal_2649 ) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_771 ( .s ({signal_2596, signal_2586}), .b ({signal_1400, signal_688}), .a ({signal_1374, signal_662}), .clk ( clk ), .r ( Fresh[595] ), .c ({signal_1500, signal_787}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_772 ( .s ({signal_2596, signal_2586}), .b ({signal_1412, signal_700}), .a ({signal_1411, signal_699}), .clk ( clk ), .r ( Fresh[596] ), .c ({signal_1501, signal_788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_773 ( .s ({signal_2596, signal_2586}), .b ({signal_1494, signal_782}), .a ({signal_1488, signal_776}), .clk ( clk ), .r ( Fresh[597] ), .c ({signal_1502, signal_789}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_774 ( .s ({signal_2596, signal_2586}), .b ({signal_1396, signal_684}), .a ({signal_1440, signal_728}), .clk ( clk ), .r ( Fresh[598] ), .c ({signal_1503, signal_790}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_775 ( .s ({signal_2596, signal_2586}), .b ({signal_1381, signal_669}), .a ({signal_1384, signal_672}), .clk ( clk ), .r ( Fresh[599] ), .c ({signal_1504, signal_791}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_776 ( .s ({signal_2596, signal_2586}), .b ({signal_1383, signal_671}), .a ({signal_1390, signal_678}), .clk ( clk ), .r ( Fresh[600] ), .c ({signal_1505, signal_792}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_777 ( .s ({signal_2596, signal_2586}), .b ({signal_1388, signal_676}), .a ({signal_1458, signal_746}), .clk ( clk ), .r ( Fresh[601] ), .c ({signal_1506, signal_793}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_778 ( .s ({signal_2596, signal_2586}), .b ({signal_1493, signal_781}), .a ({signal_1391, signal_679}), .clk ( clk ), .r ( Fresh[602] ), .c ({signal_1507, signal_794}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_779 ( .s ({signal_2596, signal_2586}), .b ({signal_1439, signal_727}), .a ({signal_1469, signal_757}), .clk ( clk ), .r ( Fresh[603] ), .c ({signal_1508, signal_795}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_780 ( .s ({signal_2596, signal_2586}), .b ({signal_1459, signal_747}), .a ({signal_1477, signal_765}), .clk ( clk ), .r ( Fresh[604] ), .c ({signal_1509, signal_796}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_781 ( .s ({signal_2596, signal_2586}), .b ({signal_1397, signal_685}), .a ({signal_1473, signal_761}), .clk ( clk ), .r ( Fresh[605] ), .c ({signal_1510, signal_797}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_782 ( .s ({signal_2596, signal_2586}), .b ({signal_1380, signal_668}), .a ({signal_1444, signal_732}), .clk ( clk ), .r ( Fresh[606] ), .c ({signal_1511, signal_798}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_783 ( .s ({signal_2596, signal_2586}), .b ({signal_1467, signal_755}), .a ({signal_1387, signal_675}), .clk ( clk ), .r ( Fresh[607] ), .c ({signal_1512, signal_799}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_784 ( .s ({signal_2596, signal_2586}), .b ({signal_1437, signal_725}), .a ({signal_1438, signal_726}), .clk ( clk ), .r ( Fresh[608] ), .c ({signal_1513, signal_800}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_785 ( .s ({signal_2596, signal_2586}), .b ({signal_1496, signal_784}), .a ({signal_1465, signal_753}), .clk ( clk ), .r ( Fresh[609] ), .c ({signal_1514, signal_801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_786 ( .s ({signal_2596, signal_2586}), .b ({signal_1419, signal_707}), .a ({signal_1451, signal_739}), .clk ( clk ), .r ( Fresh[610] ), .c ({signal_1515, signal_802}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_787 ( .s ({signal_2596, signal_2586}), .b ({signal_1415, signal_703}), .a ({signal_1377, signal_665}), .clk ( clk ), .r ( Fresh[611] ), .c ({signal_1516, signal_803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_788 ( .s ({signal_2596, signal_2586}), .b ({signal_1442, signal_730}), .a ({signal_1492, signal_780}), .clk ( clk ), .r ( Fresh[612] ), .c ({signal_1517, signal_804}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_789 ( .s ({signal_2596, signal_2586}), .b ({signal_1445, signal_733}), .a ({signal_1422, signal_710}), .clk ( clk ), .r ( Fresh[613] ), .c ({signal_1518, signal_805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_790 ( .s ({signal_2596, signal_2586}), .b ({signal_1402, signal_690}), .a ({signal_1487, signal_775}), .clk ( clk ), .r ( Fresh[614] ), .c ({signal_1519, signal_806}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_791 ( .s ({signal_2596, signal_2586}), .b ({signal_1386, signal_674}), .a ({signal_1489, signal_777}), .clk ( clk ), .r ( Fresh[615] ), .c ({signal_1520, signal_807}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_792 ( .s ({signal_2596, signal_2586}), .b ({signal_1407, signal_695}), .a ({signal_1436, signal_724}), .clk ( clk ), .r ( Fresh[616] ), .c ({signal_1521, signal_808}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_793 ( .s ({signal_2596, signal_2586}), .b ({signal_1449, signal_737}), .a ({signal_1409, signal_697}), .clk ( clk ), .r ( Fresh[617] ), .c ({signal_1522, signal_809}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_794 ( .s ({signal_2596, signal_2586}), .b ({signal_1404, signal_692}), .a ({signal_1373, signal_661}), .clk ( clk ), .r ( Fresh[618] ), .c ({signal_1523, signal_810}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_795 ( .s ({signal_2596, signal_2586}), .b ({signal_1410, signal_698}), .a ({signal_1379, signal_667}), .clk ( clk ), .r ( Fresh[619] ), .c ({signal_1524, signal_811}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_796 ( .s ({signal_2596, signal_2586}), .b ({signal_1475, signal_763}), .a ({signal_1460, signal_748}), .clk ( clk ), .r ( Fresh[620] ), .c ({signal_1525, signal_812}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_797 ( .s ({signal_2596, signal_2586}), .b ({signal_1476, signal_764}), .a ({signal_1376, signal_664}), .clk ( clk ), .r ( Fresh[621] ), .c ({signal_1526, signal_813}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_798 ( .s ({signal_2596, signal_2586}), .b ({signal_1455, signal_743}), .a ({signal_1481, signal_769}), .clk ( clk ), .r ( Fresh[622] ), .c ({signal_1527, signal_814}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_799 ( .s ({signal_2596, signal_2586}), .b ({signal_1463, signal_751}), .a ({signal_1399, signal_687}), .clk ( clk ), .r ( Fresh[623] ), .c ({signal_1528, signal_815}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_800 ( .s ({signal_2596, signal_2586}), .b ({signal_1450, signal_738}), .a ({signal_1485, signal_773}), .clk ( clk ), .r ( Fresh[624] ), .c ({signal_1529, signal_816}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_801 ( .s ({signal_2596, signal_2586}), .b ({signal_1466, signal_754}), .a ({signal_1452, signal_740}), .clk ( clk ), .r ( Fresh[625] ), .c ({signal_1530, signal_817}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_802 ( .s ({signal_2596, signal_2586}), .b ({signal_1435, signal_723}), .a ({signal_1483, signal_771}), .clk ( clk ), .r ( Fresh[626] ), .c ({signal_1531, signal_818}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_803 ( .s ({signal_2596, signal_2586}), .b ({signal_1478, signal_766}), .a ({signal_1420, signal_708}), .clk ( clk ), .r ( Fresh[627] ), .c ({signal_1532, signal_819}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_804 ( .s ({signal_2596, signal_2586}), .b ({signal_1482, signal_770}), .a ({signal_1426, signal_714}), .clk ( clk ), .r ( Fresh[628] ), .c ({signal_1533, signal_820}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_805 ( .s ({signal_2596, signal_2586}), .b ({signal_1441, signal_729}), .a ({signal_1424, signal_712}), .clk ( clk ), .r ( Fresh[629] ), .c ({signal_1534, signal_821}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_806 ( .s ({signal_2596, signal_2586}), .b ({signal_1468, signal_756}), .a ({signal_1393, signal_681}), .clk ( clk ), .r ( Fresh[630] ), .c ({signal_1535, signal_822}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_807 ( .s ({signal_2596, signal_2586}), .b ({signal_1472, signal_760}), .a ({signal_1471, signal_759}), .clk ( clk ), .r ( Fresh[631] ), .c ({signal_1536, signal_823}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_808 ( .s ({signal_2596, signal_2586}), .b ({signal_1427, signal_715}), .a ({signal_1414, signal_702}), .clk ( clk ), .r ( Fresh[632] ), .c ({signal_1537, signal_824}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_809 ( .s ({signal_2596, signal_2586}), .b ({signal_1470, signal_758}), .a ({signal_1394, signal_682}), .clk ( clk ), .r ( Fresh[633] ), .c ({signal_1538, signal_825}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_810 ( .s ({signal_2596, signal_2586}), .b ({signal_1431, signal_719}), .a ({signal_1480, signal_768}), .clk ( clk ), .r ( Fresh[634] ), .c ({signal_1539, signal_826}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_811 ( .s ({signal_2596, signal_2586}), .b ({signal_1429, signal_717}), .a ({signal_1448, signal_736}), .clk ( clk ), .r ( Fresh[635] ), .c ({signal_1540, signal_827}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_812 ( .s ({signal_2596, signal_2586}), .b ({signal_1395, signal_683}), .a ({signal_1461, signal_749}), .clk ( clk ), .r ( Fresh[636] ), .c ({signal_1541, signal_828}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_813 ( .s ({signal_2596, signal_2586}), .b ({signal_1447, signal_735}), .a ({signal_1434, signal_722}), .clk ( clk ), .r ( Fresh[637] ), .c ({signal_1542, signal_829}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_814 ( .s ({signal_2596, signal_2586}), .b ({signal_1392, signal_680}), .a ({signal_1453, signal_741}), .clk ( clk ), .r ( Fresh[638] ), .c ({signal_1543, signal_830}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_815 ( .s ({signal_2596, signal_2586}), .b ({signal_1413, signal_701}), .a ({signal_1382, signal_670}), .clk ( clk ), .r ( Fresh[639] ), .c ({signal_1544, signal_831}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_816 ( .s ({signal_2596, signal_2586}), .b ({signal_1430, signal_718}), .a ({signal_1457, signal_745}), .clk ( clk ), .r ( Fresh[640] ), .c ({signal_1545, signal_832}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_817 ( .s ({signal_2596, signal_2586}), .b ({signal_1446, signal_734}), .a ({signal_1408, signal_696}), .clk ( clk ), .r ( Fresh[641] ), .c ({signal_1546, signal_833}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_818 ( .s ({signal_2596, signal_2586}), .b ({signal_1418, signal_706}), .a ({signal_1401, signal_689}), .clk ( clk ), .r ( Fresh[642] ), .c ({signal_1547, signal_834}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_819 ( .s ({signal_2596, signal_2586}), .b ({signal_1405, signal_693}), .a ({signal_1421, signal_709}), .clk ( clk ), .r ( Fresh[643] ), .c ({signal_1548, signal_835}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_820 ( .s ({signal_2596, signal_2586}), .b ({signal_1497, signal_785}), .a ({signal_1479, signal_767}), .clk ( clk ), .r ( Fresh[644] ), .c ({signal_1549, signal_836}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_821 ( .s ({signal_2596, signal_2586}), .b ({signal_1454, signal_742}), .a ({signal_1375, signal_663}), .clk ( clk ), .r ( Fresh[645] ), .c ({signal_1550, signal_837}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_822 ( .s ({signal_2596, signal_2586}), .b ({signal_2600, signal_2598}), .a ({signal_1425, signal_713}), .clk ( clk ), .r ( Fresh[646] ), .c ({signal_1551, signal_838}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_823 ( .s ({signal_2596, signal_2586}), .b ({signal_1433, signal_721}), .a ({signal_1474, signal_762}), .clk ( clk ), .r ( Fresh[647] ), .c ({signal_1552, signal_839}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_824 ( .s ({signal_2596, signal_2586}), .b ({signal_1389, signal_677}), .a ({signal_1423, signal_711}), .clk ( clk ), .r ( Fresh[648] ), .c ({signal_1553, signal_840}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_825 ( .s ({signal_2596, signal_2586}), .b ({signal_1491, signal_779}), .a ({signal_1464, signal_752}), .clk ( clk ), .r ( Fresh[649] ), .c ({signal_1554, signal_841}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_826 ( .s ({signal_2596, signal_2586}), .b ({signal_1484, signal_772}), .a ({signal_1378, signal_666}), .clk ( clk ), .r ( Fresh[650] ), .c ({signal_1555, signal_842}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_827 ( .s ({signal_2596, signal_2586}), .b ({signal_1416, signal_704}), .a ({signal_1462, signal_750}), .clk ( clk ), .r ( Fresh[651] ), .c ({signal_1556, signal_843}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_828 ( .s ({signal_2596, signal_2586}), .b ({signal_1456, signal_744}), .a ({signal_1498, signal_786}), .clk ( clk ), .r ( Fresh[652] ), .c ({signal_1557, signal_844}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_829 ( .s ({signal_2596, signal_2586}), .b ({signal_1372, signal_660}), .a ({signal_1398, signal_686}), .clk ( clk ), .r ( Fresh[653] ), .c ({signal_1558, signal_845}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_830 ( .s ({signal_2596, signal_2586}), .b ({signal_1428, signal_716}), .a ({signal_1406, signal_694}), .clk ( clk ), .r ( Fresh[654] ), .c ({signal_1559, signal_846}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_831 ( .s ({signal_2596, signal_2586}), .b ({signal_1417, signal_705}), .a ({signal_1403, signal_691}), .clk ( clk ), .r ( Fresh[655] ), .c ({signal_1560, signal_847}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_832 ( .s ({signal_2596, signal_2586}), .b ({signal_1443, signal_731}), .a ({signal_1432, signal_720}), .clk ( clk ), .r ( Fresh[656] ), .c ({signal_1561, signal_848}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_833 ( .s ({signal_2596, signal_2586}), .b ({signal_1486, signal_774}), .a ({signal_1385, signal_673}), .clk ( clk ), .r ( Fresh[657] ), .c ({signal_1562, signal_849}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_834 ( .s ({signal_2596, signal_2586}), .b ({signal_1495, signal_783}), .a ({signal_1490, signal_778}), .clk ( clk ), .r ( Fresh[658] ), .c ({signal_1563, signal_850}) ) ;
    buf_clk cell_1166 ( .C ( clk ), .D ( signal_2611 ), .Q ( signal_2612 ) ) ;
    buf_clk cell_1178 ( .C ( clk ), .D ( signal_2623 ), .Q ( signal_2624 ) ) ;
    buf_clk cell_1190 ( .C ( clk ), .D ( signal_2635 ), .Q ( signal_2636 ) ) ;
    buf_clk cell_1204 ( .C ( clk ), .D ( signal_2649 ), .Q ( signal_2650 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_1191 ( .C ( clk ), .D ( signal_2636 ), .Q ( signal_2637 ) ) ;
    buf_clk cell_1205 ( .C ( clk ), .D ( signal_2650 ), .Q ( signal_2651 ) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_835 ( .s ({signal_2624, signal_2612}), .b ({signal_1510, signal_797}), .a ({signal_1502, signal_789}), .clk ( clk ), .r ( Fresh[659] ), .c ({signal_1565, signal_851}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_836 ( .s ({signal_2624, signal_2612}), .b ({signal_1519, signal_806}), .a ({signal_1520, signal_807}), .clk ( clk ), .r ( Fresh[660] ), .c ({signal_1566, signal_852}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_837 ( .s ({signal_2624, signal_2612}), .b ({signal_1550, signal_837}), .a ({signal_1523, signal_810}), .clk ( clk ), .r ( Fresh[661] ), .c ({signal_1567, signal_853}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_838 ( .s ({signal_2624, signal_2612}), .b ({signal_1528, signal_815}), .a ({signal_1540, signal_827}), .clk ( clk ), .r ( Fresh[662] ), .c ({signal_1568, signal_854}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_839 ( .s ({signal_2624, signal_2612}), .b ({signal_1534, signal_821}), .a ({signal_1517, signal_804}), .clk ( clk ), .r ( Fresh[663] ), .c ({signal_1569, signal_855}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_840 ( .s ({signal_2624, signal_2612}), .b ({signal_1504, signal_791}), .a ({signal_1542, signal_829}), .clk ( clk ), .r ( Fresh[664] ), .c ({signal_1570, signal_856}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_841 ( .s ({signal_2624, signal_2612}), .b ({signal_1503, signal_790}), .a ({signal_1546, signal_833}), .clk ( clk ), .r ( Fresh[665] ), .c ({signal_1571, signal_857}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_842 ( .s ({signal_2624, signal_2612}), .b ({signal_1560, signal_847}), .a ({signal_1524, signal_811}), .clk ( clk ), .r ( Fresh[666] ), .c ({signal_1572, signal_858}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_843 ( .s ({signal_2624, signal_2612}), .b ({signal_1552, signal_839}), .a ({signal_1554, signal_841}), .clk ( clk ), .r ( Fresh[667] ), .c ({signal_1573, signal_859}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_844 ( .s ({signal_2624, signal_2612}), .b ({signal_1553, signal_840}), .a ({signal_1559, signal_846}), .clk ( clk ), .r ( Fresh[668] ), .c ({signal_1574, signal_860}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_845 ( .s ({signal_2624, signal_2612}), .b ({signal_1562, signal_849}), .a ({signal_1547, signal_834}), .clk ( clk ), .r ( Fresh[669] ), .c ({signal_1575, signal_861}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_846 ( .s ({signal_2624, signal_2612}), .b ({signal_1506, signal_793}), .a ({signal_1555, signal_842}), .clk ( clk ), .r ( Fresh[670] ), .c ({signal_1576, signal_862}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_847 ( .s ({signal_2624, signal_2612}), .b ({signal_1526, signal_813}), .a ({signal_1507, signal_794}), .clk ( clk ), .r ( Fresh[671] ), .c ({signal_1577, signal_863}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_848 ( .s ({signal_2624, signal_2612}), .b ({signal_1509, signal_796}), .a ({signal_1508, signal_795}), .clk ( clk ), .r ( Fresh[672] ), .c ({signal_1578, signal_864}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_849 ( .s ({signal_2624, signal_2612}), .b ({signal_1563, signal_850}), .a ({signal_1529, signal_816}), .clk ( clk ), .r ( Fresh[673] ), .c ({signal_1579, signal_865}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_850 ( .s ({signal_2624, signal_2612}), .b ({signal_1551, signal_838}), .a ({signal_1535, signal_822}), .clk ( clk ), .r ( Fresh[674] ), .c ({signal_1580, signal_866}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_851 ( .s ({signal_2624, signal_2612}), .b ({signal_1501, signal_788}), .a ({signal_1557, signal_844}), .clk ( clk ), .r ( Fresh[675] ), .c ({signal_1581, signal_867}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_852 ( .s ({signal_2624, signal_2612}), .b ({signal_1527, signal_814}), .a ({signal_1511, signal_798}), .clk ( clk ), .r ( Fresh[676] ), .c ({signal_1582, signal_868}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_853 ( .s ({signal_2624, signal_2612}), .b ({signal_1518, signal_805}), .a ({signal_1530, signal_817}), .clk ( clk ), .r ( Fresh[677] ), .c ({signal_1583, signal_869}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_854 ( .s ({signal_2624, signal_2612}), .b ({signal_1539, signal_826}), .a ({signal_1549, signal_836}), .clk ( clk ), .r ( Fresh[678] ), .c ({signal_1584, signal_870}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_855 ( .s ({signal_2624, signal_2612}), .b ({signal_1558, signal_845}), .a ({signal_1532, signal_819}), .clk ( clk ), .r ( Fresh[679] ), .c ({signal_1585, signal_871}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_856 ( .s ({signal_2624, signal_2612}), .b ({signal_1515, signal_802}), .a ({signal_1525, signal_812}), .clk ( clk ), .r ( Fresh[680] ), .c ({signal_1586, signal_872}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_857 ( .s ({signal_2624, signal_2612}), .b ({signal_1516, signal_803}), .a ({signal_1561, signal_848}), .clk ( clk ), .r ( Fresh[681] ), .c ({signal_1587, signal_873}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_858 ( .s ({signal_2624, signal_2612}), .b ({signal_1512, signal_799}), .a ({signal_1538, signal_825}), .clk ( clk ), .r ( Fresh[682] ), .c ({signal_1588, signal_874}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_859 ( .s ({signal_2624, signal_2612}), .b ({signal_1533, signal_820}), .a ({signal_1522, signal_809}), .clk ( clk ), .r ( Fresh[683] ), .c ({signal_1589, signal_875}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_860 ( .s ({signal_2624, signal_2612}), .b ({signal_1544, signal_831}), .a ({signal_1531, signal_818}), .clk ( clk ), .r ( Fresh[684] ), .c ({signal_1590, signal_876}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_861 ( .s ({signal_2624, signal_2612}), .b ({signal_1536, signal_823}), .a ({signal_1513, signal_800}), .clk ( clk ), .r ( Fresh[685] ), .c ({signal_1591, signal_877}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_862 ( .s ({signal_2624, signal_2612}), .b ({signal_1514, signal_801}), .a ({signal_1505, signal_792}), .clk ( clk ), .r ( Fresh[686] ), .c ({signal_1592, signal_878}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_863 ( .s ({signal_2624, signal_2612}), .b ({signal_1500, signal_787}), .a ({signal_1545, signal_832}), .clk ( clk ), .r ( Fresh[687] ), .c ({signal_1593, signal_879}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_864 ( .s ({signal_2624, signal_2612}), .b ({signal_1541, signal_828}), .a ({signal_1543, signal_830}), .clk ( clk ), .r ( Fresh[688] ), .c ({signal_1594, signal_880}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_865 ( .s ({signal_2624, signal_2612}), .b ({signal_1537, signal_824}), .a ({signal_1556, signal_843}), .clk ( clk ), .r ( Fresh[689] ), .c ({signal_1595, signal_881}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_866 ( .s ({signal_2624, signal_2612}), .b ({signal_1521, signal_808}), .a ({signal_1548, signal_835}), .clk ( clk ), .r ( Fresh[690] ), .c ({signal_1596, signal_882}) ) ;
    buf_clk cell_1192 ( .C ( clk ), .D ( signal_2637 ), .Q ( signal_2638 ) ) ;
    buf_clk cell_1206 ( .C ( clk ), .D ( signal_2651 ), .Q ( signal_2652 ) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_867 ( .s ({signal_2652, signal_2638}), .b ({signal_1570, signal_856}), .a ({signal_1588, signal_874}), .clk ( clk ), .r ( Fresh[691] ), .c ({signal_1598, signal_883}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_868 ( .s ({signal_2652, signal_2638}), .b ({signal_1579, signal_865}), .a ({signal_1586, signal_872}), .clk ( clk ), .r ( Fresh[692] ), .c ({signal_1599, signal_884}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_869 ( .s ({signal_2652, signal_2638}), .b ({signal_1578, signal_864}), .a ({signal_1582, signal_868}), .clk ( clk ), .r ( Fresh[693] ), .c ({signal_1600, signal_885}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_870 ( .s ({signal_2652, signal_2638}), .b ({signal_1572, signal_858}), .a ({signal_1569, signal_855}), .clk ( clk ), .r ( Fresh[694] ), .c ({signal_1601, signal_886}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_871 ( .s ({signal_2652, signal_2638}), .b ({signal_1592, signal_878}), .a ({signal_1568, signal_854}), .clk ( clk ), .r ( Fresh[695] ), .c ({signal_1602, signal_887}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_872 ( .s ({signal_2652, signal_2638}), .b ({signal_1576, signal_862}), .a ({signal_1585, signal_871}), .clk ( clk ), .r ( Fresh[696] ), .c ({signal_1603, signal_888}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_873 ( .s ({signal_2652, signal_2638}), .b ({signal_1594, signal_880}), .a ({signal_1591, signal_877}), .clk ( clk ), .r ( Fresh[697] ), .c ({signal_1604, signal_889}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_874 ( .s ({signal_2652, signal_2638}), .b ({signal_1596, signal_882}), .a ({signal_1581, signal_867}), .clk ( clk ), .r ( Fresh[698] ), .c ({signal_1605, signal_890}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_875 ( .s ({signal_2652, signal_2638}), .b ({signal_1566, signal_852}), .a ({signal_1573, signal_859}), .clk ( clk ), .r ( Fresh[699] ), .c ({signal_1606, signal_891}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_876 ( .s ({signal_2652, signal_2638}), .b ({signal_1583, signal_869}), .a ({signal_1571, signal_857}), .clk ( clk ), .r ( Fresh[700] ), .c ({signal_1607, signal_892}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_877 ( .s ({signal_2652, signal_2638}), .b ({signal_1595, signal_881}), .a ({signal_1574, signal_860}), .clk ( clk ), .r ( Fresh[701] ), .c ({signal_1608, signal_893}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_878 ( .s ({signal_2652, signal_2638}), .b ({signal_1580, signal_866}), .a ({signal_1577, signal_863}), .clk ( clk ), .r ( Fresh[702] ), .c ({signal_1609, signal_894}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_879 ( .s ({signal_2652, signal_2638}), .b ({signal_1565, signal_851}), .a ({signal_1593, signal_879}), .clk ( clk ), .r ( Fresh[703] ), .c ({signal_1610, signal_895}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_880 ( .s ({signal_2652, signal_2638}), .b ({signal_1584, signal_870}), .a ({signal_1567, signal_853}), .clk ( clk ), .r ( Fresh[704] ), .c ({signal_1611, signal_896}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_881 ( .s ({signal_2652, signal_2638}), .b ({signal_1589, signal_875}), .a ({signal_1587, signal_873}), .clk ( clk ), .r ( Fresh[705] ), .c ({signal_1612, signal_897}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_882 ( .s ({signal_2652, signal_2638}), .b ({signal_1590, signal_876}), .a ({signal_1575, signal_861}), .clk ( clk ), .r ( Fresh[706] ), .c ({signal_1613, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_883 ( .s ( 1'b1 ), .b ({signal_1600, signal_885}), .a ({signal_1613, signal_898}), .c ({signal_1614, signal_165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_884 ( .s ( 1'b1 ), .b ({signal_1598, signal_883}), .a ({signal_1599, signal_884}), .c ({signal_1615, signal_161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_885 ( .s ( 1'b1 ), .b ({signal_1604, signal_889}), .a ({signal_1609, signal_894}), .c ({signal_1616, signal_166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_886 ( .s ( 1'b1 ), .b ({signal_1601, signal_886}), .a ({signal_1602, signal_887}), .c ({signal_1617, signal_160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_887 ( .s ( 1'b1 ), .b ({signal_1603, signal_888}), .a ({signal_1605, signal_890}), .c ({signal_1618, signal_164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_888 ( .s ( 1'b1 ), .b ({signal_1607, signal_892}), .a ({signal_1608, signal_893}), .c ({signal_1619, signal_167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_889 ( .s ( 1'b1 ), .b ({signal_1612, signal_897}), .a ({signal_1606, signal_891}), .c ({signal_1620, signal_163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_890 ( .s ( 1'b1 ), .b ({signal_1610, signal_895}), .a ({signal_1611, signal_896}), .c ({signal_1621, signal_162}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_1617, signal_160}), .Q ({Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_1615, signal_161}), .Q ({Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_1621, signal_162}), .Q ({Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_1620, signal_163}), .Q ({Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_1618, signal_164}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_1614, signal_165}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_1616, signal_166}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_1619, signal_167}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
